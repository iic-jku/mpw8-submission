magic
tech sky130A
magscale 1 2
timestamp 1670618893
<< viali >>
rect 2145 57545 2179 57579
rect 11161 57545 11195 57579
rect 13737 57545 13771 57579
rect 16221 57545 16255 57579
rect 17049 57545 17083 57579
rect 22477 57545 22511 57579
rect 25421 57545 25455 57579
rect 26617 57545 26651 57579
rect 29193 57545 29227 57579
rect 34253 57545 34287 57579
rect 41429 57545 41463 57579
rect 42625 57545 42659 57579
rect 46213 57545 46247 57579
rect 1961 57409 1995 57443
rect 3433 57409 3467 57443
rect 4353 57409 4387 57443
rect 6009 57409 6043 57443
rect 6561 57409 6595 57443
rect 8585 57409 8619 57443
rect 9137 57409 9171 57443
rect 9873 57409 9907 57443
rect 10333 57409 10367 57443
rect 11713 57409 11747 57443
rect 12725 57409 12759 57443
rect 14289 57409 14323 57443
rect 15117 57409 15151 57443
rect 16865 57409 16899 57443
rect 17509 57409 17543 57443
rect 18245 57409 18279 57443
rect 18705 57409 18739 57443
rect 19901 57409 19935 57443
rect 20637 57409 20671 57443
rect 21097 57409 21131 57443
rect 22293 57409 22327 57443
rect 23029 57409 23063 57443
rect 23489 57409 23523 57443
rect 24685 57409 24719 57443
rect 26065 57409 26099 57443
rect 27353 57409 27387 57443
rect 28273 57409 28307 57443
rect 29929 57409 29963 57443
rect 30665 57409 30699 57443
rect 31309 57409 31343 57443
rect 32321 57409 32355 57443
rect 33057 57409 33091 57443
rect 33701 57409 33735 57443
rect 35081 57409 35115 57443
rect 35541 57409 35575 57443
rect 36829 57409 36863 57443
rect 38025 57409 38059 57443
rect 38485 57409 38519 57443
rect 39221 57409 39255 57443
rect 40417 57409 40451 57443
rect 40877 57409 40911 57443
rect 41613 57409 41647 57443
rect 42809 57409 42843 57443
rect 43269 57409 43303 57443
rect 44005 57409 44039 57443
rect 44465 57409 44499 57443
rect 45385 57409 45419 57443
rect 46397 57409 46431 57443
rect 46857 57409 46891 57443
rect 47961 57409 47995 57443
rect 48789 57409 48823 57443
rect 49249 57409 49283 57443
rect 50537 57409 50571 57443
rect 51181 57409 51215 57443
rect 51641 57409 51675 57443
rect 52377 57409 52411 57443
rect 53573 57409 53607 57443
rect 54033 57409 54067 57443
rect 54769 57409 54803 57443
rect 55965 57409 55999 57443
rect 56425 57409 56459 57443
rect 57161 57409 57195 57443
rect 58357 57409 58391 57443
rect 3157 57341 3191 57375
rect 5733 57341 5767 57375
rect 8309 57341 8343 57375
rect 15301 57273 15335 57307
rect 17693 57273 17727 57307
rect 23673 57273 23707 57307
rect 30849 57273 30883 57307
rect 47777 57273 47811 57307
rect 50997 57273 51031 57307
rect 4537 57205 4571 57239
rect 9321 57205 9355 57239
rect 10517 57205 10551 57239
rect 11897 57205 11931 57239
rect 12909 57205 12943 57239
rect 14473 57205 14507 57239
rect 18889 57205 18923 57239
rect 20085 57205 20119 57239
rect 21281 57205 21315 57239
rect 24869 57205 24903 57239
rect 25881 57205 25915 57239
rect 27169 57205 27203 57239
rect 28457 57205 28491 57239
rect 29745 57205 29779 57239
rect 32505 57205 32539 57239
rect 33241 57205 33275 57239
rect 34897 57205 34931 57239
rect 35725 57205 35759 57239
rect 36645 57205 36679 57239
rect 37841 57205 37875 57239
rect 39037 57205 39071 57239
rect 40233 57205 40267 57239
rect 43821 57205 43855 57239
rect 45201 57205 45235 57239
rect 48605 57205 48639 57239
rect 50353 57205 50387 57239
rect 52193 57205 52227 57239
rect 53389 57205 53423 57239
rect 54585 57205 54619 57239
rect 55781 57205 55815 57239
rect 56977 57205 57011 57239
rect 58173 57205 58207 57239
rect 1869 57001 1903 57035
rect 3341 57001 3375 57035
rect 4261 57001 4295 57035
rect 8493 57001 8527 57035
rect 9137 57001 9171 57035
rect 12633 57001 12667 57035
rect 15025 57001 15059 57035
rect 17417 57001 17451 57035
rect 19809 57001 19843 57035
rect 22201 57001 22235 57035
rect 24593 57001 24627 57035
rect 28181 57001 28215 57035
rect 32137 57001 32171 57035
rect 35357 57001 35391 57035
rect 36553 57001 36587 57035
rect 38117 57001 38151 57035
rect 41337 57001 41371 57035
rect 45201 57001 45235 57035
rect 47593 57001 47627 57035
rect 50353 57001 50387 57035
rect 52101 57001 52135 57035
rect 54493 57001 54527 57035
rect 56425 57001 56459 57035
rect 21557 56933 21591 56967
rect 43269 56933 43303 56967
rect 6285 56865 6319 56899
rect 6745 56865 6779 56899
rect 29745 56865 29779 56899
rect 55873 56865 55907 56899
rect 7021 56797 7055 56831
rect 29837 56797 29871 56831
rect 30021 56797 30055 56831
rect 38764 56797 38798 56831
rect 38885 56797 38919 56831
rect 38996 56797 39030 56831
rect 39129 56797 39163 56831
rect 43407 56797 43441 56831
rect 43545 56797 43579 56831
rect 43820 56797 43854 56831
rect 43913 56797 43947 56831
rect 57069 56797 57103 56831
rect 57529 56797 57563 56831
rect 58357 56797 58391 56831
rect 21189 56729 21223 56763
rect 21373 56729 21407 56763
rect 43637 56729 43671 56763
rect 30205 56661 30239 56695
rect 38577 56661 38611 56695
rect 56885 56661 56919 56695
rect 57713 56661 57747 56695
rect 58173 56661 58207 56695
rect 26525 56457 26559 56491
rect 30665 56457 30699 56491
rect 34437 56457 34471 56491
rect 57161 56457 57195 56491
rect 21281 56389 21315 56423
rect 22201 56389 22235 56423
rect 25421 56389 25455 56423
rect 26249 56389 26283 56423
rect 27353 56389 27387 56423
rect 29121 56389 29155 56423
rect 30297 56389 30331 56423
rect 31309 56389 31343 56423
rect 32873 56389 32907 56423
rect 34713 56389 34747 56423
rect 34805 56389 34839 56423
rect 35817 56389 35851 56423
rect 35909 56389 35943 56423
rect 43545 56389 43579 56423
rect 56701 56389 56735 56423
rect 21097 56321 21131 56355
rect 22017 56321 22051 56355
rect 23760 56321 23794 56355
rect 23857 56321 23891 56355
rect 23949 56321 23983 56355
rect 24132 56321 24166 56355
rect 24225 56321 24259 56355
rect 24961 56321 24995 56355
rect 25237 56321 25271 56355
rect 25881 56321 25915 56355
rect 25974 56321 26008 56355
rect 26157 56321 26191 56355
rect 26387 56321 26421 56355
rect 27215 56321 27249 56355
rect 27445 56321 27479 56355
rect 27542 56321 27576 56355
rect 28733 56321 28767 56355
rect 28826 56321 28860 56355
rect 28963 56321 28997 56355
rect 29239 56321 29273 56355
rect 30021 56321 30055 56355
rect 30169 56321 30203 56355
rect 30389 56321 30423 56355
rect 30486 56321 30520 56355
rect 31125 56321 31159 56355
rect 31401 56321 31435 56355
rect 31545 56321 31579 56355
rect 32776 56321 32810 56355
rect 32965 56321 32999 56355
rect 33148 56321 33182 56355
rect 33241 56321 33275 56355
rect 34616 56321 34650 56355
rect 34988 56321 35022 56355
rect 35081 56321 35115 56355
rect 35720 56321 35754 56355
rect 36092 56321 36126 56355
rect 36185 56321 36219 56355
rect 37657 56321 37691 56355
rect 37749 56321 37783 56355
rect 37933 56321 37967 56355
rect 38025 56321 38059 56355
rect 38669 56321 38703 56355
rect 38761 56321 38795 56355
rect 38945 56321 38979 56355
rect 39037 56321 39071 56355
rect 40780 56321 40814 56355
rect 40877 56321 40911 56355
rect 40969 56321 41003 56355
rect 41152 56321 41186 56355
rect 41245 56321 41279 56355
rect 43315 56321 43349 56355
rect 43453 56321 43487 56355
rect 43728 56321 43762 56355
rect 43821 56321 43855 56355
rect 56149 56321 56183 56355
rect 58357 56321 58391 56355
rect 21465 56185 21499 56219
rect 29377 56185 29411 56219
rect 31677 56185 31711 56219
rect 35541 56185 35575 56219
rect 40601 56185 40635 56219
rect 22385 56117 22419 56151
rect 23581 56117 23615 56151
rect 25053 56117 25087 56151
rect 27721 56117 27755 56151
rect 32597 56117 32631 56151
rect 37473 56117 37507 56151
rect 38485 56117 38519 56151
rect 43177 56117 43211 56151
rect 58173 56117 58207 56151
rect 22845 55913 22879 55947
rect 24593 55913 24627 55947
rect 28825 55913 28859 55947
rect 32689 55913 32723 55947
rect 38485 55913 38519 55947
rect 57161 55913 57195 55947
rect 23949 55845 23983 55879
rect 30297 55845 30331 55879
rect 35633 55845 35667 55879
rect 41153 55845 41187 55879
rect 43269 55845 43303 55879
rect 25053 55777 25087 55811
rect 28365 55777 28399 55811
rect 30941 55777 30975 55811
rect 1869 55709 1903 55743
rect 21373 55709 21407 55743
rect 23397 55709 23431 55743
rect 23581 55709 23615 55743
rect 23673 55709 23707 55743
rect 23817 55709 23851 55743
rect 24777 55709 24811 55743
rect 24961 55709 24995 55743
rect 26985 55709 27019 55743
rect 28457 55709 28491 55743
rect 28641 55709 28675 55743
rect 29745 55709 29779 55743
rect 29929 55709 29963 55743
rect 30165 55709 30199 55743
rect 32868 55709 32902 55743
rect 32965 55709 32999 55743
rect 33240 55709 33274 55743
rect 33333 55709 33367 55743
rect 35771 55709 35805 55743
rect 35909 55709 35943 55743
rect 36184 55709 36218 55743
rect 36277 55709 36311 55743
rect 38661 55709 38695 55743
rect 38761 55709 38795 55743
rect 38945 55709 38979 55743
rect 39047 55687 39081 55721
rect 41332 55709 41366 55743
rect 41420 55709 41454 55743
rect 41704 55709 41738 55743
rect 41797 55709 41831 55743
rect 43407 55709 43441 55743
rect 43637 55709 43671 55743
rect 43820 55709 43854 55743
rect 43913 55709 43947 55743
rect 57713 55709 57747 55743
rect 58357 55709 58391 55743
rect 21189 55641 21223 55675
rect 21557 55641 21591 55675
rect 30021 55641 30055 55675
rect 33057 55641 33091 55675
rect 36001 55641 36035 55675
rect 41521 55641 41555 55675
rect 43545 55641 43579 55675
rect 1685 55573 1719 55607
rect 2329 55573 2363 55607
rect 58173 55573 58207 55607
rect 42625 55369 42659 55403
rect 58173 55369 58207 55403
rect 29561 55301 29595 55335
rect 42901 55301 42935 55335
rect 1869 55233 1903 55267
rect 2421 55233 2455 55267
rect 22017 55233 22051 55267
rect 22201 55233 22235 55267
rect 22385 55233 22419 55267
rect 38485 55233 38519 55267
rect 39589 55233 39623 55267
rect 42763 55233 42797 55267
rect 42993 55233 43027 55267
rect 43176 55233 43210 55267
rect 43269 55233 43303 55267
rect 57529 55233 57563 55267
rect 58357 55233 58391 55267
rect 1685 55029 1719 55063
rect 32413 55029 32447 55063
rect 26065 54825 26099 54859
rect 32781 54825 32815 54859
rect 32965 54825 32999 54859
rect 37473 54825 37507 54859
rect 25697 54689 25731 54723
rect 36921 54689 36955 54723
rect 21833 54621 21867 54655
rect 25881 54621 25915 54655
rect 26157 54621 26191 54655
rect 26617 54621 26651 54655
rect 26710 54621 26744 54655
rect 26893 54621 26927 54655
rect 27082 54621 27116 54655
rect 32413 54621 32447 54655
rect 35035 54621 35069 54655
rect 35448 54621 35482 54655
rect 35541 54621 35575 54655
rect 37657 54621 37691 54655
rect 37749 54621 37783 54655
rect 37933 54621 37967 54655
rect 38025 54621 38059 54655
rect 38669 54621 38703 54655
rect 39313 54621 39347 54655
rect 40601 54621 40635 54655
rect 21649 54553 21683 54587
rect 26985 54553 27019 54587
rect 35173 54553 35207 54587
rect 35265 54553 35299 54587
rect 22017 54485 22051 54519
rect 27261 54485 27295 54519
rect 31861 54485 31895 54519
rect 32781 54485 32815 54519
rect 34897 54485 34931 54519
rect 38761 54485 38795 54519
rect 40049 54485 40083 54519
rect 58357 54485 58391 54519
rect 26525 54281 26559 54315
rect 27738 54281 27772 54315
rect 31769 54281 31803 54315
rect 32505 54281 32539 54315
rect 34529 54281 34563 54315
rect 36277 54281 36311 54315
rect 38945 54281 38979 54315
rect 40325 54281 40359 54315
rect 41153 54281 41187 54315
rect 24501 54213 24535 54247
rect 25329 54213 25363 54247
rect 27353 54213 27387 54247
rect 27445 54213 27479 54247
rect 34897 54213 34931 54247
rect 40141 54213 40175 54247
rect 40785 54213 40819 54247
rect 40985 54213 41019 54247
rect 41613 54213 41647 54247
rect 34667 54179 34701 54213
rect 1869 54145 1903 54179
rect 24404 54145 24438 54179
rect 24593 54145 24627 54179
rect 24776 54145 24810 54179
rect 24869 54145 24903 54179
rect 25513 54145 25547 54179
rect 25697 54145 25731 54179
rect 25789 54145 25823 54179
rect 27169 54145 27203 54179
rect 27542 54145 27576 54179
rect 30205 54145 30239 54179
rect 32689 54145 32723 54179
rect 36453 54135 36487 54169
rect 36545 54145 36579 54179
rect 36737 54145 36771 54179
rect 36829 54145 36863 54179
rect 38301 54145 38335 54179
rect 38853 54145 38887 54179
rect 58357 54145 58391 54179
rect 29285 54077 29319 54111
rect 30113 54077 30147 54111
rect 32321 54077 32355 54111
rect 33977 54077 34011 54111
rect 1685 54009 1719 54043
rect 39773 54009 39807 54043
rect 2421 53941 2455 53975
rect 24225 53941 24259 53975
rect 29837 53941 29871 53975
rect 30021 53941 30055 53975
rect 32873 53941 32907 53975
rect 34713 53941 34747 53975
rect 40141 53941 40175 53975
rect 40969 53941 41003 53975
rect 58173 53941 58207 53975
rect 31493 53737 31527 53771
rect 31677 53737 31711 53771
rect 32321 53737 32355 53771
rect 37565 53737 37599 53771
rect 38485 53737 38519 53771
rect 40417 53737 40451 53771
rect 40601 53737 40635 53771
rect 25145 53669 25179 53703
rect 30481 53669 30515 53703
rect 40049 53669 40083 53703
rect 41061 53669 41095 53703
rect 1869 53533 1903 53567
rect 24593 53533 24627 53567
rect 24777 53533 24811 53567
rect 24966 53533 25000 53567
rect 29193 53533 29227 53567
rect 29745 53533 29779 53567
rect 30205 53533 30239 53567
rect 30573 53533 30607 53567
rect 32413 53533 32447 53567
rect 32597 53533 32631 53567
rect 33149 53533 33183 53567
rect 33885 53533 33919 53567
rect 39405 53533 39439 53567
rect 57713 53533 57747 53567
rect 58357 53533 58391 53567
rect 24869 53465 24903 53499
rect 31861 53465 31895 53499
rect 38209 53465 38243 53499
rect 40417 53465 40451 53499
rect 1685 53397 1719 53431
rect 2421 53397 2455 53431
rect 23949 53397 23983 53431
rect 31677 53397 31711 53431
rect 58173 53397 58207 53431
rect 29561 53193 29595 53227
rect 32597 53193 32631 53227
rect 40233 53193 40267 53227
rect 29929 53057 29963 53091
rect 32689 53057 32723 53091
rect 29377 52989 29411 53023
rect 29837 52989 29871 53023
rect 28825 52853 28859 52887
rect 39681 52853 39715 52887
rect 29101 52649 29135 52683
rect 1685 52581 1719 52615
rect 58173 52581 58207 52615
rect 1869 52445 1903 52479
rect 2421 52445 2455 52479
rect 57713 52445 57747 52479
rect 58357 52445 58391 52479
rect 1869 51969 1903 52003
rect 57529 51969 57563 52003
rect 58357 51969 58391 52003
rect 1685 51765 1719 51799
rect 2421 51765 2455 51799
rect 58173 51765 58207 51799
rect 58357 51221 58391 51255
rect 1869 50881 1903 50915
rect 58357 50881 58391 50915
rect 1685 50745 1719 50779
rect 2421 50677 2455 50711
rect 58173 50677 58207 50711
rect 1869 50269 1903 50303
rect 2329 50269 2363 50303
rect 57713 50269 57747 50303
rect 58357 50269 58391 50303
rect 1685 50133 1719 50167
rect 58173 50133 58207 50167
rect 1869 49181 1903 49215
rect 2421 49181 2455 49215
rect 57713 49181 57747 49215
rect 58357 49181 58391 49215
rect 1685 49045 1719 49079
rect 58173 49045 58207 49079
rect 1869 48705 1903 48739
rect 57529 48705 57563 48739
rect 58357 48705 58391 48739
rect 1685 48501 1719 48535
rect 2329 48501 2363 48535
rect 58173 48501 58207 48535
rect 58357 47957 58391 47991
rect 1869 47617 1903 47651
rect 58357 47617 58391 47651
rect 1685 47481 1719 47515
rect 2421 47413 2455 47447
rect 58173 47413 58207 47447
rect 58173 47141 58207 47175
rect 1869 47005 1903 47039
rect 57713 47005 57747 47039
rect 58357 47005 58391 47039
rect 2329 46937 2363 46971
rect 1685 46869 1719 46903
rect 1869 45917 1903 45951
rect 57713 45917 57747 45951
rect 58357 45917 58391 45951
rect 1685 45781 1719 45815
rect 2421 45781 2455 45815
rect 58173 45781 58207 45815
rect 1869 45441 1903 45475
rect 57529 45441 57563 45475
rect 58357 45441 58391 45475
rect 1685 45237 1719 45271
rect 2421 45237 2455 45271
rect 58173 45237 58207 45271
rect 58357 44693 58391 44727
rect 1869 44353 1903 44387
rect 58357 44353 58391 44387
rect 1685 44217 1719 44251
rect 2421 44149 2455 44183
rect 58173 44149 58207 44183
rect 1869 43741 1903 43775
rect 57713 43741 57747 43775
rect 58357 43741 58391 43775
rect 1685 43605 1719 43639
rect 2421 43605 2455 43639
rect 58173 43605 58207 43639
rect 1869 42653 1903 42687
rect 2421 42653 2455 42687
rect 57713 42653 57747 42687
rect 58357 42653 58391 42687
rect 1685 42517 1719 42551
rect 58173 42517 58207 42551
rect 1869 42177 1903 42211
rect 2421 42177 2455 42211
rect 57529 42177 57563 42211
rect 58357 42177 58391 42211
rect 1685 41973 1719 42007
rect 58173 41973 58207 42007
rect 58357 41429 58391 41463
rect 1869 41089 1903 41123
rect 58357 41089 58391 41123
rect 1685 40953 1719 40987
rect 2421 40885 2455 40919
rect 58173 40885 58207 40919
rect 1869 40477 1903 40511
rect 57713 40477 57747 40511
rect 58357 40477 58391 40511
rect 1685 40341 1719 40375
rect 2421 40341 2455 40375
rect 58173 40341 58207 40375
rect 58173 40137 58207 40171
rect 57529 40001 57563 40035
rect 58357 40001 58391 40035
rect 56425 39797 56459 39831
rect 1869 39389 1903 39423
rect 57253 39389 57287 39423
rect 57713 39389 57747 39423
rect 57621 39321 57655 39355
rect 57989 39321 58023 39355
rect 1685 39253 1719 39287
rect 2421 39253 2455 39287
rect 56149 39253 56183 39287
rect 56701 39253 56735 39287
rect 56885 39253 56919 39287
rect 56149 39049 56183 39083
rect 57253 39049 57287 39083
rect 58173 39049 58207 39083
rect 56517 38981 56551 39015
rect 1869 38913 1903 38947
rect 56885 38913 56919 38947
rect 56977 38913 57011 38947
rect 58357 38913 58391 38947
rect 1685 38709 1719 38743
rect 2421 38709 2455 38743
rect 55413 38709 55447 38743
rect 55965 38709 55999 38743
rect 57069 38505 57103 38539
rect 57621 38505 57655 38539
rect 55781 38165 55815 38199
rect 58357 38165 58391 38199
rect 58173 37961 58207 37995
rect 54677 37893 54711 37927
rect 55045 37893 55079 37927
rect 55505 37893 55539 37927
rect 55781 37893 55815 37927
rect 56425 37893 56459 37927
rect 1869 37825 1903 37859
rect 53941 37825 53975 37859
rect 55413 37825 55447 37859
rect 58357 37825 58391 37859
rect 1685 37689 1719 37723
rect 2421 37621 2455 37655
rect 54493 37621 54527 37655
rect 54309 37417 54343 37451
rect 57161 37281 57195 37315
rect 57713 37281 57747 37315
rect 1869 37213 1903 37247
rect 58357 37213 58391 37247
rect 1685 37077 1719 37111
rect 2421 37077 2455 37111
rect 58173 37077 58207 37111
rect 57529 36873 57563 36907
rect 58357 36737 58391 36771
rect 56609 36533 56643 36567
rect 58173 36533 58207 36567
rect 56885 36261 56919 36295
rect 1869 36125 1903 36159
rect 2421 36125 2455 36159
rect 57437 36125 57471 36159
rect 57897 36125 57931 36159
rect 56333 36057 56367 36091
rect 57805 36057 57839 36091
rect 1685 35989 1719 36023
rect 57069 35989 57103 36023
rect 58173 35989 58207 36023
rect 57529 35785 57563 35819
rect 1869 35649 1903 35683
rect 2421 35649 2455 35683
rect 56977 35649 57011 35683
rect 58357 35649 58391 35683
rect 1685 35445 1719 35479
rect 56241 35445 56275 35479
rect 58173 35445 58207 35479
rect 56977 35105 57011 35139
rect 57136 35105 57170 35139
rect 57253 35105 57287 35139
rect 57529 35105 57563 35139
rect 58173 35105 58207 35139
rect 57989 35037 58023 35071
rect 56333 34969 56367 35003
rect 55781 34901 55815 34935
rect 56701 34697 56735 34731
rect 1869 34561 1903 34595
rect 52377 34561 52411 34595
rect 55321 34561 55355 34595
rect 56241 34561 56275 34595
rect 57529 34561 57563 34595
rect 58357 34561 58391 34595
rect 2421 34493 2455 34527
rect 52101 34493 52135 34527
rect 53941 34493 53975 34527
rect 55045 34493 55079 34527
rect 55204 34493 55238 34527
rect 56057 34493 56091 34527
rect 1685 34425 1719 34459
rect 55597 34425 55631 34459
rect 54401 34357 54435 34391
rect 58173 34357 58207 34391
rect 54309 34153 54343 34187
rect 58173 34085 58207 34119
rect 1869 33949 1903 33983
rect 2329 33949 2363 33983
rect 57161 33949 57195 33983
rect 58357 33949 58391 33983
rect 1685 33813 1719 33847
rect 57713 33813 57747 33847
rect 57529 33609 57563 33643
rect 55045 33473 55079 33507
rect 58357 33473 58391 33507
rect 54769 33405 54803 33439
rect 58173 33269 58207 33303
rect 56425 32997 56459 33031
rect 1869 32861 1903 32895
rect 56977 32861 57011 32895
rect 57437 32861 57471 32895
rect 57345 32793 57379 32827
rect 1685 32725 1719 32759
rect 2421 32725 2455 32759
rect 55781 32725 55815 32759
rect 56609 32725 56643 32759
rect 57713 32725 57747 32759
rect 1869 32385 1903 32419
rect 2421 32385 2455 32419
rect 57529 32385 57563 32419
rect 58357 32385 58391 32419
rect 1685 32181 1719 32215
rect 56241 32181 56275 32215
rect 58173 32181 58207 32215
rect 55781 31909 55815 31943
rect 56885 31841 56919 31875
rect 57023 31841 57057 31875
rect 57161 31841 57195 31875
rect 57437 31841 57471 31875
rect 58081 31841 58115 31875
rect 56241 31773 56275 31807
rect 57897 31773 57931 31807
rect 57529 31433 57563 31467
rect 1869 31297 1903 31331
rect 53757 31297 53791 31331
rect 58173 31297 58207 31331
rect 53481 31229 53515 31263
rect 1685 31161 1719 31195
rect 2329 31093 2363 31127
rect 56149 31093 56183 31127
rect 58357 31093 58391 31127
rect 57713 30889 57747 30923
rect 1869 30685 1903 30719
rect 58173 30685 58207 30719
rect 1685 30549 1719 30583
rect 2421 30549 2455 30583
rect 58357 30549 58391 30583
rect 58357 30345 58391 30379
rect 12173 30277 12207 30311
rect 12909 30277 12943 30311
rect 56977 30277 57011 30311
rect 12081 30209 12115 30243
rect 12357 30141 12391 30175
rect 11069 30005 11103 30039
rect 11713 30005 11747 30039
rect 57437 30005 57471 30039
rect 9229 29665 9263 29699
rect 58357 29665 58391 29699
rect 1869 29597 1903 29631
rect 11437 29597 11471 29631
rect 56885 29597 56919 29631
rect 2421 29529 2455 29563
rect 9781 29529 9815 29563
rect 56517 29529 56551 29563
rect 57253 29529 57287 29563
rect 57345 29529 57379 29563
rect 57621 29529 57655 29563
rect 1685 29461 1719 29495
rect 11253 29461 11287 29495
rect 12541 29461 12575 29495
rect 56333 29461 56367 29495
rect 8493 29257 8527 29291
rect 9229 29257 9263 29291
rect 10701 29257 10735 29291
rect 11713 29257 11747 29291
rect 57345 29257 57379 29291
rect 58173 29257 58207 29291
rect 2421 29189 2455 29223
rect 56333 29189 56367 29223
rect 1869 29121 1903 29155
rect 8401 29121 8435 29155
rect 10609 29121 10643 29155
rect 57529 29121 57563 29155
rect 58357 29121 58391 29155
rect 7481 29053 7515 29087
rect 8677 29053 8711 29087
rect 10885 29053 10919 29087
rect 1685 28985 1719 29019
rect 10241 28985 10275 29019
rect 12265 28985 12299 29019
rect 56885 28985 56919 29019
rect 6837 28917 6871 28951
rect 8033 28917 8067 28951
rect 8585 28713 8619 28747
rect 16589 28713 16623 28747
rect 7849 28645 7883 28679
rect 11805 28645 11839 28679
rect 5917 28577 5951 28611
rect 9597 28577 9631 28611
rect 9689 28577 9723 28611
rect 12357 28577 12391 28611
rect 6193 28509 6227 28543
rect 7665 28509 7699 28543
rect 9505 28509 9539 28543
rect 10333 28509 10367 28543
rect 12265 28509 12299 28543
rect 56057 28509 56091 28543
rect 57161 28509 57195 28543
rect 57529 28509 57563 28543
rect 57621 28509 57655 28543
rect 6101 28441 6135 28475
rect 7021 28441 7055 28475
rect 13001 28441 13035 28475
rect 57897 28441 57931 28475
rect 1961 28373 1995 28407
rect 5273 28373 5307 28407
rect 6561 28373 6595 28407
rect 9137 28373 9171 28407
rect 11253 28373 11287 28407
rect 12173 28373 12207 28407
rect 56609 28373 56643 28407
rect 56793 28373 56827 28407
rect 4721 28169 4755 28203
rect 5641 28169 5675 28203
rect 8493 28169 8527 28203
rect 9137 28169 9171 28203
rect 12725 28169 12759 28203
rect 56977 28169 57011 28203
rect 57529 28169 57563 28203
rect 10149 28101 10183 28135
rect 11713 28101 11747 28135
rect 17325 28101 17359 28135
rect 1869 28033 1903 28067
rect 4813 28033 4847 28067
rect 6837 28033 6871 28067
rect 8125 28033 8159 28067
rect 8953 28033 8987 28067
rect 15945 28033 15979 28067
rect 17233 28033 17267 28067
rect 56425 28033 56459 28067
rect 58357 28033 58391 28067
rect 4537 27965 4571 27999
rect 7849 27965 7883 27999
rect 8033 27965 8067 27999
rect 17509 27965 17543 27999
rect 1685 27897 1719 27931
rect 2421 27897 2455 27931
rect 16865 27897 16899 27931
rect 58173 27897 58207 27931
rect 3433 27829 3467 27863
rect 5181 27829 5215 27863
rect 7021 27829 7055 27863
rect 9689 27829 9723 27863
rect 10793 27829 10827 27863
rect 13553 27829 13587 27863
rect 15761 27829 15795 27863
rect 18153 27829 18187 27863
rect 5917 27625 5951 27659
rect 9137 27557 9171 27591
rect 57713 27557 57747 27591
rect 2789 27489 2823 27523
rect 2881 27489 2915 27523
rect 3985 27489 4019 27523
rect 11161 27489 11195 27523
rect 11345 27489 11379 27523
rect 13277 27489 13311 27523
rect 14841 27489 14875 27523
rect 57161 27489 57195 27523
rect 57299 27489 57333 27523
rect 57437 27489 57471 27523
rect 58357 27489 58391 27523
rect 1869 27421 1903 27455
rect 5181 27421 5215 27455
rect 6377 27421 6411 27455
rect 8217 27421 8251 27455
rect 14657 27421 14691 27455
rect 16037 27421 16071 27455
rect 58173 27421 58207 27455
rect 2973 27353 3007 27387
rect 10149 27353 10183 27387
rect 12173 27353 12207 27387
rect 13185 27353 13219 27387
rect 16773 27353 16807 27387
rect 1685 27285 1719 27319
rect 3341 27285 3375 27319
rect 5365 27285 5399 27319
rect 8401 27285 8435 27319
rect 10701 27285 10735 27319
rect 11069 27285 11103 27319
rect 12725 27285 12759 27319
rect 13093 27285 13127 27319
rect 14289 27285 14323 27319
rect 14749 27285 14783 27319
rect 15485 27285 15519 27319
rect 17877 27285 17911 27319
rect 56517 27285 56551 27319
rect 5549 27081 5583 27115
rect 6561 27081 6595 27115
rect 11713 27081 11747 27115
rect 15117 27081 15151 27115
rect 56977 27081 57011 27115
rect 57529 27081 57563 27115
rect 58173 27081 58207 27115
rect 1685 27013 1719 27047
rect 11161 27013 11195 27047
rect 2513 26945 2547 26979
rect 4169 26945 4203 26979
rect 5641 26945 5675 26979
rect 7113 26945 7147 26979
rect 8769 26945 8803 26979
rect 9965 26945 9999 26979
rect 12265 26945 12299 26979
rect 13093 26945 13127 26979
rect 17325 26945 17359 26979
rect 58357 26945 58391 26979
rect 2237 26877 2271 26911
rect 2421 26877 2455 26911
rect 5365 26877 5399 26911
rect 13737 26877 13771 26911
rect 16313 26877 16347 26911
rect 17417 26877 17451 26911
rect 17601 26877 17635 26911
rect 12449 26809 12483 26843
rect 2881 26741 2915 26775
rect 3617 26741 3651 26775
rect 4353 26741 4387 26775
rect 6009 26741 6043 26775
rect 8953 26741 8987 26775
rect 10149 26741 10183 26775
rect 12909 26741 12943 26775
rect 16957 26741 16991 26775
rect 18245 26741 18279 26775
rect 10425 26537 10459 26571
rect 57161 26537 57195 26571
rect 4537 26469 4571 26503
rect 6193 26469 6227 26503
rect 11069 26469 11103 26503
rect 17049 26469 17083 26503
rect 44097 26469 44131 26503
rect 57621 26469 57655 26503
rect 58173 26469 58207 26503
rect 2329 26401 2363 26435
rect 2513 26401 2547 26435
rect 5549 26401 5583 26435
rect 5733 26401 5767 26435
rect 9873 26401 9907 26435
rect 17693 26401 17727 26435
rect 4077 26333 4111 26367
rect 7021 26333 7055 26367
rect 10885 26333 10919 26367
rect 16405 26333 16439 26367
rect 17417 26333 17451 26367
rect 44281 26333 44315 26367
rect 58357 26333 58391 26367
rect 5825 26265 5859 26299
rect 7757 26265 7791 26299
rect 9965 26265 9999 26299
rect 10057 26265 10091 26299
rect 11621 26265 11655 26299
rect 17509 26265 17543 26299
rect 18245 26265 18279 26299
rect 2605 26197 2639 26231
rect 2973 26197 3007 26231
rect 7205 26197 7239 26231
rect 16589 26197 16623 26231
rect 18797 26197 18831 26231
rect 1685 25993 1719 26027
rect 2329 25993 2363 26027
rect 3525 25993 3559 26027
rect 5917 25993 5951 26027
rect 57529 25993 57563 26027
rect 19349 25925 19383 25959
rect 1869 25857 1903 25891
rect 2881 25857 2915 25891
rect 6561 25857 6595 25891
rect 12725 25857 12759 25891
rect 17049 25857 17083 25891
rect 19257 25857 19291 25891
rect 56977 25857 57011 25891
rect 58357 25857 58391 25891
rect 19165 25789 19199 25823
rect 7205 25721 7239 25755
rect 58173 25721 58207 25755
rect 3065 25653 3099 25687
rect 4169 25653 4203 25687
rect 6745 25653 6779 25687
rect 10517 25653 10551 25687
rect 12909 25653 12943 25687
rect 16865 25653 16899 25687
rect 17969 25653 18003 25687
rect 18521 25653 18555 25687
rect 19717 25653 19751 25687
rect 20269 25653 20303 25687
rect 1685 25449 1719 25483
rect 3157 25449 3191 25483
rect 10885 25449 10919 25483
rect 5917 25381 5951 25415
rect 7665 25313 7699 25347
rect 57320 25313 57354 25347
rect 57713 25313 57747 25347
rect 58357 25313 58391 25347
rect 1869 25245 1903 25279
rect 2973 25245 3007 25279
rect 12633 25245 12667 25279
rect 19625 25245 19659 25279
rect 57161 25245 57195 25279
rect 57437 25245 57471 25279
rect 58173 25245 58207 25279
rect 2329 25177 2363 25211
rect 7389 25177 7423 25211
rect 12357 25177 12391 25211
rect 18613 25109 18647 25143
rect 19441 25109 19475 25143
rect 56517 25109 56551 25143
rect 1869 24769 1903 24803
rect 2973 24769 3007 24803
rect 5733 24769 5767 24803
rect 15393 24769 15427 24803
rect 19165 24769 19199 24803
rect 58357 24769 58391 24803
rect 5457 24701 5491 24735
rect 8309 24701 8343 24735
rect 9781 24701 9815 24735
rect 10057 24701 10091 24735
rect 15117 24701 15151 24735
rect 1685 24633 1719 24667
rect 3985 24633 4019 24667
rect 18981 24633 19015 24667
rect 58173 24633 58207 24667
rect 2421 24565 2455 24599
rect 3525 24565 3559 24599
rect 13645 24565 13679 24599
rect 18521 24565 18555 24599
rect 19625 24565 19659 24599
rect 56977 24565 57011 24599
rect 57437 24565 57471 24599
rect 12173 24361 12207 24395
rect 18521 24361 18555 24395
rect 19625 24361 19659 24395
rect 57713 24361 57747 24395
rect 58173 24293 58207 24327
rect 2789 24225 2823 24259
rect 2973 24225 3007 24259
rect 10425 24225 10459 24259
rect 10701 24225 10735 24259
rect 20269 24225 20303 24259
rect 1869 24157 1903 24191
rect 18797 24157 18831 24191
rect 57161 24157 57195 24191
rect 58357 24157 58391 24191
rect 3065 24089 3099 24123
rect 4537 24089 4571 24123
rect 20085 24089 20119 24123
rect 1685 24021 1719 24055
rect 3433 24021 3467 24055
rect 4077 24021 4111 24055
rect 19993 24021 20027 24055
rect 20821 24021 20855 24055
rect 3525 23817 3559 23851
rect 19533 23817 19567 23851
rect 58357 23817 58391 23851
rect 2237 23749 2271 23783
rect 2329 23681 2363 23715
rect 18613 23681 18647 23715
rect 2145 23613 2179 23647
rect 4169 23545 4203 23579
rect 2697 23477 2731 23511
rect 18429 23477 18463 23511
rect 20269 23477 20303 23511
rect 16037 23273 16071 23307
rect 18797 23273 18831 23307
rect 19441 23273 19475 23307
rect 58173 23273 58207 23307
rect 2513 23205 2547 23239
rect 17785 23137 17819 23171
rect 19901 23137 19935 23171
rect 20085 23137 20119 23171
rect 1869 23069 1903 23103
rect 2329 23069 2363 23103
rect 3985 23069 4019 23103
rect 57713 23069 57747 23103
rect 58357 23069 58391 23103
rect 17509 23001 17543 23035
rect 1685 22933 1719 22967
rect 3065 22933 3099 22967
rect 4169 22933 4203 22967
rect 19809 22933 19843 22967
rect 20637 22933 20671 22967
rect 2329 22729 2363 22763
rect 3709 22729 3743 22763
rect 8309 22729 8343 22763
rect 18613 22729 18647 22763
rect 58173 22729 58207 22763
rect 2237 22661 2271 22695
rect 3157 22661 3191 22695
rect 10057 22593 10091 22627
rect 57529 22593 57563 22627
rect 58357 22593 58391 22627
rect 2145 22525 2179 22559
rect 9781 22525 9815 22559
rect 16865 22525 16899 22559
rect 17141 22525 17175 22559
rect 19257 22525 19291 22559
rect 19533 22525 19567 22559
rect 2697 22389 2731 22423
rect 1685 22185 1719 22219
rect 13013 22185 13047 22219
rect 19625 22185 19659 22219
rect 2789 22049 2823 22083
rect 11529 22049 11563 22083
rect 13277 22049 13311 22083
rect 20269 22049 20303 22083
rect 58265 22049 58299 22083
rect 1869 21981 1903 22015
rect 18889 21981 18923 22015
rect 19993 21981 20027 22015
rect 57989 21981 58023 22015
rect 3433 21913 3467 21947
rect 18337 21913 18371 21947
rect 20085 21913 20119 21947
rect 20821 21845 20855 21879
rect 19441 21641 19475 21675
rect 58173 21641 58207 21675
rect 14749 21573 14783 21607
rect 2329 21505 2363 21539
rect 13001 21505 13035 21539
rect 19349 21505 19383 21539
rect 57529 21505 57563 21539
rect 58357 21505 58391 21539
rect 2053 21437 2087 21471
rect 2237 21437 2271 21471
rect 19625 21437 19659 21471
rect 2697 21301 2731 21335
rect 3249 21301 3283 21335
rect 12449 21301 12483 21335
rect 18521 21301 18555 21335
rect 18981 21301 19015 21335
rect 20269 21301 20303 21335
rect 1685 21097 1719 21131
rect 3985 21097 4019 21131
rect 6837 21097 6871 21131
rect 8321 21097 8355 21131
rect 14381 21097 14415 21131
rect 18705 21097 18739 21131
rect 58173 21097 58207 21131
rect 2513 21029 2547 21063
rect 5457 20961 5491 20995
rect 5733 20961 5767 20995
rect 8585 20961 8619 20995
rect 16129 20961 16163 20995
rect 1869 20893 1903 20927
rect 2329 20893 2363 20927
rect 2973 20893 3007 20927
rect 57713 20893 57747 20927
rect 58357 20893 58391 20927
rect 15853 20825 15887 20859
rect 11897 20757 11931 20791
rect 1685 20553 1719 20587
rect 2789 20553 2823 20587
rect 8309 20553 8343 20587
rect 14289 20553 14323 20587
rect 4997 20485 5031 20519
rect 12173 20485 12207 20519
rect 12357 20485 12391 20519
rect 19165 20485 19199 20519
rect 20361 20485 20395 20519
rect 1869 20417 1903 20451
rect 5181 20417 5215 20451
rect 9597 20417 9631 20451
rect 16037 20417 16071 20451
rect 18337 20417 18371 20451
rect 20637 20417 20671 20451
rect 21097 20417 21131 20451
rect 15761 20349 15795 20383
rect 19257 20349 19291 20383
rect 19441 20349 19475 20383
rect 10149 20281 10183 20315
rect 5825 20213 5859 20247
rect 17601 20213 17635 20247
rect 18153 20213 18187 20247
rect 18797 20213 18831 20247
rect 12633 19941 12667 19975
rect 2145 19873 2179 19907
rect 5549 19873 5583 19907
rect 7573 19873 7607 19907
rect 10885 19873 10919 19907
rect 11161 19873 11195 19907
rect 2329 19805 2363 19839
rect 57713 19805 57747 19839
rect 58357 19805 58391 19839
rect 2237 19737 2271 19771
rect 3157 19737 3191 19771
rect 7297 19737 7331 19771
rect 2697 19669 2731 19703
rect 18705 19669 18739 19703
rect 19717 19669 19751 19703
rect 58173 19669 58207 19703
rect 1685 19465 1719 19499
rect 10517 19465 10551 19499
rect 12725 19465 12759 19499
rect 17417 19465 17451 19499
rect 18613 19465 18647 19499
rect 58173 19465 58207 19499
rect 1869 19329 1903 19363
rect 8769 19329 8803 19363
rect 14473 19329 14507 19363
rect 17601 19329 17635 19363
rect 18981 19329 19015 19363
rect 58357 19329 58391 19363
rect 3065 19261 3099 19295
rect 9045 19261 9079 19295
rect 14197 19261 14231 19295
rect 19073 19261 19107 19295
rect 19257 19261 19291 19295
rect 19901 19261 19935 19295
rect 18153 19125 18187 19159
rect 20453 19125 20487 19159
rect 1685 18921 1719 18955
rect 2513 18921 2547 18955
rect 3065 18921 3099 18955
rect 16957 18921 16991 18955
rect 58357 18921 58391 18955
rect 18613 18785 18647 18819
rect 20085 18785 20119 18819
rect 1869 18717 1903 18751
rect 2329 18717 2363 18751
rect 17141 18717 17175 18751
rect 17969 18717 18003 18751
rect 18889 18717 18923 18751
rect 19809 18649 19843 18683
rect 17785 18581 17819 18615
rect 19441 18581 19475 18615
rect 19901 18581 19935 18615
rect 20637 18581 20671 18615
rect 1961 18377 1995 18411
rect 2421 18377 2455 18411
rect 6653 18377 6687 18411
rect 18337 18377 18371 18411
rect 18705 18377 18739 18411
rect 2053 18309 2087 18343
rect 8125 18309 8159 18343
rect 18797 18309 18831 18343
rect 20085 18309 20119 18343
rect 17509 18241 17543 18275
rect 57529 18241 57563 18275
rect 58357 18241 58391 18275
rect 1869 18173 1903 18207
rect 2881 18173 2915 18207
rect 4629 18173 4663 18207
rect 4905 18173 4939 18207
rect 8401 18173 8435 18207
rect 18981 18173 19015 18207
rect 17325 18105 17359 18139
rect 19625 18037 19659 18071
rect 58173 18037 58207 18071
rect 1685 17833 1719 17867
rect 3065 17833 3099 17867
rect 10057 17833 10091 17867
rect 18153 17833 18187 17867
rect 19533 17833 19567 17867
rect 11529 17697 11563 17731
rect 15209 17697 15243 17731
rect 18797 17697 18831 17731
rect 1869 17629 1903 17663
rect 2605 17629 2639 17663
rect 11805 17629 11839 17663
rect 17233 17629 17267 17663
rect 57713 17629 57747 17663
rect 58357 17629 58391 17663
rect 16957 17561 16991 17595
rect 2421 17493 2455 17527
rect 18521 17493 18555 17527
rect 18613 17493 18647 17527
rect 58173 17493 58207 17527
rect 2329 17289 2363 17323
rect 3801 17289 3835 17323
rect 11989 17289 12023 17323
rect 17785 17289 17819 17323
rect 19073 17289 19107 17323
rect 2237 17221 2271 17255
rect 3157 17153 3191 17187
rect 5365 17153 5399 17187
rect 13737 17153 13771 17187
rect 15945 17153 15979 17187
rect 18429 17153 18463 17187
rect 2053 17085 2087 17119
rect 5549 17085 5583 17119
rect 13461 17085 13495 17119
rect 15669 17085 15703 17119
rect 2697 17017 2731 17051
rect 3341 17017 3375 17051
rect 14197 17017 14231 17051
rect 18245 17017 18279 17051
rect 6561 16949 6595 16983
rect 3065 16745 3099 16779
rect 17785 16745 17819 16779
rect 5641 16609 5675 16643
rect 5917 16609 5951 16643
rect 1869 16541 1903 16575
rect 2421 16541 2455 16575
rect 17969 16541 18003 16575
rect 57713 16541 57747 16575
rect 58357 16541 58391 16575
rect 1685 16405 1719 16439
rect 2605 16405 2639 16439
rect 4169 16405 4203 16439
rect 58173 16405 58207 16439
rect 10425 16201 10459 16235
rect 18153 16201 18187 16235
rect 18797 16201 18831 16235
rect 8953 16133 8987 16167
rect 1869 16065 1903 16099
rect 13001 16065 13035 16099
rect 18337 16065 18371 16099
rect 19165 16065 19199 16099
rect 58357 16065 58391 16099
rect 8677 15997 8711 16031
rect 19257 15997 19291 16031
rect 19441 15997 19475 16031
rect 1685 15861 1719 15895
rect 2421 15861 2455 15895
rect 12541 15861 12575 15895
rect 14473 15861 14507 15895
rect 20085 15861 20119 15895
rect 58173 15861 58207 15895
rect 2789 15657 2823 15691
rect 5917 15657 5951 15691
rect 10885 15657 10919 15691
rect 18613 15657 18647 15691
rect 58357 15657 58391 15691
rect 2053 15589 2087 15623
rect 7389 15521 7423 15555
rect 9413 15521 9447 15555
rect 57253 15521 57287 15555
rect 7665 15453 7699 15487
rect 9137 15453 9171 15487
rect 19625 15453 19659 15487
rect 56977 15453 57011 15487
rect 19441 15317 19475 15351
rect 20085 15317 20119 15351
rect 56425 15317 56459 15351
rect 12357 15113 12391 15147
rect 19625 15113 19659 15147
rect 14841 15045 14875 15079
rect 19993 15045 20027 15079
rect 2329 14977 2363 15011
rect 9597 14977 9631 15011
rect 14565 14977 14599 15011
rect 16865 14977 16899 15011
rect 18889 14977 18923 15011
rect 57529 14977 57563 15011
rect 58357 14977 58391 15011
rect 2053 14909 2087 14943
rect 2237 14909 2271 14943
rect 13829 14909 13863 14943
rect 14105 14909 14139 14943
rect 17141 14909 17175 14943
rect 20085 14909 20119 14943
rect 20269 14909 20303 14943
rect 10149 14841 10183 14875
rect 2697 14773 2731 14807
rect 3157 14773 3191 14807
rect 3801 14773 3835 14807
rect 8309 14773 8343 14807
rect 20821 14773 20855 14807
rect 58173 14773 58207 14807
rect 1685 14569 1719 14603
rect 5089 14569 5123 14603
rect 18797 14569 18831 14603
rect 19441 14569 19475 14603
rect 20821 14569 20855 14603
rect 3249 14501 3283 14535
rect 6561 14433 6595 14467
rect 6837 14433 6871 14467
rect 9321 14433 9355 14467
rect 19901 14433 19935 14467
rect 19993 14433 20027 14467
rect 1869 14365 1903 14399
rect 2605 14365 2639 14399
rect 3065 14365 3099 14399
rect 21005 14365 21039 14399
rect 57713 14365 57747 14399
rect 58357 14365 58391 14399
rect 9597 14297 9631 14331
rect 11529 14297 11563 14331
rect 2421 14229 2455 14263
rect 4077 14229 4111 14263
rect 11069 14229 11103 14263
rect 12817 14229 12851 14263
rect 14381 14229 14415 14263
rect 19809 14229 19843 14263
rect 58173 14229 58207 14263
rect 3341 14025 3375 14059
rect 13277 14025 13311 14059
rect 20177 14025 20211 14059
rect 20729 14025 20763 14059
rect 58265 14025 58299 14059
rect 2329 13957 2363 13991
rect 3893 13957 3927 13991
rect 21189 13957 21223 13991
rect 3157 13889 3191 13923
rect 21097 13889 21131 13923
rect 2145 13821 2179 13855
rect 2237 13821 2271 13855
rect 11713 13821 11747 13855
rect 15025 13821 15059 13855
rect 21373 13821 21407 13855
rect 2697 13685 2731 13719
rect 14767 13685 14801 13719
rect 22017 13685 22051 13719
rect 2513 13481 2547 13515
rect 18429 13481 18463 13515
rect 2973 13413 3007 13447
rect 57161 13345 57195 13379
rect 57320 13345 57354 13379
rect 57437 13345 57471 13379
rect 57713 13345 57747 13379
rect 58173 13345 58207 13379
rect 1869 13277 1903 13311
rect 2329 13277 2363 13311
rect 16681 13277 16715 13311
rect 58357 13277 58391 13311
rect 16957 13209 16991 13243
rect 1685 13141 1719 13175
rect 56517 13141 56551 13175
rect 18429 12937 18463 12971
rect 19073 12937 19107 12971
rect 19533 12937 19567 12971
rect 57437 12937 57471 12971
rect 1869 12801 1903 12835
rect 18613 12801 18647 12835
rect 19441 12801 19475 12835
rect 58357 12801 58391 12835
rect 19717 12733 19751 12767
rect 2421 12665 2455 12699
rect 58173 12665 58207 12699
rect 1685 12597 1719 12631
rect 20361 12597 20395 12631
rect 9229 12393 9263 12427
rect 19441 12393 19475 12427
rect 57713 12393 57747 12427
rect 15853 12325 15887 12359
rect 10977 12257 11011 12291
rect 17601 12257 17635 12291
rect 55689 12189 55723 12223
rect 57161 12189 57195 12223
rect 58357 12189 58391 12223
rect 10701 12121 10735 12155
rect 17325 12121 17359 12155
rect 1961 12053 1995 12087
rect 8585 12053 8619 12087
rect 55505 12053 55539 12087
rect 58173 12053 58207 12087
rect 11069 11849 11103 11883
rect 19073 11849 19107 11883
rect 3065 11781 3099 11815
rect 13829 11781 13863 11815
rect 19717 11781 19751 11815
rect 1869 11713 1903 11747
rect 9321 11713 9355 11747
rect 19257 11713 19291 11747
rect 57529 11713 57563 11747
rect 58357 11713 58391 11747
rect 9597 11645 9631 11679
rect 14105 11645 14139 11679
rect 1685 11577 1719 11611
rect 3525 11577 3559 11611
rect 2421 11509 2455 11543
rect 12357 11509 12391 11543
rect 20729 11509 20763 11543
rect 58173 11509 58207 11543
rect 18705 11305 18739 11339
rect 56517 11305 56551 11339
rect 2697 11237 2731 11271
rect 3341 11237 3375 11271
rect 6745 11237 6779 11271
rect 19441 11237 19475 11271
rect 2145 11169 2179 11203
rect 5917 11169 5951 11203
rect 19901 11169 19935 11203
rect 20085 11169 20119 11203
rect 21557 11169 21591 11203
rect 57161 11169 57195 11203
rect 57320 11169 57354 11203
rect 57713 11169 57747 11203
rect 2329 11101 2363 11135
rect 3157 11101 3191 11135
rect 4169 11101 4203 11135
rect 6193 11101 6227 11135
rect 18889 11101 18923 11135
rect 19809 11101 19843 11135
rect 21373 11101 21407 11135
rect 57437 11101 57471 11135
rect 58173 11101 58207 11135
rect 58357 11101 58391 11135
rect 2237 11033 2271 11067
rect 21281 11033 21315 11067
rect 22201 11033 22235 11067
rect 20913 10965 20947 10999
rect 2697 10761 2731 10795
rect 19625 10761 19659 10795
rect 20177 10761 20211 10795
rect 56885 10761 56919 10795
rect 57529 10761 57563 10795
rect 13093 10693 13127 10727
rect 2329 10625 2363 10659
rect 3157 10625 3191 10659
rect 15117 10625 15151 10659
rect 19165 10625 19199 10659
rect 19257 10625 19291 10659
rect 20361 10625 20395 10659
rect 58357 10625 58391 10659
rect 2145 10557 2179 10591
rect 2237 10557 2271 10591
rect 5733 10557 5767 10591
rect 6009 10557 6043 10591
rect 14841 10557 14875 10591
rect 18981 10557 19015 10591
rect 3341 10489 3375 10523
rect 4261 10421 4295 10455
rect 12541 10421 12575 10455
rect 18337 10421 18371 10455
rect 58173 10421 58207 10455
rect 1685 10217 1719 10251
rect 3065 10217 3099 10251
rect 15025 10217 15059 10251
rect 18521 10217 18555 10251
rect 19717 10217 19751 10251
rect 58357 10217 58391 10251
rect 5825 10149 5859 10183
rect 57713 10149 57747 10183
rect 12265 10081 12299 10115
rect 16773 10081 16807 10115
rect 1869 10013 1903 10047
rect 7573 10013 7607 10047
rect 12081 10013 12115 10047
rect 57161 10013 57195 10047
rect 58173 10013 58207 10047
rect 7297 9945 7331 9979
rect 16497 9945 16531 9979
rect 2513 9877 2547 9911
rect 11713 9877 11747 9911
rect 12173 9877 12207 9911
rect 13001 9877 13035 9911
rect 56977 9673 57011 9707
rect 5733 9605 5767 9639
rect 14105 9605 14139 9639
rect 20821 9605 20855 9639
rect 1869 9537 1903 9571
rect 9965 9537 9999 9571
rect 19901 9537 19935 9571
rect 20913 9537 20947 9571
rect 57529 9537 57563 9571
rect 58173 9537 58207 9571
rect 2421 9469 2455 9503
rect 6009 9469 6043 9503
rect 9689 9469 9723 9503
rect 14381 9469 14415 9503
rect 21097 9469 21131 9503
rect 1685 9401 1719 9435
rect 4261 9401 4295 9435
rect 19717 9401 19751 9435
rect 20453 9401 20487 9435
rect 58357 9401 58391 9435
rect 8217 9333 8251 9367
rect 12633 9333 12667 9367
rect 1685 9129 1719 9163
rect 2789 9129 2823 9163
rect 5641 9129 5675 9163
rect 6377 9129 6411 9163
rect 12541 9129 12575 9163
rect 13185 9129 13219 9163
rect 14381 9129 14415 9163
rect 20269 9129 20303 9163
rect 10793 8993 10827 9027
rect 21649 8993 21683 9027
rect 56057 8993 56091 9027
rect 57161 8993 57195 9027
rect 57320 8993 57354 9027
rect 57437 8993 57471 9027
rect 57713 8993 57747 9027
rect 58173 8993 58207 9027
rect 1869 8925 1903 8959
rect 5825 8925 5859 8959
rect 10149 8925 10183 8959
rect 13001 8925 13035 8959
rect 21925 8925 21959 8959
rect 58357 8925 58391 8959
rect 11069 8857 11103 8891
rect 10333 8789 10367 8823
rect 21005 8789 21039 8823
rect 21833 8789 21867 8823
rect 22293 8789 22327 8823
rect 22753 8789 22787 8823
rect 56517 8789 56551 8823
rect 2697 8585 2731 8619
rect 3801 8585 3835 8619
rect 14473 8585 14507 8619
rect 57345 8585 57379 8619
rect 58357 8585 58391 8619
rect 12541 8517 12575 8551
rect 13001 8517 13035 8551
rect 56241 8517 56275 8551
rect 56609 8517 56643 8551
rect 2329 8449 2363 8483
rect 3157 8449 3191 8483
rect 22201 8449 22235 8483
rect 56977 8449 57011 8483
rect 57069 8449 57103 8483
rect 58173 8449 58207 8483
rect 2053 8381 2087 8415
rect 2237 8381 2271 8415
rect 3341 8313 3375 8347
rect 56057 8313 56091 8347
rect 22017 8245 22051 8279
rect 1685 8041 1719 8075
rect 4445 8041 4479 8075
rect 57069 8041 57103 8075
rect 57713 8041 57747 8075
rect 58173 8041 58207 8075
rect 3065 7973 3099 8007
rect 5917 7905 5951 7939
rect 15853 7905 15887 7939
rect 17601 7905 17635 7939
rect 22569 7905 22603 7939
rect 1869 7837 1903 7871
rect 2605 7837 2639 7871
rect 6193 7837 6227 7871
rect 17877 7837 17911 7871
rect 21741 7837 21775 7871
rect 22293 7837 22327 7871
rect 22661 7837 22695 7871
rect 58357 7837 58391 7871
rect 21189 7769 21223 7803
rect 2421 7701 2455 7735
rect 2421 7497 2455 7531
rect 2789 7497 2823 7531
rect 3893 7497 3927 7531
rect 8309 7497 8343 7531
rect 13829 7497 13863 7531
rect 19441 7497 19475 7531
rect 57529 7497 57563 7531
rect 15301 7429 15335 7463
rect 22661 7429 22695 7463
rect 58265 7429 58299 7463
rect 3249 7361 3283 7395
rect 9597 7361 9631 7395
rect 10057 7361 10091 7395
rect 15577 7361 15611 7395
rect 19625 7361 19659 7395
rect 21465 7361 21499 7395
rect 22201 7361 22235 7395
rect 22845 7361 22879 7395
rect 23581 7361 23615 7395
rect 2145 7293 2179 7327
rect 2329 7293 2363 7327
rect 3433 7157 3467 7191
rect 56977 7157 57011 7191
rect 8321 6953 8355 6987
rect 22477 6953 22511 6987
rect 57713 6953 57747 6987
rect 2237 6817 2271 6851
rect 6837 6817 6871 6851
rect 20637 6817 20671 6851
rect 57069 6817 57103 6851
rect 8585 6749 8619 6783
rect 19717 6749 19751 6783
rect 20913 6749 20947 6783
rect 22017 6749 22051 6783
rect 22937 6749 22971 6783
rect 55689 6749 55723 6783
rect 56241 6749 56275 6783
rect 56609 6749 56643 6783
rect 58357 6749 58391 6783
rect 2421 6681 2455 6715
rect 2329 6613 2363 6647
rect 2789 6613 2823 6647
rect 3341 6613 3375 6647
rect 19533 6613 19567 6647
rect 21557 6613 21591 6647
rect 58173 6613 58207 6647
rect 1685 6409 1719 6443
rect 4261 6409 4295 6443
rect 19257 6409 19291 6443
rect 19717 6409 19751 6443
rect 9597 6341 9631 6375
rect 10057 6341 10091 6375
rect 13461 6341 13495 6375
rect 18705 6341 18739 6375
rect 20177 6341 20211 6375
rect 1869 6273 1903 6307
rect 2605 6273 2639 6307
rect 13185 6273 13219 6307
rect 20085 6273 20119 6307
rect 55689 6273 55723 6307
rect 56726 6273 56760 6307
rect 56885 6273 56919 6307
rect 58357 6273 58391 6307
rect 5733 6205 5767 6239
rect 6009 6205 6043 6239
rect 12725 6205 12759 6239
rect 14933 6205 14967 6239
rect 20361 6205 20395 6239
rect 20913 6205 20947 6239
rect 55873 6205 55907 6239
rect 56609 6205 56643 6239
rect 2789 6137 2823 6171
rect 56333 6137 56367 6171
rect 3249 6069 3283 6103
rect 8309 6069 8343 6103
rect 22109 6069 22143 6103
rect 57529 6069 57563 6103
rect 58173 6069 58207 6103
rect 1685 5865 1719 5899
rect 12081 5865 12115 5899
rect 18797 5865 18831 5899
rect 19717 5865 19751 5899
rect 57161 5797 57195 5831
rect 9781 5729 9815 5763
rect 11529 5729 11563 5763
rect 20177 5729 20211 5763
rect 20361 5729 20395 5763
rect 56517 5729 56551 5763
rect 57437 5729 57471 5763
rect 57575 5729 57609 5763
rect 1869 5661 1903 5695
rect 9505 5661 9539 5695
rect 20085 5661 20119 5695
rect 56701 5661 56735 5695
rect 57713 5661 57747 5695
rect 56057 5525 56091 5559
rect 58357 5525 58391 5559
rect 12541 5321 12575 5355
rect 19625 5321 19659 5355
rect 56977 5321 57011 5355
rect 57529 5321 57563 5355
rect 58173 5321 58207 5355
rect 10057 5253 10091 5287
rect 13001 5253 13035 5287
rect 1869 5185 1903 5219
rect 56425 5185 56459 5219
rect 58357 5185 58391 5219
rect 10333 5117 10367 5151
rect 14749 5117 14783 5151
rect 1685 5049 1719 5083
rect 8585 4981 8619 5015
rect 5917 4777 5951 4811
rect 21649 4777 21683 4811
rect 57713 4777 57747 4811
rect 58173 4777 58207 4811
rect 19441 4709 19475 4743
rect 6469 4641 6503 4675
rect 8217 4641 8251 4675
rect 8493 4641 8527 4675
rect 16865 4641 16899 4675
rect 17141 4641 17175 4675
rect 18889 4641 18923 4675
rect 22661 4641 22695 4675
rect 22753 4641 22787 4675
rect 1869 4573 1903 4607
rect 57069 4573 57103 4607
rect 57529 4573 57563 4607
rect 58357 4573 58391 4607
rect 56517 4505 56551 4539
rect 1685 4437 1719 4471
rect 2789 4437 2823 4471
rect 15577 4437 15611 4471
rect 20085 4437 20119 4471
rect 22201 4437 22235 4471
rect 22569 4437 22603 4471
rect 55965 4437 55999 4471
rect 18613 4233 18647 4267
rect 19625 4233 19659 4267
rect 2329 4165 2363 4199
rect 5457 4165 5491 4199
rect 16037 4165 16071 4199
rect 16313 4097 16347 4131
rect 18797 4097 18831 4131
rect 21465 4097 21499 4131
rect 22385 4097 22419 4131
rect 23029 4097 23063 4131
rect 55873 4097 55907 4131
rect 56609 4097 56643 4131
rect 57529 4097 57563 4131
rect 58265 4097 58299 4131
rect 2145 4029 2179 4063
rect 2237 4029 2271 4063
rect 5733 4029 5767 4063
rect 14565 4029 14599 4063
rect 19717 4029 19751 4063
rect 19809 4029 19843 4063
rect 22845 3961 22879 3995
rect 57345 3961 57379 3995
rect 2697 3893 2731 3927
rect 3249 3893 3283 3927
rect 12265 3893 12299 3927
rect 16865 3893 16899 3927
rect 18061 3893 18095 3927
rect 19257 3893 19291 3927
rect 20453 3893 20487 3927
rect 22201 3893 22235 3927
rect 55321 3893 55355 3927
rect 58081 3893 58115 3927
rect 3341 3689 3375 3723
rect 5653 3689 5687 3723
rect 11161 3689 11195 3723
rect 13369 3689 13403 3723
rect 18889 3689 18923 3723
rect 22753 3689 22787 3723
rect 4169 3621 4203 3655
rect 14749 3621 14783 3655
rect 40141 3621 40175 3655
rect 2145 3553 2179 3587
rect 2237 3553 2271 3587
rect 12633 3553 12667 3587
rect 12909 3553 12943 3587
rect 16497 3553 16531 3587
rect 18337 3553 18371 3587
rect 20913 3553 20947 3587
rect 22109 3553 22143 3587
rect 22293 3553 22327 3587
rect 3157 3485 3191 3519
rect 5917 3485 5951 3519
rect 6837 3485 6871 3519
rect 17693 3485 17727 3519
rect 18521 3485 18555 3519
rect 19901 3485 19935 3519
rect 20729 3485 20763 3519
rect 22385 3485 22419 3519
rect 23213 3485 23247 3519
rect 39129 3485 39163 3519
rect 46489 3485 46523 3519
rect 48513 3485 48547 3519
rect 48973 3485 49007 3519
rect 53113 3485 53147 3519
rect 53573 3485 53607 3519
rect 54585 3485 54619 3519
rect 55689 3485 55723 3519
rect 56517 3485 56551 3519
rect 57161 3485 57195 3519
rect 57621 3485 57655 3519
rect 2329 3417 2363 3451
rect 6469 3417 6503 3451
rect 16221 3417 16255 3451
rect 47041 3417 47075 3451
rect 2697 3349 2731 3383
rect 7297 3349 7331 3383
rect 9137 3349 9171 3383
rect 17049 3349 17083 3383
rect 18429 3349 18463 3383
rect 19717 3349 19751 3383
rect 20361 3349 20395 3383
rect 20821 3349 20855 3383
rect 23397 3349 23431 3383
rect 38945 3349 38979 3383
rect 46305 3349 46339 3383
rect 48329 3349 48363 3383
rect 52929 3349 52963 3383
rect 54401 3349 54435 3383
rect 55505 3349 55539 3383
rect 56333 3349 56367 3383
rect 56977 3349 57011 3383
rect 57805 3349 57839 3383
rect 58357 3349 58391 3383
rect 4077 3145 4111 3179
rect 6561 3145 6595 3179
rect 8033 3145 8067 3179
rect 11713 3145 11747 3179
rect 19165 3145 19199 3179
rect 22569 3145 22603 3179
rect 27261 3145 27295 3179
rect 28733 3145 28767 3179
rect 29837 3145 29871 3179
rect 30941 3145 30975 3179
rect 33149 3145 33183 3179
rect 42993 3145 43027 3179
rect 43729 3145 43763 3179
rect 44833 3145 44867 3179
rect 51457 3145 51491 3179
rect 54677 3145 54711 3179
rect 55873 3145 55907 3179
rect 56517 3145 56551 3179
rect 3525 3077 3559 3111
rect 9505 3077 9539 3111
rect 12265 3077 12299 3111
rect 12633 3077 12667 3111
rect 15393 3077 15427 3111
rect 21373 3077 21407 3111
rect 32321 3077 32355 3111
rect 37933 3077 37967 3111
rect 2237 3009 2271 3043
rect 2973 3009 3007 3043
rect 5825 3009 5859 3043
rect 9781 3009 9815 3043
rect 15669 3009 15703 3043
rect 18153 3009 18187 3043
rect 19349 3009 19383 3043
rect 20085 3009 20119 3043
rect 20361 3009 20395 3043
rect 22201 3009 22235 3043
rect 22385 3009 22419 3043
rect 23029 3009 23063 3043
rect 27813 3009 27847 3043
rect 55413 3009 55447 3043
rect 56057 3009 56091 3043
rect 56701 3009 56735 3043
rect 57345 3009 57379 3043
rect 58265 3009 58299 3043
rect 5549 2941 5583 2975
rect 16313 2941 16347 2975
rect 17877 2941 17911 2975
rect 40509 2941 40543 2975
rect 50813 2941 50847 2975
rect 2421 2873 2455 2907
rect 13921 2873 13955 2907
rect 38669 2873 38703 2907
rect 58081 2873 58115 2907
rect 7481 2805 7515 2839
rect 10241 2805 10275 2839
rect 11161 2805 11195 2839
rect 13461 2805 13495 2839
rect 17417 2805 17451 2839
rect 23857 2805 23891 2839
rect 24409 2805 24443 2839
rect 25513 2805 25547 2839
rect 27997 2805 28031 2839
rect 36001 2805 36035 2839
rect 54217 2805 54251 2839
rect 57161 2805 57195 2839
rect 2605 2601 2639 2635
rect 4813 2601 4847 2635
rect 14657 2601 14691 2635
rect 15853 2601 15887 2635
rect 22477 2601 22511 2635
rect 24961 2601 24995 2635
rect 56701 2601 56735 2635
rect 6837 2533 6871 2567
rect 17141 2533 17175 2567
rect 25789 2533 25823 2567
rect 57345 2533 57379 2567
rect 9413 2465 9447 2499
rect 18889 2465 18923 2499
rect 19625 2465 19659 2499
rect 20637 2465 20671 2499
rect 23489 2465 23523 2499
rect 27997 2465 28031 2499
rect 36369 2465 36403 2499
rect 1961 2397 1995 2431
rect 2421 2397 2455 2431
rect 3433 2397 3467 2431
rect 4629 2397 4663 2431
rect 5733 2397 5767 2431
rect 7021 2397 7055 2431
rect 10149 2397 10183 2431
rect 12357 2397 12391 2431
rect 12541 2397 12575 2431
rect 13461 2397 13495 2431
rect 14749 2397 14783 2431
rect 15761 2397 15795 2431
rect 18613 2397 18647 2431
rect 20913 2397 20947 2431
rect 22293 2397 22327 2431
rect 23213 2397 23247 2431
rect 25605 2397 25639 2431
rect 28917 2397 28951 2431
rect 30021 2397 30055 2431
rect 31125 2397 31159 2431
rect 32321 2397 32355 2431
rect 33333 2397 33367 2431
rect 34989 2397 35023 2431
rect 36093 2397 36127 2431
rect 37749 2397 37783 2431
rect 38485 2397 38519 2431
rect 38945 2397 38979 2431
rect 40325 2397 40359 2431
rect 41337 2397 41371 2431
rect 42901 2397 42935 2431
rect 43637 2397 43671 2431
rect 44649 2397 44683 2431
rect 45753 2397 45787 2431
rect 46857 2397 46891 2431
rect 48053 2397 48087 2431
rect 49065 2397 49099 2431
rect 49525 2397 49559 2431
rect 50629 2397 50663 2431
rect 51365 2397 51399 2431
rect 52377 2397 52411 2431
rect 53481 2397 53515 2431
rect 54585 2397 54619 2431
rect 55781 2397 55815 2431
rect 56517 2397 56551 2431
rect 57529 2397 57563 2431
rect 58081 2397 58115 2431
rect 4169 2329 4203 2363
rect 8033 2329 8067 2363
rect 9229 2329 9263 2363
rect 10333 2329 10367 2363
rect 11069 2329 11103 2363
rect 16957 2329 16991 2363
rect 20177 2329 20211 2363
rect 24685 2329 24719 2363
rect 27169 2329 27203 2363
rect 35541 2329 35575 2363
rect 5917 2261 5951 2295
rect 8125 2261 8159 2295
rect 10977 2261 11011 2295
rect 11897 2261 11931 2295
rect 13645 2261 13679 2295
rect 26617 2261 26651 2295
rect 29101 2261 29135 2295
rect 30205 2261 30239 2295
rect 31309 2261 31343 2295
rect 32505 2261 32539 2295
rect 33517 2261 33551 2295
rect 34345 2261 34379 2295
rect 37565 2261 37599 2295
rect 38301 2261 38335 2295
rect 39129 2261 39163 2295
rect 40141 2261 40175 2295
rect 41153 2261 41187 2295
rect 41889 2261 41923 2295
rect 42717 2261 42751 2295
rect 43453 2261 43487 2295
rect 44465 2261 44499 2295
rect 45569 2261 45603 2295
rect 46673 2261 46707 2295
rect 47869 2261 47903 2295
rect 48881 2261 48915 2295
rect 50445 2261 50479 2295
rect 51181 2261 51215 2295
rect 52193 2261 52227 2295
rect 53297 2261 53331 2295
rect 54401 2261 54435 2295
rect 55597 2261 55631 2295
rect 58265 2261 58299 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 2133 57579 2191 57585
rect 2133 57545 2145 57579
rect 2179 57576 2191 57579
rect 11149 57579 11207 57585
rect 2179 57548 6914 57576
rect 2179 57545 2191 57548
rect 2133 57539 2191 57545
rect 6886 57508 6914 57548
rect 11149 57545 11161 57579
rect 11195 57576 11207 57579
rect 11422 57576 11428 57588
rect 11195 57548 11428 57576
rect 11195 57545 11207 57548
rect 11149 57539 11207 57545
rect 11422 57536 11428 57548
rect 11480 57536 11486 57588
rect 13725 57579 13783 57585
rect 13725 57545 13737 57579
rect 13771 57576 13783 57579
rect 13814 57576 13820 57588
rect 13771 57548 13820 57576
rect 13771 57545 13783 57548
rect 13725 57539 13783 57545
rect 13814 57536 13820 57548
rect 13872 57536 13878 57588
rect 16206 57576 16212 57588
rect 16167 57548 16212 57576
rect 16206 57536 16212 57548
rect 16264 57536 16270 57588
rect 17037 57579 17095 57585
rect 17037 57545 17049 57579
rect 17083 57576 17095 57579
rect 20714 57576 20720 57588
rect 17083 57548 20720 57576
rect 17083 57545 17095 57548
rect 17037 57539 17095 57545
rect 20714 57536 20720 57548
rect 20772 57536 20778 57588
rect 22465 57579 22523 57585
rect 22465 57545 22477 57579
rect 22511 57545 22523 57579
rect 22465 57539 22523 57545
rect 25409 57579 25467 57585
rect 25409 57545 25421 57579
rect 25455 57576 25467 57579
rect 25774 57576 25780 57588
rect 25455 57548 25780 57576
rect 25455 57545 25467 57548
rect 25409 57539 25467 57545
rect 20898 57508 20904 57520
rect 6886 57480 20904 57508
rect 20898 57468 20904 57480
rect 20956 57468 20962 57520
rect 22480 57508 22508 57539
rect 25774 57536 25780 57548
rect 25832 57536 25838 57588
rect 26605 57579 26663 57585
rect 26605 57545 26617 57579
rect 26651 57576 26663 57579
rect 26970 57576 26976 57588
rect 26651 57548 26976 57576
rect 26651 57545 26663 57548
rect 26605 57539 26663 57545
rect 26970 57536 26976 57548
rect 27028 57536 27034 57588
rect 29181 57579 29239 57585
rect 29181 57545 29193 57579
rect 29227 57576 29239 57579
rect 29362 57576 29368 57588
rect 29227 57548 29368 57576
rect 29227 57545 29239 57548
rect 29181 57539 29239 57545
rect 29362 57536 29368 57548
rect 29420 57536 29426 57588
rect 34146 57536 34152 57588
rect 34204 57576 34210 57588
rect 34241 57579 34299 57585
rect 34241 57576 34253 57579
rect 34204 57548 34253 57576
rect 34204 57536 34210 57548
rect 34241 57545 34253 57548
rect 34287 57545 34299 57579
rect 34241 57539 34299 57545
rect 22480 57480 25728 57508
rect 1854 57400 1860 57452
rect 1912 57440 1918 57452
rect 1949 57443 2007 57449
rect 1949 57440 1961 57443
rect 1912 57412 1961 57440
rect 1912 57400 1918 57412
rect 1949 57409 1961 57412
rect 1995 57409 2007 57443
rect 1949 57403 2007 57409
rect 3050 57400 3056 57452
rect 3108 57440 3114 57452
rect 3421 57443 3479 57449
rect 3421 57440 3433 57443
rect 3108 57412 3433 57440
rect 3108 57400 3114 57412
rect 3421 57409 3433 57412
rect 3467 57409 3479 57443
rect 3421 57403 3479 57409
rect 4246 57400 4252 57452
rect 4304 57440 4310 57452
rect 4341 57443 4399 57449
rect 4341 57440 4353 57443
rect 4304 57412 4353 57440
rect 4304 57400 4310 57412
rect 4341 57409 4353 57412
rect 4387 57440 4399 57443
rect 4614 57440 4620 57452
rect 4387 57412 4620 57440
rect 4387 57409 4399 57412
rect 4341 57403 4399 57409
rect 4614 57400 4620 57412
rect 4672 57400 4678 57452
rect 5534 57400 5540 57452
rect 5592 57440 5598 57452
rect 5997 57443 6055 57449
rect 5997 57440 6009 57443
rect 5592 57412 6009 57440
rect 5592 57400 5598 57412
rect 5997 57409 6009 57412
rect 6043 57440 6055 57443
rect 6549 57443 6607 57449
rect 6549 57440 6561 57443
rect 6043 57412 6561 57440
rect 6043 57409 6055 57412
rect 5997 57403 6055 57409
rect 6549 57409 6561 57412
rect 6595 57409 6607 57443
rect 6549 57403 6607 57409
rect 7834 57400 7840 57452
rect 7892 57440 7898 57452
rect 8478 57440 8484 57452
rect 7892 57412 8484 57440
rect 7892 57400 7898 57412
rect 8478 57400 8484 57412
rect 8536 57440 8542 57452
rect 8573 57443 8631 57449
rect 8573 57440 8585 57443
rect 8536 57412 8585 57440
rect 8536 57400 8542 57412
rect 8573 57409 8585 57412
rect 8619 57409 8631 57443
rect 8573 57403 8631 57409
rect 9030 57400 9036 57452
rect 9088 57440 9094 57452
rect 9125 57443 9183 57449
rect 9125 57440 9137 57443
rect 9088 57412 9137 57440
rect 9088 57400 9094 57412
rect 9125 57409 9137 57412
rect 9171 57409 9183 57443
rect 9125 57403 9183 57409
rect 9861 57443 9919 57449
rect 9861 57409 9873 57443
rect 9907 57440 9919 57443
rect 10226 57440 10232 57452
rect 9907 57412 10232 57440
rect 9907 57409 9919 57412
rect 9861 57403 9919 57409
rect 10226 57400 10232 57412
rect 10284 57440 10290 57452
rect 10321 57443 10379 57449
rect 10321 57440 10333 57443
rect 10284 57412 10333 57440
rect 10284 57400 10290 57412
rect 10321 57409 10333 57412
rect 10367 57409 10379 57443
rect 10321 57403 10379 57409
rect 11422 57400 11428 57452
rect 11480 57440 11486 57452
rect 11701 57443 11759 57449
rect 11701 57440 11713 57443
rect 11480 57412 11713 57440
rect 11480 57400 11486 57412
rect 11701 57409 11713 57412
rect 11747 57409 11759 57443
rect 11701 57403 11759 57409
rect 12618 57400 12624 57452
rect 12676 57440 12682 57452
rect 12713 57443 12771 57449
rect 12713 57440 12725 57443
rect 12676 57412 12725 57440
rect 12676 57400 12682 57412
rect 12713 57409 12725 57412
rect 12759 57409 12771 57443
rect 12713 57403 12771 57409
rect 13814 57400 13820 57452
rect 13872 57440 13878 57452
rect 14277 57443 14335 57449
rect 14277 57440 14289 57443
rect 13872 57412 14289 57440
rect 13872 57400 13878 57412
rect 14277 57409 14289 57412
rect 14323 57409 14335 57443
rect 14277 57403 14335 57409
rect 15010 57400 15016 57452
rect 15068 57440 15074 57452
rect 15105 57443 15163 57449
rect 15105 57440 15117 57443
rect 15068 57412 15117 57440
rect 15068 57400 15074 57412
rect 15105 57409 15117 57412
rect 15151 57409 15163 57443
rect 15105 57403 15163 57409
rect 16206 57400 16212 57452
rect 16264 57440 16270 57452
rect 16853 57443 16911 57449
rect 16853 57440 16865 57443
rect 16264 57412 16865 57440
rect 16264 57400 16270 57412
rect 16853 57409 16865 57412
rect 16899 57409 16911 57443
rect 16853 57403 16911 57409
rect 17402 57400 17408 57452
rect 17460 57440 17466 57452
rect 17497 57443 17555 57449
rect 17497 57440 17509 57443
rect 17460 57412 17509 57440
rect 17460 57400 17466 57412
rect 17497 57409 17509 57412
rect 17543 57409 17555 57443
rect 17497 57403 17555 57409
rect 18233 57443 18291 57449
rect 18233 57409 18245 57443
rect 18279 57440 18291 57443
rect 18598 57440 18604 57452
rect 18279 57412 18604 57440
rect 18279 57409 18291 57412
rect 18233 57403 18291 57409
rect 18598 57400 18604 57412
rect 18656 57440 18662 57452
rect 18693 57443 18751 57449
rect 18693 57440 18705 57443
rect 18656 57412 18705 57440
rect 18656 57400 18662 57412
rect 18693 57409 18705 57412
rect 18739 57409 18751 57443
rect 18693 57403 18751 57409
rect 19889 57443 19947 57449
rect 19889 57409 19901 57443
rect 19935 57440 19947 57443
rect 19978 57440 19984 57452
rect 19935 57412 19984 57440
rect 19935 57409 19947 57412
rect 19889 57403 19947 57409
rect 19978 57400 19984 57412
rect 20036 57400 20042 57452
rect 20625 57443 20683 57449
rect 20625 57409 20637 57443
rect 20671 57440 20683 57443
rect 20990 57440 20996 57452
rect 20671 57412 20996 57440
rect 20671 57409 20683 57412
rect 20625 57403 20683 57409
rect 20990 57400 20996 57412
rect 21048 57440 21054 57452
rect 21085 57443 21143 57449
rect 21085 57440 21097 57443
rect 21048 57412 21097 57440
rect 21048 57400 21054 57412
rect 21085 57409 21097 57412
rect 21131 57409 21143 57443
rect 21085 57403 21143 57409
rect 22186 57400 22192 57452
rect 22244 57440 22250 57452
rect 22281 57443 22339 57449
rect 22281 57440 22293 57443
rect 22244 57412 22293 57440
rect 22244 57400 22250 57412
rect 22281 57409 22293 57412
rect 22327 57409 22339 57443
rect 22281 57403 22339 57409
rect 23017 57443 23075 57449
rect 23017 57409 23029 57443
rect 23063 57440 23075 57443
rect 23382 57440 23388 57452
rect 23063 57412 23388 57440
rect 23063 57409 23075 57412
rect 23017 57403 23075 57409
rect 23382 57400 23388 57412
rect 23440 57440 23446 57452
rect 23477 57443 23535 57449
rect 23477 57440 23489 57443
rect 23440 57412 23489 57440
rect 23440 57400 23446 57412
rect 23477 57409 23489 57412
rect 23523 57409 23535 57443
rect 23477 57403 23535 57409
rect 24578 57400 24584 57452
rect 24636 57440 24642 57452
rect 24673 57443 24731 57449
rect 24673 57440 24685 57443
rect 24636 57412 24685 57440
rect 24636 57400 24642 57412
rect 24673 57409 24685 57412
rect 24719 57409 24731 57443
rect 24673 57403 24731 57409
rect 3142 57372 3148 57384
rect 3103 57344 3148 57372
rect 3142 57332 3148 57344
rect 3200 57332 3206 57384
rect 5718 57372 5724 57384
rect 5679 57344 5724 57372
rect 5718 57332 5724 57344
rect 5776 57332 5782 57384
rect 8294 57372 8300 57384
rect 8255 57344 8300 57372
rect 8294 57332 8300 57344
rect 8352 57332 8358 57384
rect 20530 57372 20536 57384
rect 15304 57344 20536 57372
rect 15304 57313 15332 57344
rect 20530 57332 20536 57344
rect 20588 57332 20594 57384
rect 24946 57372 24952 57384
rect 22066 57344 24952 57372
rect 15289 57307 15347 57313
rect 15289 57273 15301 57307
rect 15335 57273 15347 57307
rect 15289 57267 15347 57273
rect 17681 57307 17739 57313
rect 17681 57273 17693 57307
rect 17727 57304 17739 57307
rect 22066 57304 22094 57344
rect 24946 57332 24952 57344
rect 25004 57332 25010 57384
rect 25700 57372 25728 57480
rect 25792 57440 25820 57536
rect 26053 57443 26111 57449
rect 26053 57440 26065 57443
rect 25792 57412 26065 57440
rect 26053 57409 26065 57412
rect 26099 57409 26111 57443
rect 26988 57440 27016 57536
rect 27341 57443 27399 57449
rect 27341 57440 27353 57443
rect 26988 57412 27353 57440
rect 26053 57403 26111 57409
rect 27341 57409 27353 57412
rect 27387 57409 27399 57443
rect 27341 57403 27399 57409
rect 28166 57400 28172 57452
rect 28224 57440 28230 57452
rect 28261 57443 28319 57449
rect 28261 57440 28273 57443
rect 28224 57412 28273 57440
rect 28224 57400 28230 57412
rect 28261 57409 28273 57412
rect 28307 57409 28319 57443
rect 29380 57440 29408 57536
rect 29917 57443 29975 57449
rect 29917 57440 29929 57443
rect 29380 57412 29929 57440
rect 28261 57403 28319 57409
rect 29917 57409 29929 57412
rect 29963 57409 29975 57443
rect 29917 57403 29975 57409
rect 30558 57400 30564 57452
rect 30616 57440 30622 57452
rect 30653 57443 30711 57449
rect 30653 57440 30665 57443
rect 30616 57412 30665 57440
rect 30616 57400 30622 57412
rect 30653 57409 30665 57412
rect 30699 57440 30711 57443
rect 31297 57443 31355 57449
rect 31297 57440 31309 57443
rect 30699 57412 31309 57440
rect 30699 57409 30711 57412
rect 30653 57403 30711 57409
rect 31297 57409 31309 57412
rect 31343 57409 31355 57443
rect 31297 57403 31355 57409
rect 31754 57400 31760 57452
rect 31812 57440 31818 57452
rect 32122 57440 32128 57452
rect 31812 57412 32128 57440
rect 31812 57400 31818 57412
rect 32122 57400 32128 57412
rect 32180 57440 32186 57452
rect 32309 57443 32367 57449
rect 32309 57440 32321 57443
rect 32180 57412 32321 57440
rect 32180 57400 32186 57412
rect 32309 57409 32321 57412
rect 32355 57409 32367 57443
rect 32309 57403 32367 57409
rect 32950 57400 32956 57452
rect 33008 57440 33014 57452
rect 33045 57443 33103 57449
rect 33045 57440 33057 57443
rect 33008 57412 33057 57440
rect 33008 57400 33014 57412
rect 33045 57409 33057 57412
rect 33091 57440 33103 57443
rect 33689 57443 33747 57449
rect 33689 57440 33701 57443
rect 33091 57412 33701 57440
rect 33091 57409 33103 57412
rect 33045 57403 33103 57409
rect 33689 57409 33701 57412
rect 33735 57409 33747 57443
rect 34256 57440 34284 57539
rect 38746 57536 38752 57588
rect 38804 57576 38810 57588
rect 41417 57579 41475 57585
rect 41417 57576 41429 57579
rect 38804 57548 41429 57576
rect 38804 57536 38810 57548
rect 41417 57545 41429 57548
rect 41463 57545 41475 57579
rect 41417 57539 41475 57545
rect 42613 57579 42671 57585
rect 42613 57545 42625 57579
rect 42659 57545 42671 57579
rect 42613 57539 42671 57545
rect 38838 57468 38844 57520
rect 38896 57508 38902 57520
rect 42628 57508 42656 57539
rect 42702 57536 42708 57588
rect 42760 57576 42766 57588
rect 46201 57579 46259 57585
rect 46201 57576 46213 57579
rect 42760 57548 46213 57576
rect 42760 57536 42766 57548
rect 46201 57545 46213 57548
rect 46247 57545 46259 57579
rect 46201 57539 46259 57545
rect 38896 57480 42656 57508
rect 38896 57468 38902 57480
rect 35069 57443 35127 57449
rect 35069 57440 35081 57443
rect 34256 57412 35081 57440
rect 33689 57403 33747 57409
rect 35069 57409 35081 57412
rect 35115 57409 35127 57443
rect 35069 57403 35127 57409
rect 35342 57400 35348 57452
rect 35400 57440 35406 57452
rect 35529 57443 35587 57449
rect 35529 57440 35541 57443
rect 35400 57412 35541 57440
rect 35400 57400 35406 57412
rect 35529 57409 35541 57412
rect 35575 57409 35587 57443
rect 35529 57403 35587 57409
rect 36538 57400 36544 57452
rect 36596 57440 36602 57452
rect 36817 57443 36875 57449
rect 36817 57440 36829 57443
rect 36596 57412 36829 57440
rect 36596 57400 36602 57412
rect 36817 57409 36829 57412
rect 36863 57409 36875 57443
rect 36817 57403 36875 57409
rect 37734 57400 37740 57452
rect 37792 57440 37798 57452
rect 38013 57443 38071 57449
rect 38013 57440 38025 57443
rect 37792 57412 38025 57440
rect 37792 57400 37798 57412
rect 38013 57409 38025 57412
rect 38059 57440 38071 57443
rect 38473 57443 38531 57449
rect 38473 57440 38485 57443
rect 38059 57412 38485 57440
rect 38059 57409 38071 57412
rect 38013 57403 38071 57409
rect 38473 57409 38485 57412
rect 38519 57409 38531 57443
rect 38473 57403 38531 57409
rect 38930 57400 38936 57452
rect 38988 57440 38994 57452
rect 39209 57443 39267 57449
rect 39209 57440 39221 57443
rect 38988 57412 39221 57440
rect 38988 57400 38994 57412
rect 39209 57409 39221 57412
rect 39255 57409 39267 57443
rect 39209 57403 39267 57409
rect 40126 57400 40132 57452
rect 40184 57440 40190 57452
rect 40405 57443 40463 57449
rect 40405 57440 40417 57443
rect 40184 57412 40417 57440
rect 40184 57400 40190 57412
rect 40405 57409 40417 57412
rect 40451 57440 40463 57443
rect 40865 57443 40923 57449
rect 40865 57440 40877 57443
rect 40451 57412 40877 57440
rect 40451 57409 40463 57412
rect 40405 57403 40463 57409
rect 40865 57409 40877 57412
rect 40911 57409 40923 57443
rect 40865 57403 40923 57409
rect 41322 57400 41328 57452
rect 41380 57440 41386 57452
rect 41601 57443 41659 57449
rect 41601 57440 41613 57443
rect 41380 57412 41613 57440
rect 41380 57400 41386 57412
rect 41601 57409 41613 57412
rect 41647 57409 41659 57443
rect 42794 57440 42800 57452
rect 42755 57412 42800 57440
rect 41601 57403 41659 57409
rect 42794 57400 42800 57412
rect 42852 57440 42858 57452
rect 43257 57443 43315 57449
rect 43257 57440 43269 57443
rect 42852 57412 43269 57440
rect 42852 57400 42858 57412
rect 43257 57409 43269 57412
rect 43303 57409 43315 57443
rect 43257 57403 43315 57409
rect 43714 57400 43720 57452
rect 43772 57440 43778 57452
rect 43993 57443 44051 57449
rect 43993 57440 44005 57443
rect 43772 57412 44005 57440
rect 43772 57400 43778 57412
rect 43993 57409 44005 57412
rect 44039 57440 44051 57443
rect 44453 57443 44511 57449
rect 44453 57440 44465 57443
rect 44039 57412 44465 57440
rect 44039 57409 44051 57412
rect 43993 57403 44051 57409
rect 44453 57409 44465 57412
rect 44499 57409 44511 57443
rect 44453 57403 44511 57409
rect 44910 57400 44916 57452
rect 44968 57440 44974 57452
rect 45373 57443 45431 57449
rect 45373 57440 45385 57443
rect 44968 57412 45385 57440
rect 44968 57400 44974 57412
rect 45373 57409 45385 57412
rect 45419 57409 45431 57443
rect 45373 57403 45431 57409
rect 46106 57400 46112 57452
rect 46164 57440 46170 57452
rect 46385 57443 46443 57449
rect 46385 57440 46397 57443
rect 46164 57412 46397 57440
rect 46164 57400 46170 57412
rect 46385 57409 46397 57412
rect 46431 57440 46443 57443
rect 46845 57443 46903 57449
rect 46845 57440 46857 57443
rect 46431 57412 46857 57440
rect 46431 57409 46443 57412
rect 46385 57403 46443 57409
rect 46845 57409 46857 57412
rect 46891 57409 46903 57443
rect 46845 57403 46903 57409
rect 47302 57400 47308 57452
rect 47360 57440 47366 57452
rect 47949 57443 48007 57449
rect 47949 57440 47961 57443
rect 47360 57412 47961 57440
rect 47360 57400 47366 57412
rect 47949 57409 47961 57412
rect 47995 57409 48007 57443
rect 47949 57403 48007 57409
rect 48498 57400 48504 57452
rect 48556 57440 48562 57452
rect 48777 57443 48835 57449
rect 48777 57440 48789 57443
rect 48556 57412 48789 57440
rect 48556 57400 48562 57412
rect 48777 57409 48789 57412
rect 48823 57440 48835 57443
rect 49237 57443 49295 57449
rect 49237 57440 49249 57443
rect 48823 57412 49249 57440
rect 48823 57409 48835 57412
rect 48777 57403 48835 57409
rect 49237 57409 49249 57412
rect 49283 57409 49295 57443
rect 49237 57403 49295 57409
rect 49694 57400 49700 57452
rect 49752 57440 49758 57452
rect 50338 57440 50344 57452
rect 49752 57412 50344 57440
rect 49752 57400 49758 57412
rect 50338 57400 50344 57412
rect 50396 57440 50402 57452
rect 50525 57443 50583 57449
rect 50525 57440 50537 57443
rect 50396 57412 50537 57440
rect 50396 57400 50402 57412
rect 50525 57409 50537 57412
rect 50571 57409 50583 57443
rect 50525 57403 50583 57409
rect 51074 57400 51080 57452
rect 51132 57440 51138 57452
rect 51169 57443 51227 57449
rect 51169 57440 51181 57443
rect 51132 57412 51181 57440
rect 51132 57400 51138 57412
rect 51169 57409 51181 57412
rect 51215 57440 51227 57443
rect 51629 57443 51687 57449
rect 51629 57440 51641 57443
rect 51215 57412 51641 57440
rect 51215 57409 51227 57412
rect 51169 57403 51227 57409
rect 51629 57409 51641 57412
rect 51675 57409 51687 57443
rect 51629 57403 51687 57409
rect 52086 57400 52092 57452
rect 52144 57440 52150 57452
rect 52365 57443 52423 57449
rect 52365 57440 52377 57443
rect 52144 57412 52377 57440
rect 52144 57400 52150 57412
rect 52365 57409 52377 57412
rect 52411 57409 52423 57443
rect 52365 57403 52423 57409
rect 53282 57400 53288 57452
rect 53340 57440 53346 57452
rect 53561 57443 53619 57449
rect 53561 57440 53573 57443
rect 53340 57412 53573 57440
rect 53340 57400 53346 57412
rect 53561 57409 53573 57412
rect 53607 57440 53619 57443
rect 54021 57443 54079 57449
rect 54021 57440 54033 57443
rect 53607 57412 54033 57440
rect 53607 57409 53619 57412
rect 53561 57403 53619 57409
rect 54021 57409 54033 57412
rect 54067 57409 54079 57443
rect 54021 57403 54079 57409
rect 54478 57400 54484 57452
rect 54536 57440 54542 57452
rect 54757 57443 54815 57449
rect 54757 57440 54769 57443
rect 54536 57412 54769 57440
rect 54536 57400 54542 57412
rect 54757 57409 54769 57412
rect 54803 57409 54815 57443
rect 54757 57403 54815 57409
rect 55674 57400 55680 57452
rect 55732 57440 55738 57452
rect 55953 57443 56011 57449
rect 55953 57440 55965 57443
rect 55732 57412 55965 57440
rect 55732 57400 55738 57412
rect 55953 57409 55965 57412
rect 55999 57440 56011 57443
rect 56413 57443 56471 57449
rect 56413 57440 56425 57443
rect 55999 57412 56425 57440
rect 55999 57409 56011 57412
rect 55953 57403 56011 57409
rect 56413 57409 56425 57412
rect 56459 57409 56471 57443
rect 56413 57403 56471 57409
rect 56870 57400 56876 57452
rect 56928 57440 56934 57452
rect 57149 57443 57207 57449
rect 57149 57440 57161 57443
rect 56928 57412 57161 57440
rect 56928 57400 56934 57412
rect 57149 57409 57161 57412
rect 57195 57409 57207 57443
rect 57149 57403 57207 57409
rect 58066 57400 58072 57452
rect 58124 57440 58130 57452
rect 58345 57443 58403 57449
rect 58345 57440 58357 57443
rect 58124 57412 58357 57440
rect 58124 57400 58130 57412
rect 58345 57409 58357 57412
rect 58391 57409 58403 57443
rect 58345 57403 58403 57409
rect 30374 57372 30380 57384
rect 25700 57344 30380 57372
rect 30374 57332 30380 57344
rect 30432 57332 30438 57384
rect 38378 57332 38384 57384
rect 38436 57372 38442 57384
rect 38436 57344 42748 57372
rect 38436 57332 38442 57344
rect 17727 57276 22094 57304
rect 23661 57307 23719 57313
rect 17727 57273 17739 57276
rect 17681 57267 17739 57273
rect 23661 57273 23673 57307
rect 23707 57304 23719 57307
rect 25038 57304 25044 57316
rect 23707 57276 25044 57304
rect 23707 57273 23719 57276
rect 23661 57267 23719 57273
rect 25038 57264 25044 57276
rect 25096 57264 25102 57316
rect 30837 57307 30895 57313
rect 30837 57273 30849 57307
rect 30883 57304 30895 57307
rect 30883 57276 31754 57304
rect 30883 57273 30895 57276
rect 30837 57267 30895 57273
rect 4525 57239 4583 57245
rect 4525 57205 4537 57239
rect 4571 57236 4583 57239
rect 5442 57236 5448 57248
rect 4571 57208 5448 57236
rect 4571 57205 4583 57208
rect 4525 57199 4583 57205
rect 5442 57196 5448 57208
rect 5500 57196 5506 57248
rect 9306 57236 9312 57248
rect 9267 57208 9312 57236
rect 9306 57196 9312 57208
rect 9364 57196 9370 57248
rect 10502 57236 10508 57248
rect 10463 57208 10508 57236
rect 10502 57196 10508 57208
rect 10560 57196 10566 57248
rect 11882 57236 11888 57248
rect 11843 57208 11888 57236
rect 11882 57196 11888 57208
rect 11940 57196 11946 57248
rect 12894 57236 12900 57248
rect 12855 57208 12900 57236
rect 12894 57196 12900 57208
rect 12952 57196 12958 57248
rect 14458 57236 14464 57248
rect 14419 57208 14464 57236
rect 14458 57196 14464 57208
rect 14516 57196 14522 57248
rect 18874 57236 18880 57248
rect 18835 57208 18880 57236
rect 18874 57196 18880 57208
rect 18932 57196 18938 57248
rect 20070 57236 20076 57248
rect 20031 57208 20076 57236
rect 20070 57196 20076 57208
rect 20128 57196 20134 57248
rect 21266 57236 21272 57248
rect 21227 57208 21272 57236
rect 21266 57196 21272 57208
rect 21324 57196 21330 57248
rect 24854 57236 24860 57248
rect 24815 57208 24860 57236
rect 24854 57196 24860 57208
rect 24912 57196 24918 57248
rect 25866 57236 25872 57248
rect 25827 57208 25872 57236
rect 25866 57196 25872 57208
rect 25924 57196 25930 57248
rect 26142 57196 26148 57248
rect 26200 57236 26206 57248
rect 27157 57239 27215 57245
rect 27157 57236 27169 57239
rect 26200 57208 27169 57236
rect 26200 57196 26206 57208
rect 27157 57205 27169 57208
rect 27203 57205 27215 57239
rect 27157 57199 27215 57205
rect 28350 57196 28356 57248
rect 28408 57236 28414 57248
rect 28445 57239 28503 57245
rect 28445 57236 28457 57239
rect 28408 57208 28457 57236
rect 28408 57196 28414 57208
rect 28445 57205 28457 57208
rect 28491 57205 28503 57239
rect 29730 57236 29736 57248
rect 29691 57208 29736 57236
rect 28445 57199 28503 57205
rect 29730 57196 29736 57208
rect 29788 57196 29794 57248
rect 31726 57236 31754 57276
rect 36446 57264 36452 57316
rect 36504 57304 36510 57316
rect 36504 57276 39160 57304
rect 36504 57264 36510 57276
rect 32306 57236 32312 57248
rect 31726 57208 32312 57236
rect 32306 57196 32312 57208
rect 32364 57196 32370 57248
rect 32493 57239 32551 57245
rect 32493 57205 32505 57239
rect 32539 57236 32551 57239
rect 32950 57236 32956 57248
rect 32539 57208 32956 57236
rect 32539 57205 32551 57208
rect 32493 57199 32551 57205
rect 32950 57196 32956 57208
rect 33008 57196 33014 57248
rect 33226 57236 33232 57248
rect 33187 57208 33232 57236
rect 33226 57196 33232 57208
rect 33284 57196 33290 57248
rect 34698 57196 34704 57248
rect 34756 57236 34762 57248
rect 34885 57239 34943 57245
rect 34885 57236 34897 57239
rect 34756 57208 34897 57236
rect 34756 57196 34762 57208
rect 34885 57205 34897 57208
rect 34931 57205 34943 57239
rect 34885 57199 34943 57205
rect 35713 57239 35771 57245
rect 35713 57205 35725 57239
rect 35759 57236 35771 57239
rect 35802 57236 35808 57248
rect 35759 57208 35808 57236
rect 35759 57205 35771 57208
rect 35713 57199 35771 57205
rect 35802 57196 35808 57208
rect 35860 57196 35866 57248
rect 35894 57196 35900 57248
rect 35952 57236 35958 57248
rect 36633 57239 36691 57245
rect 36633 57236 36645 57239
rect 35952 57208 36645 57236
rect 35952 57196 35958 57208
rect 36633 57205 36645 57208
rect 36679 57205 36691 57239
rect 36633 57199 36691 57205
rect 37642 57196 37648 57248
rect 37700 57236 37706 57248
rect 37829 57239 37887 57245
rect 37829 57236 37841 57239
rect 37700 57208 37841 57236
rect 37700 57196 37706 57208
rect 37829 57205 37841 57208
rect 37875 57205 37887 57239
rect 37829 57199 37887 57205
rect 38654 57196 38660 57248
rect 38712 57236 38718 57248
rect 39025 57239 39083 57245
rect 39025 57236 39037 57239
rect 38712 57208 39037 57236
rect 38712 57196 38718 57208
rect 39025 57205 39037 57208
rect 39071 57205 39083 57239
rect 39132 57236 39160 57276
rect 40221 57239 40279 57245
rect 40221 57236 40233 57239
rect 39132 57208 40233 57236
rect 39025 57199 39083 57205
rect 40221 57205 40233 57208
rect 40267 57205 40279 57239
rect 42720 57236 42748 57344
rect 44542 57332 44548 57384
rect 44600 57372 44606 57384
rect 44600 57344 47808 57372
rect 44600 57332 44606 57344
rect 42794 57264 42800 57316
rect 42852 57304 42858 57316
rect 42852 57276 43944 57304
rect 42852 57264 42858 57276
rect 43809 57239 43867 57245
rect 43809 57236 43821 57239
rect 42720 57208 43821 57236
rect 40221 57199 40279 57205
rect 43809 57205 43821 57208
rect 43855 57205 43867 57239
rect 43916 57236 43944 57276
rect 44634 57264 44640 57316
rect 44692 57304 44698 57316
rect 47780 57313 47808 57344
rect 47765 57307 47823 57313
rect 44692 57276 45554 57304
rect 44692 57264 44698 57276
rect 45189 57239 45247 57245
rect 45189 57236 45201 57239
rect 43916 57208 45201 57236
rect 43809 57199 43867 57205
rect 45189 57205 45201 57208
rect 45235 57205 45247 57239
rect 45526 57236 45554 57276
rect 47765 57273 47777 57307
rect 47811 57273 47823 57307
rect 50985 57307 51043 57313
rect 50985 57304 50997 57307
rect 47765 57267 47823 57273
rect 47872 57276 50997 57304
rect 47872 57236 47900 57276
rect 50985 57273 50997 57276
rect 51031 57273 51043 57307
rect 50985 57267 51043 57273
rect 48590 57236 48596 57248
rect 45526 57208 47900 57236
rect 48551 57208 48596 57236
rect 45189 57199 45247 57205
rect 48590 57196 48596 57208
rect 48648 57196 48654 57248
rect 48682 57196 48688 57248
rect 48740 57236 48746 57248
rect 50341 57239 50399 57245
rect 50341 57236 50353 57239
rect 48740 57208 50353 57236
rect 48740 57196 48746 57208
rect 50341 57205 50353 57208
rect 50387 57205 50399 57239
rect 52178 57236 52184 57248
rect 52139 57208 52184 57236
rect 50341 57199 50399 57205
rect 52178 57196 52184 57208
rect 52236 57196 52242 57248
rect 53374 57236 53380 57248
rect 53335 57208 53380 57236
rect 53374 57196 53380 57208
rect 53432 57196 53438 57248
rect 54570 57236 54576 57248
rect 54531 57208 54576 57236
rect 54570 57196 54576 57208
rect 54628 57196 54634 57248
rect 55766 57236 55772 57248
rect 55727 57208 55772 57236
rect 55766 57196 55772 57208
rect 55824 57196 55830 57248
rect 56962 57236 56968 57248
rect 56923 57208 56968 57236
rect 56962 57196 56968 57208
rect 57020 57196 57026 57248
rect 58158 57236 58164 57248
rect 58119 57208 58164 57236
rect 58158 57196 58164 57208
rect 58216 57196 58222 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 1854 57032 1860 57044
rect 1815 57004 1860 57032
rect 1854 56992 1860 57004
rect 1912 56992 1918 57044
rect 3050 56992 3056 57044
rect 3108 57032 3114 57044
rect 3329 57035 3387 57041
rect 3329 57032 3341 57035
rect 3108 57004 3341 57032
rect 3108 56992 3114 57004
rect 3329 57001 3341 57004
rect 3375 57001 3387 57035
rect 3329 56995 3387 57001
rect 4249 57035 4307 57041
rect 4249 57001 4261 57035
rect 4295 57032 4307 57035
rect 4614 57032 4620 57044
rect 4295 57004 4620 57032
rect 4295 57001 4307 57004
rect 4249 56995 4307 57001
rect 4614 56992 4620 57004
rect 4672 56992 4678 57044
rect 8478 57032 8484 57044
rect 8439 57004 8484 57032
rect 8478 56992 8484 57004
rect 8536 56992 8542 57044
rect 9030 56992 9036 57044
rect 9088 57032 9094 57044
rect 9125 57035 9183 57041
rect 9125 57032 9137 57035
rect 9088 57004 9137 57032
rect 9088 56992 9094 57004
rect 9125 57001 9137 57004
rect 9171 57001 9183 57035
rect 12618 57032 12624 57044
rect 12579 57004 12624 57032
rect 9125 56995 9183 57001
rect 12618 56992 12624 57004
rect 12676 56992 12682 57044
rect 15010 57032 15016 57044
rect 14971 57004 15016 57032
rect 15010 56992 15016 57004
rect 15068 56992 15074 57044
rect 17402 57032 17408 57044
rect 17363 57004 17408 57032
rect 17402 56992 17408 57004
rect 17460 56992 17466 57044
rect 19797 57035 19855 57041
rect 19797 57001 19809 57035
rect 19843 57032 19855 57035
rect 19978 57032 19984 57044
rect 19843 57004 19984 57032
rect 19843 57001 19855 57004
rect 19797 56995 19855 57001
rect 19978 56992 19984 57004
rect 20036 56992 20042 57044
rect 22186 57032 22192 57044
rect 22147 57004 22192 57032
rect 22186 56992 22192 57004
rect 22244 56992 22250 57044
rect 24578 57032 24584 57044
rect 24539 57004 24584 57032
rect 24578 56992 24584 57004
rect 24636 56992 24642 57044
rect 28166 57032 28172 57044
rect 28127 57004 28172 57032
rect 28166 56992 28172 57004
rect 28224 56992 28230 57044
rect 32122 57032 32128 57044
rect 32083 57004 32128 57032
rect 32122 56992 32128 57004
rect 32180 56992 32186 57044
rect 35342 57032 35348 57044
rect 35303 57004 35348 57032
rect 35342 56992 35348 57004
rect 35400 56992 35406 57044
rect 36538 57032 36544 57044
rect 36499 57004 36544 57032
rect 36538 56992 36544 57004
rect 36596 56992 36602 57044
rect 38105 57035 38163 57041
rect 38105 57001 38117 57035
rect 38151 57032 38163 57035
rect 38930 57032 38936 57044
rect 38151 57004 38936 57032
rect 38151 57001 38163 57004
rect 38105 56995 38163 57001
rect 38930 56992 38936 57004
rect 38988 56992 38994 57044
rect 41322 57032 41328 57044
rect 41283 57004 41328 57032
rect 41322 56992 41328 57004
rect 41380 56992 41386 57044
rect 44910 56992 44916 57044
rect 44968 57032 44974 57044
rect 45189 57035 45247 57041
rect 45189 57032 45201 57035
rect 44968 57004 45201 57032
rect 44968 56992 44974 57004
rect 45189 57001 45201 57004
rect 45235 57001 45247 57035
rect 45189 56995 45247 57001
rect 47302 56992 47308 57044
rect 47360 57032 47366 57044
rect 47581 57035 47639 57041
rect 47581 57032 47593 57035
rect 47360 57004 47593 57032
rect 47360 56992 47366 57004
rect 47581 57001 47593 57004
rect 47627 57001 47639 57035
rect 50338 57032 50344 57044
rect 50299 57004 50344 57032
rect 47581 56995 47639 57001
rect 50338 56992 50344 57004
rect 50396 56992 50402 57044
rect 52086 57032 52092 57044
rect 52047 57004 52092 57032
rect 52086 56992 52092 57004
rect 52144 56992 52150 57044
rect 54478 57032 54484 57044
rect 54439 57004 54484 57032
rect 54478 56992 54484 57004
rect 54536 56992 54542 57044
rect 56413 57035 56471 57041
rect 56413 57001 56425 57035
rect 56459 57032 56471 57035
rect 56870 57032 56876 57044
rect 56459 57004 56876 57032
rect 56459 57001 56471 57004
rect 56413 56995 56471 57001
rect 56870 56992 56876 57004
rect 56928 56992 56934 57044
rect 9306 56924 9312 56976
rect 9364 56964 9370 56976
rect 17218 56964 17224 56976
rect 9364 56936 17224 56964
rect 9364 56924 9370 56936
rect 17218 56924 17224 56936
rect 17276 56924 17282 56976
rect 21545 56967 21603 56973
rect 21545 56933 21557 56967
rect 21591 56964 21603 56967
rect 29178 56964 29184 56976
rect 21591 56936 29184 56964
rect 21591 56933 21603 56936
rect 21545 56927 21603 56933
rect 29178 56924 29184 56936
rect 29236 56924 29242 56976
rect 37826 56924 37832 56976
rect 37884 56964 37890 56976
rect 43257 56967 43315 56973
rect 43257 56964 43269 56967
rect 37884 56936 43269 56964
rect 37884 56924 37890 56936
rect 43257 56933 43269 56936
rect 43303 56933 43315 56967
rect 43257 56927 43315 56933
rect 44726 56924 44732 56976
rect 44784 56964 44790 56976
rect 48590 56964 48596 56976
rect 44784 56936 48596 56964
rect 44784 56924 44790 56936
rect 48590 56924 48596 56936
rect 48648 56924 48654 56976
rect 6273 56899 6331 56905
rect 6273 56865 6285 56899
rect 6319 56896 6331 56899
rect 6638 56896 6644 56908
rect 6319 56868 6644 56896
rect 6319 56865 6331 56868
rect 6273 56859 6331 56865
rect 6638 56856 6644 56868
rect 6696 56896 6702 56908
rect 6733 56899 6791 56905
rect 6733 56896 6745 56899
rect 6696 56868 6745 56896
rect 6696 56856 6702 56868
rect 6733 56865 6745 56868
rect 6779 56865 6791 56899
rect 6733 56859 6791 56865
rect 10502 56856 10508 56908
rect 10560 56896 10566 56908
rect 17954 56896 17960 56908
rect 10560 56868 17960 56896
rect 10560 56856 10566 56868
rect 17954 56856 17960 56868
rect 18012 56856 18018 56908
rect 20070 56856 20076 56908
rect 20128 56896 20134 56908
rect 26234 56896 26240 56908
rect 20128 56868 26240 56896
rect 20128 56856 20134 56868
rect 26234 56856 26240 56868
rect 26292 56856 26298 56908
rect 29730 56896 29736 56908
rect 29691 56868 29736 56896
rect 29730 56856 29736 56868
rect 29788 56856 29794 56908
rect 48682 56896 48688 56908
rect 43824 56868 48688 56896
rect 7006 56828 7012 56840
rect 6967 56800 7012 56828
rect 7006 56788 7012 56800
rect 7064 56788 7070 56840
rect 11882 56788 11888 56840
rect 11940 56828 11946 56840
rect 19334 56828 19340 56840
rect 11940 56800 19340 56828
rect 11940 56788 11946 56800
rect 19334 56788 19340 56800
rect 19392 56788 19398 56840
rect 21266 56788 21272 56840
rect 21324 56828 21330 56840
rect 29362 56828 29368 56840
rect 21324 56800 29368 56828
rect 21324 56788 21330 56800
rect 29362 56788 29368 56800
rect 29420 56788 29426 56840
rect 29822 56828 29828 56840
rect 29783 56800 29828 56828
rect 29822 56788 29828 56800
rect 29880 56788 29886 56840
rect 30009 56831 30067 56837
rect 30009 56797 30021 56831
rect 30055 56797 30067 56831
rect 38746 56828 38752 56840
rect 38710 56800 38752 56828
rect 30009 56791 30067 56797
rect 12894 56720 12900 56772
rect 12952 56760 12958 56772
rect 20806 56760 20812 56772
rect 12952 56732 20812 56760
rect 12952 56720 12958 56732
rect 20806 56720 20812 56732
rect 20864 56720 20870 56772
rect 21174 56760 21180 56772
rect 21135 56732 21180 56760
rect 21174 56720 21180 56732
rect 21232 56720 21238 56772
rect 21361 56763 21419 56769
rect 21361 56729 21373 56763
rect 21407 56729 21419 56763
rect 21361 56723 21419 56729
rect 14458 56652 14464 56704
rect 14516 56692 14522 56704
rect 21376 56692 21404 56723
rect 29454 56720 29460 56772
rect 29512 56760 29518 56772
rect 30024 56760 30052 56791
rect 38746 56788 38752 56800
rect 38804 56788 38810 56840
rect 38873 56831 38931 56837
rect 38873 56828 38885 56831
rect 38856 56797 38885 56828
rect 38919 56797 38931 56831
rect 38856 56791 38931 56797
rect 38984 56831 39042 56837
rect 38984 56797 38996 56831
rect 39030 56828 39042 56831
rect 39030 56818 39068 56828
rect 38984 56791 39028 56797
rect 38856 56760 38884 56791
rect 39022 56766 39028 56791
rect 39080 56766 39086 56818
rect 39114 56788 39120 56840
rect 39172 56828 39178 56840
rect 39172 56800 39217 56828
rect 39172 56788 39178 56800
rect 43346 56788 43352 56840
rect 43404 56837 43410 56840
rect 43824 56837 43852 56868
rect 48682 56856 48688 56868
rect 48740 56856 48746 56908
rect 55861 56899 55919 56905
rect 55861 56865 55873 56899
rect 55907 56896 55919 56899
rect 55907 56868 58388 56896
rect 55907 56865 55919 56868
rect 55861 56859 55919 56865
rect 58360 56840 58388 56868
rect 43404 56831 43453 56837
rect 43404 56797 43407 56831
rect 43441 56797 43453 56831
rect 43404 56791 43453 56797
rect 43533 56831 43591 56837
rect 43533 56797 43545 56831
rect 43579 56828 43591 56831
rect 43808 56831 43866 56837
rect 43579 56800 43760 56828
rect 43579 56797 43591 56800
rect 43533 56791 43591 56797
rect 43404 56788 43410 56791
rect 43622 56760 43628 56772
rect 29512 56732 30052 56760
rect 38764 56732 38884 56760
rect 43583 56732 43628 56760
rect 29512 56720 29518 56732
rect 38764 56704 38792 56732
rect 43622 56720 43628 56732
rect 43680 56720 43686 56772
rect 43732 56760 43760 56800
rect 43808 56797 43820 56831
rect 43854 56797 43866 56831
rect 43808 56791 43866 56797
rect 43898 56788 43904 56840
rect 43956 56828 43962 56840
rect 57054 56828 57060 56840
rect 43956 56800 44001 56828
rect 57015 56800 57060 56828
rect 43956 56788 43962 56800
rect 57054 56788 57060 56800
rect 57112 56788 57118 56840
rect 57514 56828 57520 56840
rect 57475 56800 57520 56828
rect 57514 56788 57520 56800
rect 57572 56788 57578 56840
rect 58342 56828 58348 56840
rect 58303 56800 58348 56828
rect 58342 56788 58348 56800
rect 58400 56788 58406 56840
rect 56962 56760 56968 56772
rect 43732 56732 56968 56760
rect 56962 56720 56968 56732
rect 57020 56720 57026 56772
rect 30190 56692 30196 56704
rect 14516 56664 21404 56692
rect 30151 56664 30196 56692
rect 14516 56652 14522 56664
rect 30190 56652 30196 56664
rect 30248 56652 30254 56704
rect 35986 56652 35992 56704
rect 36044 56692 36050 56704
rect 38565 56695 38623 56701
rect 38565 56692 38577 56695
rect 36044 56664 38577 56692
rect 36044 56652 36050 56664
rect 38565 56661 38577 56664
rect 38611 56661 38623 56695
rect 38565 56655 38623 56661
rect 38746 56652 38752 56704
rect 38804 56652 38810 56704
rect 56870 56692 56876 56704
rect 56831 56664 56876 56692
rect 56870 56652 56876 56664
rect 56928 56652 56934 56704
rect 57698 56692 57704 56704
rect 57659 56664 57704 56692
rect 57698 56652 57704 56664
rect 57756 56652 57762 56704
rect 58161 56695 58219 56701
rect 58161 56661 58173 56695
rect 58207 56692 58219 56695
rect 59170 56692 59176 56704
rect 58207 56664 59176 56692
rect 58207 56661 58219 56664
rect 58161 56655 58219 56661
rect 59170 56652 59176 56664
rect 59228 56652 59234 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 17218 56448 17224 56500
rect 17276 56488 17282 56500
rect 17276 56460 22094 56488
rect 17276 56448 17282 56460
rect 17954 56380 17960 56432
rect 18012 56420 18018 56432
rect 21269 56423 21327 56429
rect 21269 56420 21281 56423
rect 18012 56392 21281 56420
rect 18012 56380 18018 56392
rect 21269 56389 21281 56392
rect 21315 56389 21327 56423
rect 22066 56420 22094 56460
rect 24946 56448 24952 56500
rect 25004 56488 25010 56500
rect 26513 56491 26571 56497
rect 25004 56460 26280 56488
rect 25004 56448 25010 56460
rect 22189 56423 22247 56429
rect 22189 56420 22201 56423
rect 22066 56392 22201 56420
rect 21269 56383 21327 56389
rect 22189 56389 22201 56392
rect 22235 56389 22247 56423
rect 25314 56420 25320 56432
rect 22189 56383 22247 56389
rect 24135 56392 25320 56420
rect 21085 56355 21143 56361
rect 21085 56321 21097 56355
rect 21131 56352 21143 56355
rect 21174 56352 21180 56364
rect 21131 56324 21180 56352
rect 21131 56321 21143 56324
rect 21085 56315 21143 56321
rect 21174 56312 21180 56324
rect 21232 56352 21238 56364
rect 21910 56352 21916 56364
rect 21232 56324 21916 56352
rect 21232 56312 21238 56324
rect 21910 56312 21916 56324
rect 21968 56352 21974 56364
rect 23750 56361 23756 56364
rect 22005 56355 22063 56361
rect 22005 56352 22017 56355
rect 21968 56324 22017 56352
rect 21968 56312 21974 56324
rect 22005 56321 22017 56324
rect 22051 56321 22063 56355
rect 23748 56352 23756 56361
rect 23711 56324 23756 56352
rect 22005 56315 22063 56321
rect 23748 56315 23756 56324
rect 23750 56312 23756 56315
rect 23808 56312 23814 56364
rect 24135 56361 24163 56392
rect 25314 56380 25320 56392
rect 25372 56380 25378 56432
rect 26252 56429 26280 56460
rect 26513 56457 26525 56491
rect 26559 56488 26571 56491
rect 26559 56460 27384 56488
rect 26559 56457 26571 56460
rect 26513 56451 26571 56457
rect 27356 56429 27384 56460
rect 27430 56448 27436 56500
rect 27488 56488 27494 56500
rect 30466 56488 30472 56500
rect 27488 56460 30472 56488
rect 27488 56448 27494 56460
rect 25409 56423 25467 56429
rect 25409 56389 25421 56423
rect 25455 56420 25467 56423
rect 26237 56423 26295 56429
rect 25455 56392 26004 56420
rect 25455 56389 25467 56392
rect 25409 56383 25467 56389
rect 23845 56355 23903 56361
rect 23845 56321 23857 56355
rect 23891 56321 23903 56355
rect 23845 56315 23903 56321
rect 23937 56355 23995 56361
rect 23937 56321 23949 56355
rect 23983 56321 23995 56355
rect 23937 56315 23995 56321
rect 24120 56355 24178 56361
rect 24120 56321 24132 56355
rect 24166 56321 24178 56355
rect 24120 56315 24178 56321
rect 20714 56244 20720 56296
rect 20772 56284 20778 56296
rect 23860 56284 23888 56315
rect 20772 56256 23888 56284
rect 23952 56284 23980 56315
rect 24210 56312 24216 56364
rect 24268 56352 24274 56364
rect 24268 56324 24313 56352
rect 24268 56312 24274 56324
rect 24854 56312 24860 56364
rect 24912 56352 24918 56364
rect 24949 56355 25007 56361
rect 24949 56352 24961 56355
rect 24912 56324 24961 56352
rect 24912 56312 24918 56324
rect 24949 56321 24961 56324
rect 24995 56321 25007 56355
rect 25222 56352 25228 56364
rect 25183 56324 25228 56352
rect 24949 56315 25007 56321
rect 25222 56312 25228 56324
rect 25280 56312 25286 56364
rect 25774 56312 25780 56364
rect 25832 56352 25838 56364
rect 25976 56361 26004 56392
rect 26237 56389 26249 56423
rect 26283 56389 26295 56423
rect 26237 56383 26295 56389
rect 27341 56423 27399 56429
rect 27341 56389 27353 56423
rect 27387 56389 27399 56423
rect 27341 56383 27399 56389
rect 29109 56423 29167 56429
rect 29109 56389 29121 56423
rect 29155 56420 29167 56423
rect 29362 56420 29368 56432
rect 29155 56392 29368 56420
rect 29155 56389 29167 56392
rect 29109 56383 29167 56389
rect 29362 56380 29368 56392
rect 29420 56380 29426 56432
rect 26418 56361 26424 56364
rect 25869 56355 25927 56361
rect 25869 56352 25881 56355
rect 25832 56324 25881 56352
rect 25832 56312 25838 56324
rect 25869 56321 25881 56324
rect 25915 56321 25927 56355
rect 25869 56315 25927 56321
rect 25962 56355 26020 56361
rect 25962 56321 25974 56355
rect 26008 56321 26020 56355
rect 25962 56315 26020 56321
rect 26145 56355 26203 56361
rect 26145 56321 26157 56355
rect 26191 56321 26203 56355
rect 26145 56315 26203 56321
rect 26375 56355 26424 56361
rect 26375 56321 26387 56355
rect 26421 56321 26424 56355
rect 26375 56315 26424 56321
rect 24578 56284 24584 56296
rect 23952 56256 24584 56284
rect 20772 56244 20778 56256
rect 24578 56244 24584 56256
rect 24636 56244 24642 56296
rect 26160 56284 26188 56315
rect 26418 56312 26424 56315
rect 26476 56312 26482 56364
rect 27203 56355 27261 56361
rect 27203 56352 27215 56355
rect 27126 56324 27215 56352
rect 26878 56284 26884 56296
rect 25148 56256 26096 56284
rect 26160 56256 26884 56284
rect 21453 56219 21511 56225
rect 21453 56185 21465 56219
rect 21499 56216 21511 56219
rect 25148 56216 25176 56256
rect 21499 56188 25176 56216
rect 26068 56216 26096 56256
rect 26878 56244 26884 56256
rect 26936 56244 26942 56296
rect 27126 56216 27154 56324
rect 27203 56321 27215 56324
rect 27249 56321 27261 56355
rect 27203 56315 27261 56321
rect 27433 56355 27491 56361
rect 27433 56321 27445 56355
rect 27479 56321 27491 56355
rect 27433 56315 27491 56321
rect 27338 56244 27344 56296
rect 27396 56284 27402 56296
rect 27448 56284 27476 56315
rect 27522 56312 27528 56364
rect 27580 56361 27586 56364
rect 27580 56352 27588 56361
rect 28721 56355 28779 56361
rect 27580 56324 27625 56352
rect 27580 56315 27588 56324
rect 28721 56321 28733 56355
rect 28767 56321 28779 56355
rect 28721 56315 28779 56321
rect 27580 56312 27586 56315
rect 27396 56256 27476 56284
rect 27396 56244 27402 56256
rect 28534 56244 28540 56296
rect 28592 56284 28598 56296
rect 28736 56284 28764 56315
rect 28810 56312 28816 56364
rect 28868 56352 28874 56364
rect 28868 56324 28913 56352
rect 28868 56312 28874 56324
rect 28948 56318 28954 56370
rect 29006 56352 29012 56370
rect 29227 56355 29285 56361
rect 29006 56324 29045 56352
rect 29006 56318 29012 56324
rect 29227 56321 29239 56355
rect 29273 56352 29285 56355
rect 29656 56352 29684 56460
rect 30466 56448 30472 56460
rect 30524 56448 30530 56500
rect 30653 56491 30711 56497
rect 30653 56457 30665 56491
rect 30699 56488 30711 56491
rect 30699 56460 31340 56488
rect 30699 56457 30711 56460
rect 30653 56451 30711 56457
rect 30285 56423 30343 56429
rect 30285 56389 30297 56423
rect 30331 56420 30343 56423
rect 31018 56420 31024 56432
rect 30331 56392 31024 56420
rect 30331 56389 30343 56392
rect 30285 56383 30343 56389
rect 31018 56380 31024 56392
rect 31076 56380 31082 56432
rect 31312 56429 31340 56460
rect 31386 56448 31392 56500
rect 31444 56488 31450 56500
rect 34425 56491 34483 56497
rect 34425 56488 34437 56491
rect 31444 56460 34437 56488
rect 31444 56448 31450 56460
rect 34425 56457 34437 56460
rect 34471 56457 34483 56491
rect 34425 56451 34483 56457
rect 34974 56448 34980 56500
rect 35032 56488 35038 56500
rect 35986 56488 35992 56500
rect 35032 56460 35992 56488
rect 35032 56448 35038 56460
rect 35986 56448 35992 56460
rect 36044 56448 36050 56500
rect 38010 56448 38016 56500
rect 38068 56488 38074 56500
rect 44634 56488 44640 56500
rect 38068 56460 39068 56488
rect 38068 56448 38074 56460
rect 31297 56423 31355 56429
rect 31297 56389 31309 56423
rect 31343 56389 31355 56423
rect 31297 56383 31355 56389
rect 32306 56380 32312 56432
rect 32364 56420 32370 56432
rect 32861 56423 32919 56429
rect 32861 56420 32873 56423
rect 32364 56392 32873 56420
rect 32364 56380 32370 56392
rect 32861 56389 32873 56392
rect 32907 56389 32919 56423
rect 34514 56420 34520 56432
rect 32861 56383 32919 56389
rect 33152 56392 34520 56420
rect 30190 56361 30196 56364
rect 29273 56324 29684 56352
rect 30009 56355 30067 56361
rect 29273 56321 29285 56324
rect 28951 56315 29009 56318
rect 29227 56315 29285 56321
rect 30009 56321 30021 56355
rect 30055 56321 30067 56355
rect 30009 56315 30067 56321
rect 30157 56355 30196 56361
rect 30157 56321 30169 56355
rect 30157 56315 30196 56321
rect 30024 56284 30052 56315
rect 30190 56312 30196 56315
rect 30248 56312 30254 56364
rect 30374 56352 30380 56364
rect 30335 56324 30380 56352
rect 30374 56312 30380 56324
rect 30432 56312 30438 56364
rect 30466 56312 30472 56364
rect 30524 56361 30530 56364
rect 30524 56352 30532 56361
rect 30524 56324 30569 56352
rect 30524 56315 30532 56324
rect 30524 56312 30530 56315
rect 30650 56312 30656 56364
rect 30708 56352 30714 56364
rect 31113 56355 31171 56361
rect 31113 56352 31125 56355
rect 30708 56324 31125 56352
rect 30708 56312 30714 56324
rect 31113 56321 31125 56324
rect 31159 56321 31171 56355
rect 31113 56315 31171 56321
rect 31202 56312 31208 56364
rect 31260 56352 31266 56364
rect 31389 56355 31447 56361
rect 31389 56352 31401 56355
rect 31260 56324 31401 56352
rect 31260 56312 31266 56324
rect 31389 56321 31401 56324
rect 31435 56321 31447 56355
rect 31389 56315 31447 56321
rect 31533 56355 31591 56361
rect 31533 56321 31545 56355
rect 31579 56352 31591 56355
rect 31662 56352 31668 56364
rect 31579 56324 31668 56352
rect 31579 56321 31591 56324
rect 31533 56315 31591 56321
rect 31662 56312 31668 56324
rect 31720 56312 31726 56364
rect 32766 56361 32772 56364
rect 32764 56352 32772 56361
rect 32727 56324 32772 56352
rect 32764 56315 32772 56324
rect 32766 56312 32772 56315
rect 32824 56312 32830 56364
rect 32953 56355 33011 56361
rect 32953 56321 32965 56355
rect 32999 56352 33011 56355
rect 33042 56352 33048 56364
rect 32999 56324 33048 56352
rect 32999 56321 33011 56324
rect 32953 56315 33011 56321
rect 33042 56312 33048 56324
rect 33100 56312 33106 56364
rect 33152 56361 33180 56392
rect 34514 56380 34520 56392
rect 34572 56380 34578 56432
rect 34698 56420 34704 56432
rect 34659 56392 34704 56420
rect 34698 56380 34704 56392
rect 34756 56380 34762 56432
rect 34793 56423 34851 56429
rect 34793 56389 34805 56423
rect 34839 56420 34851 56423
rect 35802 56420 35808 56432
rect 34839 56392 35664 56420
rect 35763 56392 35808 56420
rect 34839 56389 34851 56392
rect 34793 56383 34851 56389
rect 33136 56355 33194 56361
rect 33136 56321 33148 56355
rect 33182 56321 33194 56355
rect 33136 56315 33194 56321
rect 33229 56355 33287 56361
rect 33229 56321 33241 56355
rect 33275 56352 33287 56355
rect 33318 56352 33324 56364
rect 33275 56324 33324 56352
rect 33275 56321 33287 56324
rect 33229 56315 33287 56321
rect 33318 56312 33324 56324
rect 33376 56312 33382 56364
rect 34606 56361 34612 56364
rect 34604 56352 34612 56361
rect 34567 56324 34612 56352
rect 34604 56315 34612 56324
rect 34606 56312 34612 56315
rect 34664 56312 34670 56364
rect 34974 56352 34980 56364
rect 34935 56324 34980 56352
rect 34974 56312 34980 56324
rect 35032 56312 35038 56364
rect 35066 56312 35072 56364
rect 35124 56352 35130 56364
rect 35526 56352 35532 56364
rect 35124 56324 35532 56352
rect 35124 56312 35130 56324
rect 35526 56312 35532 56324
rect 35584 56312 35590 56364
rect 30834 56284 30840 56296
rect 28592 56256 30840 56284
rect 28592 56244 28598 56256
rect 30834 56244 30840 56256
rect 30892 56244 30898 56296
rect 35636 56284 35664 56392
rect 35802 56380 35808 56392
rect 35860 56380 35866 56432
rect 35897 56423 35955 56429
rect 35897 56389 35909 56423
rect 35943 56420 35955 56423
rect 37826 56420 37832 56432
rect 35943 56392 37832 56420
rect 35943 56389 35955 56392
rect 35897 56383 35955 56389
rect 37826 56380 37832 56392
rect 37884 56380 37890 56432
rect 37936 56392 38976 56420
rect 35710 56361 35716 56364
rect 35708 56315 35716 56361
rect 35768 56352 35774 56364
rect 36078 56352 36084 56364
rect 35768 56324 35808 56352
rect 36039 56324 36084 56352
rect 35710 56312 35716 56315
rect 35768 56312 35774 56324
rect 36078 56312 36084 56324
rect 36136 56312 36142 56364
rect 36170 56312 36176 56364
rect 36228 56352 36234 56364
rect 37642 56352 37648 56364
rect 36228 56324 36273 56352
rect 37603 56324 37648 56352
rect 36228 56312 36234 56324
rect 37642 56312 37648 56324
rect 37700 56312 37706 56364
rect 37734 56312 37740 56364
rect 37792 56352 37798 56364
rect 37936 56361 37964 56392
rect 38948 56364 38976 56392
rect 39040 56364 39068 56460
rect 43732 56460 44640 56488
rect 42702 56420 42708 56432
rect 41156 56392 42708 56420
rect 37921 56355 37979 56361
rect 37792 56324 37837 56352
rect 37792 56312 37798 56324
rect 37921 56321 37933 56355
rect 37967 56321 37979 56355
rect 37921 56315 37979 56321
rect 38010 56312 38016 56364
rect 38068 56352 38074 56364
rect 38654 56352 38660 56364
rect 38068 56324 38113 56352
rect 38615 56324 38660 56352
rect 38068 56312 38074 56324
rect 38654 56312 38660 56324
rect 38712 56312 38718 56364
rect 38746 56312 38752 56364
rect 38804 56352 38810 56364
rect 38930 56352 38936 56364
rect 38804 56324 38849 56352
rect 38891 56324 38936 56352
rect 38804 56312 38810 56324
rect 38930 56312 38936 56324
rect 38988 56312 38994 56364
rect 39022 56312 39028 56364
rect 39080 56352 39086 56364
rect 40770 56361 40776 56364
rect 40768 56352 40776 56361
rect 39080 56324 39125 56352
rect 40731 56324 40776 56352
rect 39080 56312 39086 56324
rect 40768 56315 40776 56324
rect 40770 56312 40776 56315
rect 40828 56312 40834 56364
rect 40865 56355 40923 56361
rect 40865 56321 40877 56355
rect 40911 56321 40923 56355
rect 40865 56315 40923 56321
rect 40494 56284 40500 56296
rect 35636 56256 40500 56284
rect 40494 56244 40500 56256
rect 40552 56244 40558 56296
rect 28626 56216 28632 56228
rect 26068 56188 27154 56216
rect 27264 56188 28632 56216
rect 21499 56185 21511 56188
rect 21453 56179 21511 56185
rect 22373 56151 22431 56157
rect 22373 56117 22385 56151
rect 22419 56148 22431 56151
rect 23382 56148 23388 56160
rect 22419 56120 23388 56148
rect 22419 56117 22431 56120
rect 22373 56111 22431 56117
rect 23382 56108 23388 56120
rect 23440 56108 23446 56160
rect 23566 56148 23572 56160
rect 23527 56120 23572 56148
rect 23566 56108 23572 56120
rect 23624 56108 23630 56160
rect 25041 56151 25099 56157
rect 25041 56117 25053 56151
rect 25087 56148 25099 56151
rect 25130 56148 25136 56160
rect 25087 56120 25136 56148
rect 25087 56117 25099 56120
rect 25041 56111 25099 56117
rect 25130 56108 25136 56120
rect 25188 56108 25194 56160
rect 25314 56108 25320 56160
rect 25372 56148 25378 56160
rect 27264 56148 27292 56188
rect 28626 56176 28632 56188
rect 28684 56176 28690 56228
rect 29365 56219 29423 56225
rect 29365 56185 29377 56219
rect 29411 56216 29423 56219
rect 31665 56219 31723 56225
rect 29411 56188 29500 56216
rect 29411 56185 29423 56188
rect 29365 56179 29423 56185
rect 25372 56120 27292 56148
rect 27709 56151 27767 56157
rect 25372 56108 25378 56120
rect 27709 56117 27721 56151
rect 27755 56148 27767 56151
rect 28718 56148 28724 56160
rect 27755 56120 28724 56148
rect 27755 56117 27767 56120
rect 27709 56111 27767 56117
rect 28718 56108 28724 56120
rect 28776 56108 28782 56160
rect 29472 56148 29500 56188
rect 31665 56185 31677 56219
rect 31711 56216 31723 56219
rect 33134 56216 33140 56228
rect 31711 56188 33140 56216
rect 31711 56185 31723 56188
rect 31665 56179 31723 56185
rect 33134 56176 33140 56188
rect 33192 56176 33198 56228
rect 33318 56176 33324 56228
rect 33376 56216 33382 56228
rect 35066 56216 35072 56228
rect 33376 56188 35072 56216
rect 33376 56176 33382 56188
rect 35066 56176 35072 56188
rect 35124 56176 35130 56228
rect 35158 56176 35164 56228
rect 35216 56216 35222 56228
rect 35529 56219 35587 56225
rect 35529 56216 35541 56219
rect 35216 56188 35541 56216
rect 35216 56176 35222 56188
rect 35529 56185 35541 56188
rect 35575 56185 35587 56219
rect 35529 56179 35587 56185
rect 35618 56176 35624 56228
rect 35676 56216 35682 56228
rect 40589 56219 40647 56225
rect 40589 56216 40601 56219
rect 35676 56188 40601 56216
rect 35676 56176 35682 56188
rect 40589 56185 40601 56188
rect 40635 56185 40647 56219
rect 40880 56216 40908 56315
rect 40954 56312 40960 56364
rect 41012 56352 41018 56364
rect 41156 56361 41184 56392
rect 42702 56380 42708 56392
rect 42760 56380 42766 56432
rect 42978 56380 42984 56432
rect 43036 56420 43042 56432
rect 43533 56423 43591 56429
rect 43533 56420 43545 56423
rect 43036 56392 43545 56420
rect 43036 56380 43042 56392
rect 43533 56389 43545 56392
rect 43579 56420 43591 56423
rect 43622 56420 43628 56432
rect 43579 56392 43628 56420
rect 43579 56389 43591 56392
rect 43533 56383 43591 56389
rect 43622 56380 43628 56392
rect 43680 56380 43686 56432
rect 41140 56355 41198 56361
rect 41012 56324 41057 56352
rect 41012 56312 41018 56324
rect 41140 56321 41152 56355
rect 41186 56321 41198 56355
rect 41140 56315 41198 56321
rect 41230 56312 41236 56364
rect 41288 56352 41294 56364
rect 41288 56324 41333 56352
rect 41288 56312 41294 56324
rect 42610 56312 42616 56364
rect 42668 56352 42674 56364
rect 43346 56361 43352 56364
rect 43303 56355 43352 56361
rect 43303 56352 43315 56355
rect 42668 56324 43315 56352
rect 42668 56312 42674 56324
rect 43303 56321 43315 56324
rect 43349 56321 43352 56355
rect 43303 56315 43352 56321
rect 43346 56312 43352 56315
rect 43404 56312 43410 56364
rect 43732 56361 43760 56460
rect 44634 56448 44640 56460
rect 44692 56448 44698 56500
rect 57054 56448 57060 56500
rect 57112 56488 57118 56500
rect 57149 56491 57207 56497
rect 57149 56488 57161 56491
rect 57112 56460 57161 56488
rect 57112 56448 57118 56460
rect 57149 56457 57161 56460
rect 57195 56457 57207 56491
rect 57149 56451 57207 56457
rect 56689 56423 56747 56429
rect 56689 56389 56701 56423
rect 56735 56420 56747 56423
rect 57514 56420 57520 56432
rect 56735 56392 57520 56420
rect 56735 56389 56747 56392
rect 56689 56383 56747 56389
rect 57514 56380 57520 56392
rect 57572 56380 57578 56432
rect 43441 56355 43499 56361
rect 43441 56321 43453 56355
rect 43487 56321 43499 56355
rect 43441 56315 43499 56321
rect 43716 56355 43774 56361
rect 43716 56321 43728 56355
rect 43762 56321 43774 56355
rect 43716 56315 43774 56321
rect 43809 56355 43867 56361
rect 43809 56321 43821 56355
rect 43855 56352 43867 56355
rect 43898 56352 43904 56364
rect 43855 56324 43904 56352
rect 43855 56321 43867 56324
rect 43809 56315 43867 56321
rect 43456 56284 43484 56315
rect 43898 56312 43904 56324
rect 43956 56312 43962 56364
rect 56137 56355 56195 56361
rect 56137 56321 56149 56355
rect 56183 56352 56195 56355
rect 58066 56352 58072 56364
rect 56183 56324 58072 56352
rect 56183 56321 56195 56324
rect 56137 56315 56195 56321
rect 58066 56312 58072 56324
rect 58124 56312 58130 56364
rect 58345 56355 58403 56361
rect 58345 56321 58357 56355
rect 58391 56352 58403 56355
rect 58434 56352 58440 56364
rect 58391 56324 58440 56352
rect 58391 56321 58403 56324
rect 58345 56315 58403 56321
rect 58434 56312 58440 56324
rect 58492 56312 58498 56364
rect 58158 56284 58164 56296
rect 43456 56256 58164 56284
rect 58158 56244 58164 56256
rect 58216 56244 58222 56296
rect 53374 56216 53380 56228
rect 40880 56188 53380 56216
rect 40589 56179 40647 56185
rect 53374 56176 53380 56188
rect 53432 56176 53438 56228
rect 29914 56148 29920 56160
rect 29472 56120 29920 56148
rect 29914 56108 29920 56120
rect 29972 56108 29978 56160
rect 32582 56148 32588 56160
rect 32543 56120 32588 56148
rect 32582 56108 32588 56120
rect 32640 56108 32646 56160
rect 33042 56108 33048 56160
rect 33100 56148 33106 56160
rect 37461 56151 37519 56157
rect 37461 56148 37473 56151
rect 33100 56120 37473 56148
rect 33100 56108 33106 56120
rect 37461 56117 37473 56120
rect 37507 56117 37519 56151
rect 37461 56111 37519 56117
rect 37550 56108 37556 56160
rect 37608 56148 37614 56160
rect 38473 56151 38531 56157
rect 38473 56148 38485 56151
rect 37608 56120 38485 56148
rect 37608 56108 37614 56120
rect 38473 56117 38485 56120
rect 38519 56117 38531 56151
rect 38473 56111 38531 56117
rect 38654 56108 38660 56160
rect 38712 56148 38718 56160
rect 41138 56148 41144 56160
rect 38712 56120 41144 56148
rect 38712 56108 38718 56120
rect 41138 56108 41144 56120
rect 41196 56108 41202 56160
rect 43162 56148 43168 56160
rect 43123 56120 43168 56148
rect 43162 56108 43168 56120
rect 43220 56108 43226 56160
rect 58158 56148 58164 56160
rect 58119 56120 58164 56148
rect 58158 56108 58164 56120
rect 58216 56108 58222 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 20898 55904 20904 55956
rect 20956 55944 20962 55956
rect 22833 55947 22891 55953
rect 22833 55944 22845 55947
rect 20956 55916 22845 55944
rect 20956 55904 20962 55916
rect 22833 55913 22845 55916
rect 22879 55944 22891 55947
rect 23658 55944 23664 55956
rect 22879 55916 23664 55944
rect 22879 55913 22891 55916
rect 22833 55907 22891 55913
rect 23658 55904 23664 55916
rect 23716 55904 23722 55956
rect 24578 55944 24584 55956
rect 24539 55916 24584 55944
rect 24578 55904 24584 55916
rect 24636 55904 24642 55956
rect 28810 55944 28816 55956
rect 24688 55916 28580 55944
rect 28771 55916 28816 55944
rect 23934 55876 23940 55888
rect 23895 55848 23940 55876
rect 23934 55836 23940 55848
rect 23992 55836 23998 55888
rect 8294 55768 8300 55820
rect 8352 55808 8358 55820
rect 24688 55808 24716 55916
rect 25222 55876 25228 55888
rect 8352 55780 24716 55808
rect 24780 55848 25228 55876
rect 8352 55768 8358 55780
rect 1857 55743 1915 55749
rect 1857 55709 1869 55743
rect 1903 55740 1915 55743
rect 1903 55712 2360 55740
rect 1903 55709 1915 55712
rect 1857 55703 1915 55709
rect 2332 55616 2360 55712
rect 20530 55700 20536 55752
rect 20588 55740 20594 55752
rect 21361 55743 21419 55749
rect 21361 55740 21373 55743
rect 20588 55712 21373 55740
rect 20588 55700 20594 55712
rect 21361 55709 21373 55712
rect 21407 55709 21419 55743
rect 23382 55740 23388 55752
rect 23343 55712 23388 55740
rect 21361 55703 21419 55709
rect 23382 55700 23388 55712
rect 23440 55700 23446 55752
rect 23566 55740 23572 55752
rect 23527 55712 23572 55740
rect 23566 55700 23572 55712
rect 23624 55700 23630 55752
rect 23658 55700 23664 55752
rect 23716 55740 23722 55752
rect 23805 55743 23863 55749
rect 23716 55712 23761 55740
rect 23716 55700 23722 55712
rect 23805 55709 23817 55743
rect 23851 55740 23863 55743
rect 24670 55740 24676 55752
rect 23851 55712 24676 55740
rect 23851 55709 23863 55712
rect 23805 55703 23863 55709
rect 24670 55700 24676 55712
rect 24728 55700 24734 55752
rect 24780 55749 24808 55848
rect 25222 55836 25228 55848
rect 25280 55836 25286 55888
rect 25406 55836 25412 55888
rect 25464 55876 25470 55888
rect 25774 55876 25780 55888
rect 25464 55848 25780 55876
rect 25464 55836 25470 55848
rect 25774 55836 25780 55848
rect 25832 55876 25838 55888
rect 26602 55876 26608 55888
rect 25832 55848 26608 55876
rect 25832 55836 25838 55848
rect 26602 55836 26608 55848
rect 26660 55836 26666 55888
rect 25038 55808 25044 55820
rect 24999 55780 25044 55808
rect 25038 55768 25044 55780
rect 25096 55768 25102 55820
rect 28350 55808 28356 55820
rect 28311 55780 28356 55808
rect 28350 55768 28356 55780
rect 28408 55768 28414 55820
rect 28552 55808 28580 55916
rect 28810 55904 28816 55916
rect 28868 55904 28874 55956
rect 28902 55904 28908 55956
rect 28960 55944 28966 55956
rect 32677 55947 32735 55953
rect 32677 55944 32689 55947
rect 28960 55916 32689 55944
rect 28960 55904 28966 55916
rect 32677 55913 32689 55916
rect 32723 55913 32735 55947
rect 32677 55907 32735 55913
rect 36078 55904 36084 55956
rect 36136 55944 36142 55956
rect 38473 55947 38531 55953
rect 38473 55944 38485 55947
rect 36136 55916 38485 55944
rect 36136 55904 36142 55916
rect 38473 55913 38485 55916
rect 38519 55913 38531 55947
rect 38473 55907 38531 55913
rect 38608 55904 38614 55956
rect 38666 55904 38672 55956
rect 40954 55904 40960 55956
rect 41012 55944 41018 55956
rect 41506 55944 41512 55956
rect 41012 55916 41512 55944
rect 41012 55904 41018 55916
rect 41506 55904 41512 55916
rect 41564 55904 41570 55956
rect 57149 55947 57207 55953
rect 57149 55913 57161 55947
rect 57195 55944 57207 55947
rect 58434 55944 58440 55956
rect 57195 55916 58440 55944
rect 57195 55913 57207 55916
rect 57149 55907 57207 55913
rect 58434 55904 58440 55916
rect 58492 55904 58498 55956
rect 30282 55876 30288 55888
rect 29012 55848 30144 55876
rect 30243 55848 30288 55876
rect 29012 55808 29040 55848
rect 28552 55780 29040 55808
rect 30116 55808 30144 55848
rect 30282 55836 30288 55848
rect 30340 55836 30346 55888
rect 31018 55836 31024 55888
rect 31076 55876 31082 55888
rect 35621 55879 35679 55885
rect 35621 55876 35633 55879
rect 31076 55848 35633 55876
rect 31076 55836 31082 55848
rect 35621 55845 35633 55848
rect 35667 55845 35679 55879
rect 37550 55876 37556 55888
rect 35621 55839 35679 55845
rect 36188 55848 37556 55876
rect 30929 55811 30987 55817
rect 30929 55808 30941 55811
rect 30116 55780 30941 55808
rect 30929 55777 30941 55780
rect 30975 55808 30987 55811
rect 31202 55808 31208 55820
rect 30975 55780 31208 55808
rect 30975 55777 30987 55780
rect 30929 55771 30987 55777
rect 31202 55768 31208 55780
rect 31260 55768 31266 55820
rect 36188 55808 36216 55848
rect 37550 55836 37556 55848
rect 37608 55836 37614 55888
rect 38286 55836 38292 55888
rect 38344 55876 38350 55888
rect 38626 55876 38654 55904
rect 41138 55876 41144 55888
rect 38344 55848 38654 55876
rect 41099 55848 41144 55876
rect 38344 55836 38350 55848
rect 41138 55836 41144 55848
rect 41196 55836 41202 55888
rect 43257 55879 43315 55885
rect 43257 55876 43269 55879
rect 41248 55848 43269 55876
rect 38838 55808 38844 55820
rect 33244 55780 36216 55808
rect 38672 55780 38844 55808
rect 24765 55743 24823 55749
rect 24765 55709 24777 55743
rect 24811 55709 24823 55743
rect 24765 55703 24823 55709
rect 24949 55743 25007 55749
rect 24949 55709 24961 55743
rect 24995 55740 25007 55743
rect 25130 55740 25136 55752
rect 24995 55712 25136 55740
rect 24995 55709 25007 55712
rect 24949 55703 25007 55709
rect 25130 55700 25136 55712
rect 25188 55740 25194 55752
rect 25774 55740 25780 55752
rect 25188 55712 25780 55740
rect 25188 55700 25194 55712
rect 25774 55700 25780 55712
rect 25832 55700 25838 55752
rect 26970 55740 26976 55752
rect 26931 55712 26976 55740
rect 26970 55700 26976 55712
rect 27028 55740 27034 55752
rect 27338 55740 27344 55752
rect 27028 55712 27344 55740
rect 27028 55700 27034 55712
rect 27338 55700 27344 55712
rect 27396 55700 27402 55752
rect 28442 55740 28448 55752
rect 28403 55712 28448 55740
rect 28442 55700 28448 55712
rect 28500 55700 28506 55752
rect 28629 55743 28687 55749
rect 28629 55709 28641 55743
rect 28675 55709 28687 55743
rect 28629 55703 28687 55709
rect 21177 55675 21235 55681
rect 21177 55641 21189 55675
rect 21223 55641 21235 55675
rect 21177 55635 21235 55641
rect 21545 55675 21603 55681
rect 21545 55641 21557 55675
rect 21591 55672 21603 55675
rect 28350 55672 28356 55684
rect 21591 55644 28356 55672
rect 21591 55641 21603 55644
rect 21545 55635 21603 55641
rect 1670 55604 1676 55616
rect 1631 55576 1676 55604
rect 1670 55564 1676 55576
rect 1728 55564 1734 55616
rect 2314 55604 2320 55616
rect 2275 55576 2320 55604
rect 2314 55564 2320 55576
rect 2372 55564 2378 55616
rect 21192 55604 21220 55635
rect 28350 55632 28356 55644
rect 28408 55632 28414 55684
rect 28644 55672 28672 55703
rect 29178 55700 29184 55752
rect 29236 55740 29242 55752
rect 29733 55743 29791 55749
rect 29733 55740 29745 55743
rect 29236 55712 29745 55740
rect 29236 55700 29242 55712
rect 29733 55709 29745 55712
rect 29779 55709 29791 55743
rect 29914 55740 29920 55752
rect 29875 55712 29920 55740
rect 29733 55703 29791 55709
rect 29914 55700 29920 55712
rect 29972 55700 29978 55752
rect 32858 55749 32864 55752
rect 30153 55743 30211 55749
rect 30153 55709 30165 55743
rect 30199 55740 30211 55743
rect 32856 55740 32864 55749
rect 30199 55712 31754 55740
rect 32819 55712 32864 55740
rect 30199 55709 30236 55712
rect 30153 55703 30236 55709
rect 29454 55672 29460 55684
rect 28644 55644 29460 55672
rect 21910 55604 21916 55616
rect 21192 55576 21916 55604
rect 21910 55564 21916 55576
rect 21968 55564 21974 55616
rect 25222 55564 25228 55616
rect 25280 55604 25286 55616
rect 25958 55604 25964 55616
rect 25280 55576 25964 55604
rect 25280 55564 25286 55576
rect 25958 55564 25964 55576
rect 26016 55604 26022 55616
rect 28644 55604 28672 55644
rect 29454 55632 29460 55644
rect 29512 55632 29518 55684
rect 30006 55672 30012 55684
rect 29967 55644 30012 55672
rect 30006 55632 30012 55644
rect 30064 55632 30070 55684
rect 26016 55576 28672 55604
rect 26016 55564 26022 55576
rect 28810 55564 28816 55616
rect 28868 55604 28874 55616
rect 30208 55604 30236 55703
rect 31726 55684 31754 55712
rect 32856 55703 32864 55712
rect 32858 55700 32864 55703
rect 32916 55700 32922 55752
rect 32950 55700 32956 55752
rect 33008 55740 33014 55752
rect 33244 55749 33272 55780
rect 33228 55743 33286 55749
rect 33008 55712 33053 55740
rect 33008 55700 33014 55712
rect 33228 55709 33240 55743
rect 33274 55709 33286 55743
rect 33228 55703 33286 55709
rect 33318 55700 33324 55752
rect 33376 55740 33382 55752
rect 33376 55712 33421 55740
rect 33376 55700 33382 55712
rect 34606 55700 34612 55752
rect 34664 55740 34670 55752
rect 35710 55740 35716 55752
rect 34664 55712 35716 55740
rect 34664 55700 34670 55712
rect 35710 55700 35716 55712
rect 35768 55749 35774 55752
rect 35768 55743 35817 55749
rect 35768 55709 35771 55743
rect 35805 55709 35817 55743
rect 35768 55703 35817 55709
rect 35768 55700 35774 55703
rect 35894 55700 35900 55752
rect 35952 55740 35958 55752
rect 36172 55743 36230 55749
rect 35952 55712 35997 55740
rect 35952 55700 35958 55712
rect 36172 55709 36184 55743
rect 36218 55709 36230 55743
rect 36172 55703 36230 55709
rect 31726 55644 31760 55684
rect 31754 55632 31760 55644
rect 31812 55632 31818 55684
rect 33045 55675 33103 55681
rect 33045 55641 33057 55675
rect 33091 55672 33103 55675
rect 35618 55672 35624 55684
rect 33091 55644 35624 55672
rect 33091 55641 33103 55644
rect 33045 55635 33103 55641
rect 35618 55632 35624 55644
rect 35676 55632 35682 55684
rect 35989 55675 36047 55681
rect 35989 55641 36001 55675
rect 36035 55641 36047 55675
rect 36188 55672 36216 55703
rect 36262 55700 36268 55752
rect 36320 55740 36326 55752
rect 36320 55712 36365 55740
rect 36320 55700 36326 55712
rect 37734 55700 37740 55752
rect 37792 55740 37798 55752
rect 38470 55740 38476 55752
rect 37792 55712 38476 55740
rect 37792 55700 37798 55712
rect 38470 55700 38476 55712
rect 38528 55700 38534 55752
rect 38672 55749 38700 55780
rect 38838 55768 38844 55780
rect 38896 55768 38902 55820
rect 41248 55808 41276 55848
rect 43257 55845 43269 55848
rect 43303 55845 43315 55879
rect 43257 55839 43315 55845
rect 52178 55808 52184 55820
rect 40972 55780 41276 55808
rect 41616 55780 52184 55808
rect 38649 55743 38707 55749
rect 38649 55709 38661 55743
rect 38695 55709 38707 55743
rect 38749 55743 38807 55749
rect 38749 55730 38761 55743
rect 38795 55730 38807 55743
rect 38933 55743 38991 55749
rect 38649 55703 38707 55709
rect 37458 55672 37464 55684
rect 36188 55644 37464 55672
rect 35989 55635 36047 55641
rect 28868 55576 30236 55604
rect 36004 55604 36032 55635
rect 37458 55632 37464 55644
rect 37516 55632 37522 55684
rect 38746 55678 38752 55730
rect 38804 55678 38810 55730
rect 38933 55709 38945 55743
rect 38979 55709 38991 55743
rect 38933 55703 38991 55709
rect 39035 55721 39093 55727
rect 38488 55644 38654 55672
rect 38488 55604 38516 55644
rect 36004 55576 38516 55604
rect 38626 55604 38654 55644
rect 38838 55632 38844 55684
rect 38896 55672 38902 55684
rect 38948 55672 38976 55703
rect 39035 55687 39047 55721
rect 39081 55687 39093 55721
rect 40494 55700 40500 55752
rect 40552 55740 40558 55752
rect 40972 55740 41000 55780
rect 40552 55712 41000 55740
rect 40552 55700 40558 55712
rect 41046 55700 41052 55752
rect 41104 55740 41110 55752
rect 41320 55743 41378 55749
rect 41320 55740 41332 55743
rect 41104 55734 41184 55740
rect 41294 55734 41332 55740
rect 41104 55712 41332 55734
rect 41104 55700 41110 55712
rect 41156 55709 41332 55712
rect 41366 55709 41378 55743
rect 41156 55706 41378 55709
rect 41320 55703 41378 55706
rect 41408 55743 41466 55749
rect 41408 55709 41420 55743
rect 41454 55740 41466 55743
rect 41616 55740 41644 55780
rect 52178 55768 52184 55780
rect 52236 55768 52242 55820
rect 41454 55712 41644 55740
rect 41692 55743 41750 55749
rect 41454 55709 41466 55712
rect 41408 55703 41466 55709
rect 41692 55709 41704 55743
rect 41738 55709 41750 55743
rect 41692 55703 41750 55709
rect 39035 55684 39093 55687
rect 38896 55644 38976 55672
rect 38896 55632 38902 55644
rect 39022 55632 39028 55684
rect 39080 55681 39093 55684
rect 39080 55632 39086 55681
rect 41506 55672 41512 55684
rect 41467 55644 41512 55672
rect 41506 55632 41512 55644
rect 41564 55632 41570 55684
rect 41708 55672 41736 55703
rect 41782 55700 41788 55752
rect 41840 55740 41846 55752
rect 41840 55712 41885 55740
rect 41840 55700 41846 55712
rect 42610 55700 42616 55752
rect 42668 55740 42674 55752
rect 43395 55743 43453 55749
rect 43395 55740 43407 55743
rect 42668 55712 43407 55740
rect 42668 55700 42674 55712
rect 43395 55709 43407 55712
rect 43441 55709 43453 55743
rect 43622 55740 43628 55752
rect 43583 55712 43628 55740
rect 43395 55703 43453 55709
rect 43622 55700 43628 55712
rect 43680 55700 43686 55752
rect 43808 55743 43866 55749
rect 43808 55709 43820 55743
rect 43854 55709 43866 55743
rect 43808 55703 43866 55709
rect 42794 55672 42800 55684
rect 41708 55644 42800 55672
rect 42794 55632 42800 55644
rect 42852 55632 42858 55684
rect 43533 55675 43591 55681
rect 43533 55641 43545 55675
rect 43579 55641 43591 55675
rect 43824 55672 43852 55703
rect 43898 55700 43904 55752
rect 43956 55740 43962 55752
rect 57701 55743 57759 55749
rect 43956 55712 44001 55740
rect 43956 55700 43962 55712
rect 57701 55709 57713 55743
rect 57747 55740 57759 55743
rect 58342 55740 58348 55752
rect 57747 55712 58348 55740
rect 57747 55709 57759 55712
rect 57701 55703 57759 55709
rect 58342 55700 58348 55712
rect 58400 55700 58406 55752
rect 44726 55672 44732 55684
rect 43824 55644 44732 55672
rect 43533 55635 43591 55641
rect 43162 55604 43168 55616
rect 38626 55576 43168 55604
rect 28868 55564 28874 55576
rect 43162 55564 43168 55576
rect 43220 55564 43226 55616
rect 43548 55604 43576 55635
rect 44726 55632 44732 55644
rect 44784 55632 44790 55684
rect 55766 55672 55772 55684
rect 45526 55644 55772 55672
rect 45526 55604 45554 55644
rect 55766 55632 55772 55644
rect 55824 55632 55830 55684
rect 43548 55576 45554 55604
rect 58161 55607 58219 55613
rect 58161 55573 58173 55607
rect 58207 55604 58219 55607
rect 59538 55604 59544 55616
rect 58207 55576 59544 55604
rect 58207 55573 58219 55576
rect 58161 55567 58219 55573
rect 59538 55564 59544 55576
rect 59596 55564 59602 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 25774 55360 25780 55412
rect 25832 55400 25838 55412
rect 28442 55400 28448 55412
rect 25832 55372 28448 55400
rect 25832 55360 25838 55372
rect 28442 55360 28448 55372
rect 28500 55400 28506 55412
rect 28994 55400 29000 55412
rect 28500 55372 29000 55400
rect 28500 55360 28506 55372
rect 28994 55360 29000 55372
rect 29052 55400 29058 55412
rect 29822 55400 29828 55412
rect 29052 55372 29828 55400
rect 29052 55360 29058 55372
rect 29822 55360 29828 55372
rect 29880 55360 29886 55412
rect 34514 55360 34520 55412
rect 34572 55400 34578 55412
rect 38286 55400 38292 55412
rect 34572 55372 38292 55400
rect 34572 55360 34578 55372
rect 38286 55360 38292 55372
rect 38344 55360 38350 55412
rect 42613 55403 42671 55409
rect 42613 55400 42625 55403
rect 38856 55372 42625 55400
rect 7006 55292 7012 55344
rect 7064 55332 7070 55344
rect 29549 55335 29607 55341
rect 29549 55332 29561 55335
rect 7064 55304 29561 55332
rect 7064 55292 7070 55304
rect 29549 55301 29561 55304
rect 29595 55332 29607 55335
rect 30006 55332 30012 55344
rect 29595 55304 30012 55332
rect 29595 55301 29607 55304
rect 29549 55295 29607 55301
rect 30006 55292 30012 55304
rect 30064 55292 30070 55344
rect 1857 55267 1915 55273
rect 1857 55233 1869 55267
rect 1903 55264 1915 55267
rect 2406 55264 2412 55276
rect 1903 55236 2412 55264
rect 1903 55233 1915 55236
rect 1857 55227 1915 55233
rect 2406 55224 2412 55236
rect 2464 55224 2470 55276
rect 20806 55224 20812 55276
rect 20864 55264 20870 55276
rect 20864 55236 21864 55264
rect 20864 55224 20870 55236
rect 21836 55196 21864 55236
rect 21910 55224 21916 55276
rect 21968 55264 21974 55276
rect 22005 55267 22063 55273
rect 22005 55264 22017 55267
rect 21968 55236 22017 55264
rect 21968 55224 21974 55236
rect 22005 55233 22017 55236
rect 22051 55233 22063 55267
rect 22189 55267 22247 55273
rect 22189 55264 22201 55267
rect 22005 55227 22063 55233
rect 22112 55236 22201 55264
rect 22112 55196 22140 55236
rect 22189 55233 22201 55236
rect 22235 55233 22247 55267
rect 22189 55227 22247 55233
rect 22373 55267 22431 55273
rect 22373 55233 22385 55267
rect 22419 55264 22431 55267
rect 26050 55264 26056 55276
rect 22419 55236 26056 55264
rect 22419 55233 22431 55236
rect 22373 55227 22431 55233
rect 26050 55224 26056 55236
rect 26108 55224 26114 55276
rect 26602 55224 26608 55276
rect 26660 55264 26666 55276
rect 28534 55264 28540 55276
rect 26660 55236 28540 55264
rect 26660 55224 26666 55236
rect 28534 55224 28540 55236
rect 28592 55224 28598 55276
rect 38473 55267 38531 55273
rect 38473 55233 38485 55267
rect 38519 55264 38531 55267
rect 38746 55264 38752 55276
rect 38519 55236 38752 55264
rect 38519 55233 38531 55236
rect 38473 55227 38531 55233
rect 38746 55224 38752 55236
rect 38804 55224 38810 55276
rect 21836 55168 22140 55196
rect 35618 55156 35624 55208
rect 35676 55196 35682 55208
rect 38856 55196 38884 55372
rect 42613 55369 42625 55372
rect 42659 55369 42671 55403
rect 43346 55400 43352 55412
rect 42613 55363 42671 55369
rect 42812 55372 43352 55400
rect 40310 55292 40316 55344
rect 40368 55332 40374 55344
rect 41230 55332 41236 55344
rect 40368 55304 41236 55332
rect 40368 55292 40374 55304
rect 41230 55292 41236 55304
rect 41288 55332 41294 55344
rect 41782 55332 41788 55344
rect 41288 55304 41788 55332
rect 41288 55292 41294 55304
rect 41782 55292 41788 55304
rect 41840 55332 41846 55344
rect 42812 55332 42840 55372
rect 43346 55360 43352 55372
rect 43404 55400 43410 55412
rect 43898 55400 43904 55412
rect 43404 55372 43904 55400
rect 43404 55360 43410 55372
rect 43898 55360 43904 55372
rect 43956 55360 43962 55412
rect 56686 55360 56692 55412
rect 56744 55400 56750 55412
rect 58161 55403 58219 55409
rect 58161 55400 58173 55403
rect 56744 55372 58173 55400
rect 56744 55360 56750 55372
rect 58161 55369 58173 55372
rect 58207 55369 58219 55403
rect 58161 55363 58219 55369
rect 41840 55304 42840 55332
rect 42889 55335 42947 55341
rect 41840 55292 41846 55304
rect 42889 55301 42901 55335
rect 42935 55332 42947 55335
rect 54570 55332 54576 55344
rect 42935 55304 54576 55332
rect 42935 55301 42947 55304
rect 42889 55295 42947 55301
rect 54570 55292 54576 55304
rect 54628 55292 54634 55344
rect 39574 55264 39580 55276
rect 39535 55236 39580 55264
rect 39574 55224 39580 55236
rect 39632 55224 39638 55276
rect 40862 55224 40868 55276
rect 40920 55264 40926 55276
rect 42610 55264 42616 55276
rect 40920 55236 42616 55264
rect 40920 55224 40926 55236
rect 42610 55224 42616 55236
rect 42668 55264 42674 55276
rect 42751 55267 42809 55273
rect 42751 55264 42763 55267
rect 42668 55236 42763 55264
rect 42668 55224 42674 55236
rect 42751 55233 42763 55236
rect 42797 55233 42809 55267
rect 42978 55264 42984 55276
rect 42891 55236 42984 55264
rect 42751 55227 42809 55233
rect 42978 55224 42984 55236
rect 43036 55224 43042 55276
rect 43164 55267 43222 55273
rect 43164 55264 43176 55267
rect 43143 55236 43176 55264
rect 43164 55233 43176 55236
rect 43210 55233 43222 55267
rect 43164 55227 43222 55233
rect 43257 55267 43315 55273
rect 43257 55233 43269 55267
rect 43303 55264 43315 55267
rect 43346 55264 43352 55276
rect 43303 55236 43352 55264
rect 43303 55233 43315 55236
rect 43257 55227 43315 55233
rect 35676 55168 38884 55196
rect 35676 55156 35682 55168
rect 41506 55156 41512 55208
rect 41564 55196 41570 55208
rect 42996 55196 43024 55224
rect 41564 55168 43024 55196
rect 43180 55196 43208 55227
rect 43346 55224 43352 55236
rect 43404 55224 43410 55276
rect 44542 55264 44548 55276
rect 43456 55236 44548 55264
rect 43456 55196 43484 55236
rect 44542 55224 44548 55236
rect 44600 55224 44606 55276
rect 57517 55267 57575 55273
rect 57517 55233 57529 55267
rect 57563 55264 57575 55267
rect 57974 55264 57980 55276
rect 57563 55236 57980 55264
rect 57563 55233 57575 55236
rect 57517 55227 57575 55233
rect 57974 55224 57980 55236
rect 58032 55264 58038 55276
rect 58345 55267 58403 55273
rect 58345 55264 58357 55267
rect 58032 55236 58357 55264
rect 58032 55224 58038 55236
rect 58345 55233 58357 55236
rect 58391 55233 58403 55267
rect 58345 55227 58403 55233
rect 43180 55168 43484 55196
rect 41564 55156 41570 55168
rect 1670 55060 1676 55072
rect 1631 55032 1676 55060
rect 1670 55020 1676 55032
rect 1728 55020 1734 55072
rect 32398 55060 32404 55072
rect 32359 55032 32404 55060
rect 32398 55020 32404 55032
rect 32456 55020 32462 55072
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 25774 54816 25780 54868
rect 25832 54856 25838 54868
rect 26053 54859 26111 54865
rect 26053 54856 26065 54859
rect 25832 54828 26065 54856
rect 25832 54816 25838 54828
rect 26053 54825 26065 54828
rect 26099 54825 26111 54859
rect 26053 54819 26111 54825
rect 32769 54859 32827 54865
rect 32769 54825 32781 54859
rect 32815 54825 32827 54859
rect 32769 54819 32827 54825
rect 32490 54788 32496 54800
rect 22066 54760 32496 54788
rect 19334 54612 19340 54664
rect 19392 54652 19398 54664
rect 21821 54655 21879 54661
rect 21821 54652 21833 54655
rect 19392 54624 21833 54652
rect 19392 54612 19398 54624
rect 21821 54621 21833 54624
rect 21867 54621 21879 54655
rect 21821 54615 21879 54621
rect 21637 54587 21695 54593
rect 21637 54553 21649 54587
rect 21683 54584 21695 54587
rect 21910 54584 21916 54596
rect 21683 54556 21916 54584
rect 21683 54553 21695 54556
rect 21637 54547 21695 54553
rect 21910 54544 21916 54556
rect 21968 54584 21974 54596
rect 22066 54584 22094 54760
rect 32490 54748 32496 54760
rect 32548 54748 32554 54800
rect 25685 54723 25743 54729
rect 25685 54689 25697 54723
rect 25731 54720 25743 54723
rect 31386 54720 31392 54732
rect 25731 54692 26740 54720
rect 25731 54689 25743 54692
rect 25685 54683 25743 54689
rect 25869 54655 25927 54661
rect 25869 54621 25881 54655
rect 25915 54652 25927 54655
rect 25958 54652 25964 54664
rect 25915 54624 25964 54652
rect 25915 54621 25927 54624
rect 25869 54615 25927 54621
rect 25958 54612 25964 54624
rect 26016 54612 26022 54664
rect 26142 54612 26148 54664
rect 26200 54652 26206 54664
rect 26602 54652 26608 54664
rect 26200 54624 26245 54652
rect 26563 54624 26608 54652
rect 26200 54612 26206 54624
rect 26602 54612 26608 54624
rect 26660 54612 26666 54664
rect 26712 54661 26740 54692
rect 26896 54692 31392 54720
rect 26896 54661 26924 54692
rect 31386 54680 31392 54692
rect 31444 54680 31450 54732
rect 32784 54720 32812 54819
rect 32858 54816 32864 54868
rect 32916 54856 32922 54868
rect 32953 54859 33011 54865
rect 32953 54856 32965 54859
rect 32916 54828 32965 54856
rect 32916 54816 32922 54828
rect 32953 54825 32965 54828
rect 32999 54856 33011 54859
rect 34606 54856 34612 54868
rect 32999 54828 34612 54856
rect 32999 54825 33011 54828
rect 32953 54819 33011 54825
rect 34606 54816 34612 54828
rect 34664 54816 34670 54868
rect 37458 54856 37464 54868
rect 37419 54828 37464 54856
rect 37458 54816 37464 54828
rect 37516 54816 37522 54868
rect 31864 54692 32812 54720
rect 26698 54655 26756 54661
rect 26698 54621 26710 54655
rect 26744 54621 26756 54655
rect 26698 54615 26756 54621
rect 26881 54655 26939 54661
rect 26881 54621 26893 54655
rect 26927 54621 26939 54655
rect 26881 54615 26939 54621
rect 27070 54655 27128 54661
rect 27070 54621 27082 54655
rect 27116 54621 27128 54655
rect 27070 54615 27128 54621
rect 21968 54556 22094 54584
rect 21968 54544 21974 54556
rect 26234 54544 26240 54596
rect 26292 54584 26298 54596
rect 26973 54587 27031 54593
rect 26973 54584 26985 54587
rect 26292 54556 26985 54584
rect 26292 54544 26298 54556
rect 26973 54553 26985 54556
rect 27019 54553 27031 54587
rect 26973 54547 27031 54553
rect 27080 54584 27108 54615
rect 27430 54584 27436 54596
rect 27080 54556 27436 54584
rect 22005 54519 22063 54525
rect 22005 54485 22017 54519
rect 22051 54516 22063 54519
rect 22922 54516 22928 54528
rect 22051 54488 22928 54516
rect 22051 54485 22063 54488
rect 22005 54479 22063 54485
rect 22922 54476 22928 54488
rect 22980 54476 22986 54528
rect 23750 54476 23756 54528
rect 23808 54516 23814 54528
rect 24394 54516 24400 54528
rect 23808 54488 24400 54516
rect 23808 54476 23814 54488
rect 24394 54476 24400 54488
rect 24452 54516 24458 54528
rect 27080 54516 27108 54556
rect 27430 54544 27436 54556
rect 27488 54544 27494 54596
rect 31864 54528 31892 54692
rect 34698 54680 34704 54732
rect 34756 54720 34762 54732
rect 36909 54723 36967 54729
rect 36909 54720 36921 54723
rect 34756 54692 36921 54720
rect 34756 54680 34762 54692
rect 36909 54689 36921 54692
rect 36955 54720 36967 54723
rect 37550 54720 37556 54732
rect 36955 54692 37556 54720
rect 36955 54689 36967 54692
rect 36909 54683 36967 54689
rect 37550 54680 37556 54692
rect 37608 54680 37614 54732
rect 38378 54720 38384 54732
rect 37660 54692 38384 54720
rect 32398 54652 32404 54664
rect 32359 54624 32404 54652
rect 32398 54612 32404 54624
rect 32456 54612 32462 54664
rect 34606 54612 34612 54664
rect 34664 54652 34670 54664
rect 35023 54655 35081 54661
rect 35023 54652 35035 54655
rect 34664 54624 35035 54652
rect 34664 54612 34670 54624
rect 35023 54621 35035 54624
rect 35069 54621 35081 54655
rect 35434 54652 35440 54664
rect 35395 54624 35440 54652
rect 35023 54615 35081 54621
rect 35434 54612 35440 54624
rect 35492 54612 35498 54664
rect 35526 54612 35532 54664
rect 35584 54652 35590 54664
rect 37660 54661 37688 54692
rect 38378 54680 38384 54692
rect 38436 54680 38442 54732
rect 37645 54655 37703 54661
rect 35584 54624 35629 54652
rect 35584 54612 35590 54624
rect 37645 54621 37657 54655
rect 37691 54621 37703 54655
rect 37645 54615 37703 54621
rect 37737 54655 37795 54661
rect 37737 54621 37749 54655
rect 37783 54621 37795 54655
rect 37918 54652 37924 54664
rect 37879 54624 37924 54652
rect 37737 54615 37795 54621
rect 33226 54544 33232 54596
rect 33284 54584 33290 54596
rect 35161 54587 35219 54593
rect 35161 54584 35173 54587
rect 33284 54556 35173 54584
rect 33284 54544 33290 54556
rect 35161 54553 35173 54556
rect 35207 54553 35219 54587
rect 35161 54547 35219 54553
rect 35253 54587 35311 54593
rect 35253 54553 35265 54587
rect 35299 54584 35311 54587
rect 35618 54584 35624 54596
rect 35299 54556 35624 54584
rect 35299 54553 35311 54556
rect 35253 54547 35311 54553
rect 35618 54544 35624 54556
rect 35676 54544 35682 54596
rect 37550 54544 37556 54596
rect 37608 54584 37614 54596
rect 37752 54584 37780 54615
rect 37918 54612 37924 54624
rect 37976 54612 37982 54664
rect 38010 54612 38016 54664
rect 38068 54652 38074 54664
rect 38654 54652 38660 54664
rect 38068 54624 38113 54652
rect 38615 54624 38660 54652
rect 38068 54612 38074 54624
rect 38654 54612 38660 54624
rect 38712 54652 38718 54664
rect 39301 54655 39359 54661
rect 39301 54652 39313 54655
rect 38712 54624 39313 54652
rect 38712 54612 38718 54624
rect 39301 54621 39313 54624
rect 39347 54652 39359 54655
rect 40589 54655 40647 54661
rect 40589 54652 40601 54655
rect 39347 54624 40601 54652
rect 39347 54621 39359 54624
rect 39301 54615 39359 54621
rect 40589 54621 40601 54624
rect 40635 54621 40647 54655
rect 40589 54615 40647 54621
rect 39574 54584 39580 54596
rect 37608 54556 39580 54584
rect 37608 54544 37614 54556
rect 39574 54544 39580 54556
rect 39632 54544 39638 54596
rect 24452 54488 27108 54516
rect 27249 54519 27307 54525
rect 24452 54476 24458 54488
rect 27249 54485 27261 54519
rect 27295 54516 27307 54519
rect 27338 54516 27344 54528
rect 27295 54488 27344 54516
rect 27295 54485 27307 54488
rect 27249 54479 27307 54485
rect 27338 54476 27344 54488
rect 27396 54476 27402 54528
rect 31846 54516 31852 54528
rect 31807 54488 31852 54516
rect 31846 54476 31852 54488
rect 31904 54476 31910 54528
rect 32766 54516 32772 54528
rect 32727 54488 32772 54516
rect 32766 54476 32772 54488
rect 32824 54476 32830 54528
rect 34882 54516 34888 54528
rect 34843 54488 34888 54516
rect 34882 54476 34888 54488
rect 34940 54476 34946 54528
rect 37918 54476 37924 54528
rect 37976 54516 37982 54528
rect 38749 54519 38807 54525
rect 38749 54516 38761 54519
rect 37976 54488 38761 54516
rect 37976 54476 37982 54488
rect 38749 54485 38761 54488
rect 38795 54516 38807 54519
rect 38930 54516 38936 54528
rect 38795 54488 38936 54516
rect 38795 54485 38807 54488
rect 38749 54479 38807 54485
rect 38930 54476 38936 54488
rect 38988 54476 38994 54528
rect 39666 54476 39672 54528
rect 39724 54516 39730 54528
rect 40037 54519 40095 54525
rect 40037 54516 40049 54519
rect 39724 54488 40049 54516
rect 39724 54476 39730 54488
rect 40037 54485 40049 54488
rect 40083 54485 40095 54519
rect 58342 54516 58348 54528
rect 58303 54488 58348 54516
rect 40037 54479 40095 54485
rect 58342 54476 58348 54488
rect 58400 54476 58406 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 26513 54315 26571 54321
rect 26513 54312 26525 54315
rect 6886 54284 26525 54312
rect 1857 54179 1915 54185
rect 1857 54145 1869 54179
rect 1903 54176 1915 54179
rect 1903 54148 2452 54176
rect 1903 54145 1915 54148
rect 1857 54139 1915 54145
rect 1670 54040 1676 54052
rect 1631 54012 1676 54040
rect 1670 54000 1676 54012
rect 1728 54000 1734 54052
rect 2424 53981 2452 54148
rect 2409 53975 2467 53981
rect 2409 53941 2421 53975
rect 2455 53972 2467 53975
rect 2866 53972 2872 53984
rect 2455 53944 2872 53972
rect 2455 53941 2467 53944
rect 2409 53935 2467 53941
rect 2866 53932 2872 53944
rect 2924 53932 2930 53984
rect 5718 53932 5724 53984
rect 5776 53972 5782 53984
rect 6886 53972 6914 54284
rect 26513 54281 26525 54284
rect 26559 54312 26571 54315
rect 27726 54315 27784 54321
rect 26559 54284 27476 54312
rect 26559 54281 26571 54284
rect 26513 54275 26571 54281
rect 18874 54204 18880 54256
rect 18932 54244 18938 54256
rect 24489 54247 24547 54253
rect 24489 54244 24501 54247
rect 18932 54216 24501 54244
rect 18932 54204 18938 54216
rect 24489 54213 24501 54216
rect 24535 54213 24547 54247
rect 25317 54247 25375 54253
rect 25317 54244 25329 54247
rect 24489 54207 24547 54213
rect 24780 54216 25329 54244
rect 24394 54185 24400 54188
rect 24392 54176 24400 54185
rect 24355 54148 24400 54176
rect 24392 54139 24400 54148
rect 24394 54136 24400 54139
rect 24452 54136 24458 54188
rect 24780 54185 24808 54216
rect 25317 54213 25329 54216
rect 25363 54213 25375 54247
rect 25958 54244 25964 54256
rect 25317 54207 25375 54213
rect 25516 54216 25964 54244
rect 24581 54179 24639 54185
rect 24581 54145 24593 54179
rect 24627 54145 24639 54179
rect 24581 54139 24639 54145
rect 24764 54179 24822 54185
rect 24764 54145 24776 54179
rect 24810 54145 24822 54179
rect 24764 54139 24822 54145
rect 24857 54179 24915 54185
rect 24857 54145 24869 54179
rect 24903 54176 24915 54179
rect 25406 54176 25412 54188
rect 24903 54148 25412 54176
rect 24903 54145 24915 54148
rect 24857 54139 24915 54145
rect 24596 54040 24624 54139
rect 25406 54136 25412 54148
rect 25464 54136 25470 54188
rect 25516 54185 25544 54216
rect 25958 54204 25964 54216
rect 26016 54204 26022 54256
rect 27338 54244 27344 54256
rect 27299 54216 27344 54244
rect 27338 54204 27344 54216
rect 27396 54204 27402 54256
rect 27448 54253 27476 54284
rect 27726 54281 27738 54315
rect 27772 54312 27784 54315
rect 30926 54312 30932 54324
rect 27772 54284 30932 54312
rect 27772 54281 27784 54284
rect 27726 54275 27784 54281
rect 30926 54272 30932 54284
rect 30984 54272 30990 54324
rect 31757 54315 31815 54321
rect 31757 54281 31769 54315
rect 31803 54312 31815 54315
rect 31846 54312 31852 54324
rect 31803 54284 31852 54312
rect 31803 54281 31815 54284
rect 31757 54275 31815 54281
rect 31846 54272 31852 54284
rect 31904 54272 31910 54324
rect 32490 54312 32496 54324
rect 32451 54284 32496 54312
rect 32490 54272 32496 54284
rect 32548 54272 32554 54324
rect 34517 54315 34575 54321
rect 34517 54281 34529 54315
rect 34563 54312 34575 54315
rect 35342 54312 35348 54324
rect 34563 54284 35348 54312
rect 34563 54281 34575 54284
rect 34517 54275 34575 54281
rect 35342 54272 35348 54284
rect 35400 54272 35406 54324
rect 35434 54272 35440 54324
rect 35492 54312 35498 54324
rect 36265 54315 36323 54321
rect 36265 54312 36277 54315
rect 35492 54284 36277 54312
rect 35492 54272 35498 54284
rect 36265 54281 36277 54284
rect 36311 54281 36323 54315
rect 36265 54275 36323 54281
rect 38010 54272 38016 54324
rect 38068 54312 38074 54324
rect 38933 54315 38991 54321
rect 38933 54312 38945 54315
rect 38068 54284 38945 54312
rect 38068 54272 38074 54284
rect 38933 54281 38945 54284
rect 38979 54312 38991 54315
rect 39022 54312 39028 54324
rect 38979 54284 39028 54312
rect 38979 54281 38991 54284
rect 38933 54275 38991 54281
rect 39022 54272 39028 54284
rect 39080 54272 39086 54324
rect 40310 54312 40316 54324
rect 40271 54284 40316 54312
rect 40310 54272 40316 54284
rect 40368 54272 40374 54324
rect 40862 54272 40868 54324
rect 40920 54312 40926 54324
rect 41141 54315 41199 54321
rect 41141 54312 41153 54315
rect 40920 54284 41153 54312
rect 40920 54272 40926 54284
rect 41141 54281 41153 54284
rect 41187 54281 41199 54315
rect 41141 54275 41199 54281
rect 27433 54247 27491 54253
rect 27433 54213 27445 54247
rect 27479 54213 27491 54247
rect 27433 54207 27491 54213
rect 32306 54204 32312 54256
rect 32364 54244 32370 54256
rect 32582 54244 32588 54256
rect 32364 54216 32588 54244
rect 32364 54204 32370 54216
rect 32582 54204 32588 54216
rect 32640 54204 32646 54256
rect 34885 54247 34943 54253
rect 34655 54213 34713 54219
rect 25501 54179 25559 54185
rect 25501 54145 25513 54179
rect 25547 54145 25559 54179
rect 25682 54176 25688 54188
rect 25643 54148 25688 54176
rect 25501 54139 25559 54145
rect 25682 54136 25688 54148
rect 25740 54136 25746 54188
rect 25777 54179 25835 54185
rect 25777 54145 25789 54179
rect 25823 54176 25835 54179
rect 25866 54176 25872 54188
rect 25823 54148 25872 54176
rect 25823 54145 25835 54148
rect 25777 54139 25835 54145
rect 25866 54136 25872 54148
rect 25924 54136 25930 54188
rect 26050 54136 26056 54188
rect 26108 54176 26114 54188
rect 27157 54179 27215 54185
rect 27157 54176 27169 54179
rect 26108 54148 27169 54176
rect 26108 54136 26114 54148
rect 27157 54145 27169 54148
rect 27203 54145 27215 54179
rect 27522 54176 27528 54188
rect 27580 54185 27586 54188
rect 27440 54148 27528 54176
rect 27157 54139 27215 54145
rect 27522 54136 27528 54148
rect 27580 54139 27588 54185
rect 30193 54179 30251 54185
rect 30193 54145 30205 54179
rect 30239 54176 30251 54179
rect 30558 54176 30564 54188
rect 30239 54148 30564 54176
rect 30239 54145 30251 54148
rect 30193 54139 30251 54145
rect 27580 54136 27586 54139
rect 30558 54136 30564 54148
rect 30616 54136 30622 54188
rect 32674 54176 32680 54188
rect 31864 54148 32680 54176
rect 24670 54068 24676 54120
rect 24728 54108 24734 54120
rect 27545 54108 27573 54136
rect 31864 54120 31892 54148
rect 32674 54136 32680 54148
rect 32732 54136 32738 54188
rect 34655 54179 34667 54213
rect 34701 54188 34713 54213
rect 34885 54213 34897 54247
rect 34931 54244 34943 54247
rect 37918 54244 37924 54256
rect 34931 54216 37924 54244
rect 34931 54213 34943 54216
rect 34885 54207 34943 54213
rect 35360 54188 35388 54216
rect 34701 54179 34704 54188
rect 34655 54176 34704 54179
rect 33980 54148 34704 54176
rect 24728 54080 27573 54108
rect 29273 54111 29331 54117
rect 24728 54068 24734 54080
rect 29273 54077 29285 54111
rect 29319 54108 29331 54111
rect 29730 54108 29736 54120
rect 29319 54080 29736 54108
rect 29319 54077 29331 54080
rect 29273 54071 29331 54077
rect 29730 54068 29736 54080
rect 29788 54108 29794 54120
rect 30101 54111 30159 54117
rect 30101 54108 30113 54111
rect 29788 54080 30113 54108
rect 29788 54068 29794 54080
rect 30101 54077 30113 54080
rect 30147 54108 30159 54111
rect 31846 54108 31852 54120
rect 30147 54080 31852 54108
rect 30147 54077 30159 54080
rect 30101 54071 30159 54077
rect 31846 54068 31852 54080
rect 31904 54068 31910 54120
rect 32306 54108 32312 54120
rect 32267 54080 32312 54108
rect 32306 54068 32312 54080
rect 32364 54068 32370 54120
rect 32398 54068 32404 54120
rect 32456 54108 32462 54120
rect 33980 54117 34008 54148
rect 34698 54136 34704 54148
rect 34756 54176 34762 54188
rect 34756 54148 34817 54176
rect 34756 54136 34762 54148
rect 35342 54136 35348 54188
rect 35400 54136 35406 54188
rect 36538 54185 36544 54188
rect 36441 54169 36499 54175
rect 36441 54135 36453 54169
rect 36487 54135 36499 54169
rect 36533 54139 36544 54185
rect 36596 54176 36602 54188
rect 36740 54185 36768 54216
rect 37918 54204 37924 54216
rect 37976 54204 37982 54256
rect 36725 54179 36783 54185
rect 36596 54148 36633 54176
rect 36538 54136 36544 54139
rect 36596 54136 36602 54148
rect 36725 54145 36737 54179
rect 36771 54145 36783 54179
rect 36725 54139 36783 54145
rect 36814 54136 36820 54188
rect 36872 54176 36878 54188
rect 38028 54176 38056 54272
rect 38654 54204 38660 54256
rect 38712 54244 38718 54256
rect 40129 54247 40187 54253
rect 40129 54244 40141 54247
rect 38712 54216 40141 54244
rect 38712 54204 38718 54216
rect 40129 54213 40141 54216
rect 40175 54244 40187 54247
rect 40773 54247 40831 54253
rect 40773 54244 40785 54247
rect 40175 54216 40785 54244
rect 40175 54213 40187 54216
rect 40129 54207 40187 54213
rect 40773 54213 40785 54216
rect 40819 54213 40831 54247
rect 40973 54247 41031 54253
rect 40973 54244 40985 54247
rect 40773 54207 40831 54213
rect 40880 54216 40985 54244
rect 36872 54148 38056 54176
rect 38289 54179 38347 54185
rect 36872 54136 36878 54148
rect 38289 54145 38301 54179
rect 38335 54176 38347 54179
rect 38841 54179 38899 54185
rect 38841 54176 38853 54179
rect 38335 54148 38853 54176
rect 38335 54145 38347 54148
rect 38289 54139 38347 54145
rect 38841 54145 38853 54148
rect 38887 54176 38899 54179
rect 39666 54176 39672 54188
rect 38887 54148 39672 54176
rect 38887 54145 38899 54148
rect 38841 54139 38899 54145
rect 39666 54136 39672 54148
rect 39724 54136 39730 54188
rect 36441 54129 36499 54135
rect 33965 54111 34023 54117
rect 33965 54108 33977 54111
rect 32456 54080 33977 54108
rect 32456 54068 32462 54080
rect 33965 54077 33977 54080
rect 34011 54077 34023 54111
rect 33965 54071 34023 54077
rect 36464 54052 36492 54129
rect 39574 54068 39580 54120
rect 39632 54108 39638 54120
rect 40880 54108 40908 54216
rect 40973 54213 40985 54216
rect 41019 54244 41031 54247
rect 41601 54247 41659 54253
rect 41601 54244 41613 54247
rect 41019 54216 41613 54244
rect 41019 54213 41031 54216
rect 40973 54207 41031 54213
rect 41601 54213 41613 54216
rect 41647 54213 41659 54247
rect 41601 54207 41659 54213
rect 58342 54176 58348 54188
rect 58303 54148 58348 54176
rect 58342 54136 58348 54148
rect 58400 54136 58406 54188
rect 39632 54080 40908 54108
rect 39632 54068 39638 54080
rect 34882 54040 34888 54052
rect 24596 54012 34888 54040
rect 34882 54000 34888 54012
rect 34940 54000 34946 54052
rect 36446 54000 36452 54052
rect 36504 54000 36510 54052
rect 39666 54000 39672 54052
rect 39724 54040 39730 54052
rect 39761 54043 39819 54049
rect 39761 54040 39773 54043
rect 39724 54012 39773 54040
rect 39724 54000 39730 54012
rect 39761 54009 39773 54012
rect 39807 54040 39819 54043
rect 39807 54012 41000 54040
rect 39807 54009 39819 54012
rect 39761 54003 39819 54009
rect 5776 53944 6914 53972
rect 24213 53975 24271 53981
rect 5776 53932 5782 53944
rect 24213 53941 24225 53975
rect 24259 53972 24271 53975
rect 24762 53972 24768 53984
rect 24259 53944 24768 53972
rect 24259 53941 24271 53944
rect 24213 53935 24271 53941
rect 24762 53932 24768 53944
rect 24820 53932 24826 53984
rect 29454 53932 29460 53984
rect 29512 53972 29518 53984
rect 29825 53975 29883 53981
rect 29825 53972 29837 53975
rect 29512 53944 29837 53972
rect 29512 53932 29518 53944
rect 29825 53941 29837 53944
rect 29871 53941 29883 53975
rect 29825 53935 29883 53941
rect 29914 53932 29920 53984
rect 29972 53972 29978 53984
rect 30009 53975 30067 53981
rect 30009 53972 30021 53975
rect 29972 53944 30021 53972
rect 29972 53932 29978 53944
rect 30009 53941 30021 53944
rect 30055 53941 30067 53975
rect 30009 53935 30067 53941
rect 32306 53932 32312 53984
rect 32364 53972 32370 53984
rect 32861 53975 32919 53981
rect 32861 53972 32873 53975
rect 32364 53944 32873 53972
rect 32364 53932 32370 53944
rect 32861 53941 32873 53944
rect 32907 53972 32919 53975
rect 34701 53975 34759 53981
rect 34701 53972 34713 53975
rect 32907 53944 34713 53972
rect 32907 53941 32919 53944
rect 32861 53935 32919 53941
rect 34701 53941 34713 53944
rect 34747 53972 34759 53975
rect 36814 53972 36820 53984
rect 34747 53944 36820 53972
rect 34747 53941 34759 53944
rect 34701 53935 34759 53941
rect 36814 53932 36820 53944
rect 36872 53932 36878 53984
rect 39574 53932 39580 53984
rect 39632 53972 39638 53984
rect 40972 53981 41000 54012
rect 40129 53975 40187 53981
rect 40129 53972 40141 53975
rect 39632 53944 40141 53972
rect 39632 53932 39638 53944
rect 40129 53941 40141 53944
rect 40175 53941 40187 53975
rect 40129 53935 40187 53941
rect 40957 53975 41015 53981
rect 40957 53941 40969 53975
rect 41003 53941 41015 53975
rect 40957 53935 41015 53941
rect 58161 53975 58219 53981
rect 58161 53941 58173 53975
rect 58207 53972 58219 53975
rect 58894 53972 58900 53984
rect 58207 53944 58900 53972
rect 58207 53941 58219 53944
rect 58161 53935 58219 53941
rect 58894 53932 58900 53944
rect 58952 53932 58958 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 30834 53728 30840 53780
rect 30892 53768 30898 53780
rect 31481 53771 31539 53777
rect 31481 53768 31493 53771
rect 30892 53740 31493 53768
rect 30892 53728 30898 53740
rect 31481 53737 31493 53740
rect 31527 53737 31539 53771
rect 31481 53731 31539 53737
rect 31665 53771 31723 53777
rect 31665 53737 31677 53771
rect 31711 53737 31723 53771
rect 31665 53731 31723 53737
rect 25133 53703 25191 53709
rect 25133 53669 25145 53703
rect 25179 53700 25191 53703
rect 29822 53700 29828 53712
rect 25179 53672 29828 53700
rect 25179 53669 25191 53672
rect 25133 53663 25191 53669
rect 29822 53660 29828 53672
rect 29880 53660 29886 53712
rect 30466 53700 30472 53712
rect 30427 53672 30472 53700
rect 30466 53660 30472 53672
rect 30524 53660 30530 53712
rect 24670 53592 24676 53644
rect 24728 53632 24734 53644
rect 31680 53632 31708 53731
rect 31754 53728 31760 53780
rect 31812 53768 31818 53780
rect 32309 53771 32367 53777
rect 32309 53768 32321 53771
rect 31812 53740 32321 53768
rect 31812 53728 31818 53740
rect 32309 53737 32321 53740
rect 32355 53737 32367 53771
rect 37550 53768 37556 53780
rect 37511 53740 37556 53768
rect 32309 53731 32367 53737
rect 37550 53728 37556 53740
rect 37608 53728 37614 53780
rect 38470 53768 38476 53780
rect 38431 53740 38476 53768
rect 38470 53728 38476 53740
rect 38528 53728 38534 53780
rect 39666 53728 39672 53780
rect 39724 53768 39730 53780
rect 40405 53771 40463 53777
rect 40405 53768 40417 53771
rect 39724 53740 40417 53768
rect 39724 53728 39730 53740
rect 40405 53737 40417 53740
rect 40451 53737 40463 53771
rect 40405 53731 40463 53737
rect 40589 53771 40647 53777
rect 40589 53737 40601 53771
rect 40635 53768 40647 53771
rect 41506 53768 41512 53780
rect 40635 53740 41512 53768
rect 40635 53737 40647 53740
rect 40589 53731 40647 53737
rect 32582 53660 32588 53712
rect 32640 53700 32646 53712
rect 32640 53672 32899 53700
rect 32640 53660 32646 53672
rect 32766 53632 32772 53644
rect 24728 53604 24900 53632
rect 24728 53592 24734 53604
rect 1857 53567 1915 53573
rect 1857 53533 1869 53567
rect 1903 53564 1915 53567
rect 1903 53536 2452 53564
rect 1903 53533 1915 53536
rect 1857 53527 1915 53533
rect 1670 53428 1676 53440
rect 1631 53400 1676 53428
rect 1670 53388 1676 53400
rect 1728 53388 1734 53440
rect 2424 53437 2452 53536
rect 22922 53524 22928 53576
rect 22980 53564 22986 53576
rect 24581 53567 24639 53573
rect 24581 53564 24593 53567
rect 22980 53536 24593 53564
rect 22980 53524 22986 53536
rect 24581 53533 24593 53536
rect 24627 53533 24639 53567
rect 24762 53564 24768 53576
rect 24723 53536 24768 53564
rect 24581 53527 24639 53533
rect 24762 53524 24768 53536
rect 24820 53524 24826 53576
rect 24872 53564 24900 53604
rect 30208 53604 32772 53632
rect 24954 53567 25012 53573
rect 24954 53564 24966 53567
rect 24872 53536 24966 53564
rect 24954 53533 24966 53536
rect 25000 53533 25012 53567
rect 24954 53527 25012 53533
rect 29181 53567 29239 53573
rect 29181 53533 29193 53567
rect 29227 53564 29239 53567
rect 29730 53564 29736 53576
rect 29227 53536 29736 53564
rect 29227 53533 29239 53536
rect 29181 53527 29239 53533
rect 29730 53524 29736 53536
rect 29788 53524 29794 53576
rect 29914 53524 29920 53576
rect 29972 53564 29978 53576
rect 30208 53573 30236 53604
rect 32766 53592 32772 53604
rect 32824 53592 32830 53644
rect 32871 53632 32899 53672
rect 36538 53660 36544 53712
rect 36596 53700 36602 53712
rect 38488 53700 38516 53728
rect 36596 53672 38516 53700
rect 36596 53660 36602 53672
rect 39574 53660 39580 53712
rect 39632 53700 39638 53712
rect 40037 53703 40095 53709
rect 40037 53700 40049 53703
rect 39632 53672 40049 53700
rect 39632 53660 39638 53672
rect 40037 53669 40049 53672
rect 40083 53669 40095 53703
rect 40420 53700 40448 53731
rect 41506 53728 41512 53740
rect 41564 53728 41570 53780
rect 41049 53703 41107 53709
rect 41049 53700 41061 53703
rect 40420 53672 41061 53700
rect 40037 53663 40095 53669
rect 41049 53669 41061 53672
rect 41095 53669 41107 53703
rect 41049 53663 41107 53669
rect 36556 53632 36584 53660
rect 32871 53604 36584 53632
rect 30193 53567 30251 53573
rect 30193 53564 30205 53567
rect 29972 53536 30205 53564
rect 29972 53524 29978 53536
rect 30193 53533 30205 53536
rect 30239 53533 30251 53567
rect 30558 53564 30564 53576
rect 30471 53536 30564 53564
rect 30193 53527 30251 53533
rect 30558 53524 30564 53536
rect 30616 53564 30622 53576
rect 30616 53536 31708 53564
rect 30616 53524 30622 53536
rect 24857 53499 24915 53505
rect 24857 53496 24869 53499
rect 23952 53468 24869 53496
rect 2409 53431 2467 53437
rect 2409 53397 2421 53431
rect 2455 53428 2467 53431
rect 2498 53428 2504 53440
rect 2455 53400 2504 53428
rect 2455 53397 2467 53400
rect 2409 53391 2467 53397
rect 2498 53388 2504 53400
rect 2556 53388 2562 53440
rect 5442 53388 5448 53440
rect 5500 53428 5506 53440
rect 23952 53437 23980 53468
rect 24857 53465 24869 53468
rect 24903 53465 24915 53499
rect 24857 53459 24915 53465
rect 31680 53437 31708 53536
rect 32306 53524 32312 53576
rect 32364 53564 32370 53576
rect 32401 53567 32459 53573
rect 32401 53564 32413 53567
rect 32364 53536 32413 53564
rect 32364 53524 32370 53536
rect 32401 53533 32413 53536
rect 32447 53533 32459 53567
rect 32582 53564 32588 53576
rect 32543 53536 32588 53564
rect 32401 53527 32459 53533
rect 32582 53524 32588 53536
rect 32640 53524 32646 53576
rect 32674 53524 32680 53576
rect 32732 53564 32738 53576
rect 33137 53567 33195 53573
rect 33137 53564 33149 53567
rect 32732 53536 33149 53564
rect 32732 53524 32738 53536
rect 33137 53533 33149 53536
rect 33183 53564 33195 53567
rect 33873 53567 33931 53573
rect 33873 53564 33885 53567
rect 33183 53536 33885 53564
rect 33183 53533 33195 53536
rect 33137 53527 33195 53533
rect 33873 53533 33885 53536
rect 33919 53564 33931 53567
rect 38654 53564 38660 53576
rect 33919 53536 38660 53564
rect 33919 53533 33931 53536
rect 33873 53527 33931 53533
rect 38654 53524 38660 53536
rect 38712 53564 38718 53576
rect 39393 53567 39451 53573
rect 39393 53564 39405 53567
rect 38712 53536 39405 53564
rect 38712 53524 38718 53536
rect 39393 53533 39405 53536
rect 39439 53533 39451 53567
rect 39393 53527 39451 53533
rect 57701 53567 57759 53573
rect 57701 53533 57713 53567
rect 57747 53564 57759 53567
rect 58342 53564 58348 53576
rect 57747 53536 58348 53564
rect 57747 53533 57759 53536
rect 57701 53527 57759 53533
rect 31849 53499 31907 53505
rect 31849 53465 31861 53499
rect 31895 53496 31907 53499
rect 35342 53496 35348 53508
rect 31895 53468 35348 53496
rect 31895 53465 31907 53468
rect 31849 53459 31907 53465
rect 35342 53456 35348 53468
rect 35400 53456 35406 53508
rect 37550 53456 37556 53508
rect 37608 53496 37614 53508
rect 38197 53499 38255 53505
rect 38197 53496 38209 53499
rect 37608 53468 38209 53496
rect 37608 53456 37614 53468
rect 38197 53465 38209 53468
rect 38243 53465 38255 53499
rect 39408 53496 39436 53527
rect 58342 53524 58348 53536
rect 58400 53524 58406 53576
rect 40405 53499 40463 53505
rect 40405 53496 40417 53499
rect 39408 53468 40417 53496
rect 38197 53459 38255 53465
rect 40405 53465 40417 53468
rect 40451 53465 40463 53499
rect 40405 53459 40463 53465
rect 23937 53431 23995 53437
rect 23937 53428 23949 53431
rect 5500 53400 23949 53428
rect 5500 53388 5506 53400
rect 23937 53397 23949 53400
rect 23983 53397 23995 53431
rect 23937 53391 23995 53397
rect 31665 53431 31723 53437
rect 31665 53397 31677 53431
rect 31711 53428 31723 53431
rect 32582 53428 32588 53440
rect 31711 53400 32588 53428
rect 31711 53397 31723 53400
rect 31665 53391 31723 53397
rect 32582 53388 32588 53400
rect 32640 53388 32646 53440
rect 58161 53431 58219 53437
rect 58161 53397 58173 53431
rect 58207 53428 58219 53431
rect 58526 53428 58532 53440
rect 58207 53400 58532 53428
rect 58207 53397 58219 53400
rect 58161 53391 58219 53397
rect 58526 53388 58532 53400
rect 58584 53388 58590 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 28994 53184 29000 53236
rect 29052 53224 29058 53236
rect 29549 53227 29607 53233
rect 29549 53224 29561 53227
rect 29052 53196 29561 53224
rect 29052 53184 29058 53196
rect 29549 53193 29561 53196
rect 29595 53193 29607 53227
rect 29549 53187 29607 53193
rect 32585 53227 32643 53233
rect 32585 53193 32597 53227
rect 32631 53224 32643 53227
rect 32766 53224 32772 53236
rect 32631 53196 32772 53224
rect 32631 53193 32643 53196
rect 32585 53187 32643 53193
rect 32766 53184 32772 53196
rect 32824 53184 32830 53236
rect 39574 53184 39580 53236
rect 39632 53224 39638 53236
rect 40221 53227 40279 53233
rect 40221 53224 40233 53227
rect 39632 53196 40233 53224
rect 39632 53184 39638 53196
rect 40221 53193 40233 53196
rect 40267 53193 40279 53227
rect 40221 53187 40279 53193
rect 32398 53156 32404 53168
rect 29380 53128 32404 53156
rect 2406 53048 2412 53100
rect 2464 53088 2470 53100
rect 10594 53088 10600 53100
rect 2464 53060 10600 53088
rect 2464 53048 2470 53060
rect 10594 53048 10600 53060
rect 10652 53048 10658 53100
rect 29380 53029 29408 53128
rect 32398 53116 32404 53128
rect 32456 53116 32462 53168
rect 29914 53088 29920 53100
rect 29875 53060 29920 53088
rect 29914 53048 29920 53060
rect 29972 53048 29978 53100
rect 32306 53048 32312 53100
rect 32364 53088 32370 53100
rect 32677 53091 32735 53097
rect 32677 53088 32689 53091
rect 32364 53060 32689 53088
rect 32364 53048 32370 53060
rect 32677 53057 32689 53060
rect 32723 53057 32735 53091
rect 32677 53051 32735 53057
rect 29365 53023 29423 53029
rect 29365 53020 29377 53023
rect 28828 52992 29377 53020
rect 28828 52896 28856 52992
rect 29365 52989 29377 52992
rect 29411 52989 29423 53023
rect 29365 52983 29423 52989
rect 29730 52980 29736 53032
rect 29788 53020 29794 53032
rect 29825 53023 29883 53029
rect 29825 53020 29837 53023
rect 29788 52992 29837 53020
rect 29788 52980 29794 52992
rect 29825 52989 29837 52992
rect 29871 52989 29883 53023
rect 29825 52983 29883 52989
rect 28810 52884 28816 52896
rect 28771 52856 28816 52884
rect 28810 52844 28816 52856
rect 28868 52844 28874 52896
rect 39666 52884 39672 52896
rect 39627 52856 39672 52884
rect 39666 52844 39672 52856
rect 39724 52844 39730 52896
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 29089 52683 29147 52689
rect 29089 52649 29101 52683
rect 29135 52680 29147 52683
rect 29730 52680 29736 52692
rect 29135 52652 29736 52680
rect 29135 52649 29147 52652
rect 29089 52643 29147 52649
rect 29730 52640 29736 52652
rect 29788 52640 29794 52692
rect 1670 52612 1676 52624
rect 1631 52584 1676 52612
rect 1670 52572 1676 52584
rect 1728 52572 1734 52624
rect 58161 52615 58219 52621
rect 58161 52581 58173 52615
rect 58207 52612 58219 52615
rect 58710 52612 58716 52624
rect 58207 52584 58716 52612
rect 58207 52581 58219 52584
rect 58161 52575 58219 52581
rect 58710 52572 58716 52584
rect 58768 52572 58774 52624
rect 1857 52479 1915 52485
rect 1857 52445 1869 52479
rect 1903 52476 1915 52479
rect 2409 52479 2467 52485
rect 2409 52476 2421 52479
rect 1903 52448 2421 52476
rect 1903 52445 1915 52448
rect 1857 52439 1915 52445
rect 2409 52445 2421 52448
rect 2455 52476 2467 52479
rect 2774 52476 2780 52488
rect 2455 52448 2780 52476
rect 2455 52445 2467 52448
rect 2409 52439 2467 52445
rect 2774 52436 2780 52448
rect 2832 52436 2838 52488
rect 55490 52436 55496 52488
rect 55548 52476 55554 52488
rect 56870 52476 56876 52488
rect 55548 52448 56876 52476
rect 55548 52436 55554 52448
rect 56870 52436 56876 52448
rect 56928 52436 56934 52488
rect 57701 52479 57759 52485
rect 57701 52445 57713 52479
rect 57747 52476 57759 52479
rect 58342 52476 58348 52488
rect 57747 52448 58348 52476
rect 57747 52445 57759 52448
rect 57701 52439 57759 52445
rect 58342 52436 58348 52448
rect 58400 52436 58406 52488
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1857 52003 1915 52009
rect 1857 51969 1869 52003
rect 1903 52000 1915 52003
rect 57517 52003 57575 52009
rect 1903 51972 2452 52000
rect 1903 51969 1915 51972
rect 1857 51963 1915 51969
rect 1670 51796 1676 51808
rect 1631 51768 1676 51796
rect 1670 51756 1676 51768
rect 1728 51756 1734 51808
rect 2424 51805 2452 51972
rect 57517 51969 57529 52003
rect 57563 52000 57575 52003
rect 58342 52000 58348 52012
rect 57563 51972 58348 52000
rect 57563 51969 57575 51972
rect 57517 51963 57575 51969
rect 58342 51960 58348 51972
rect 58400 51960 58406 52012
rect 2409 51799 2467 51805
rect 2409 51765 2421 51799
rect 2455 51796 2467 51799
rect 4798 51796 4804 51808
rect 2455 51768 4804 51796
rect 2455 51765 2467 51768
rect 2409 51759 2467 51765
rect 4798 51756 4804 51768
rect 4856 51756 4862 51808
rect 58161 51799 58219 51805
rect 58161 51765 58173 51799
rect 58207 51796 58219 51799
rect 59078 51796 59084 51808
rect 58207 51768 59084 51796
rect 58207 51765 58219 51768
rect 58161 51759 58219 51765
rect 59078 51756 59084 51768
rect 59136 51756 59142 51808
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 58342 51252 58348 51264
rect 58303 51224 58348 51252
rect 58342 51212 58348 51224
rect 58400 51212 58406 51264
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 2498 51008 2504 51060
rect 2556 51048 2562 51060
rect 3602 51048 3608 51060
rect 2556 51020 3608 51048
rect 2556 51008 2562 51020
rect 3602 51008 3608 51020
rect 3660 51008 3666 51060
rect 1857 50915 1915 50921
rect 1857 50881 1869 50915
rect 1903 50912 1915 50915
rect 58342 50912 58348 50924
rect 1903 50884 2452 50912
rect 58303 50884 58348 50912
rect 1903 50881 1915 50884
rect 1857 50875 1915 50881
rect 1670 50776 1676 50788
rect 1631 50748 1676 50776
rect 1670 50736 1676 50748
rect 1728 50736 1734 50788
rect 2424 50717 2452 50884
rect 58342 50872 58348 50884
rect 58400 50872 58406 50924
rect 2409 50711 2467 50717
rect 2409 50677 2421 50711
rect 2455 50708 2467 50711
rect 2590 50708 2596 50720
rect 2455 50680 2596 50708
rect 2455 50677 2467 50680
rect 2409 50671 2467 50677
rect 2590 50668 2596 50680
rect 2648 50668 2654 50720
rect 58161 50711 58219 50717
rect 58161 50677 58173 50711
rect 58207 50708 58219 50711
rect 58802 50708 58808 50720
rect 58207 50680 58808 50708
rect 58207 50677 58219 50680
rect 58161 50671 58219 50677
rect 58802 50668 58808 50680
rect 58860 50668 58866 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 2774 50328 2780 50380
rect 2832 50368 2838 50380
rect 19058 50368 19064 50380
rect 2832 50340 19064 50368
rect 2832 50328 2838 50340
rect 19058 50328 19064 50340
rect 19116 50328 19122 50380
rect 1857 50303 1915 50309
rect 1857 50269 1869 50303
rect 1903 50300 1915 50303
rect 1946 50300 1952 50312
rect 1903 50272 1952 50300
rect 1903 50269 1915 50272
rect 1857 50263 1915 50269
rect 1946 50260 1952 50272
rect 2004 50300 2010 50312
rect 2317 50303 2375 50309
rect 2317 50300 2329 50303
rect 2004 50272 2329 50300
rect 2004 50260 2010 50272
rect 2317 50269 2329 50272
rect 2363 50269 2375 50303
rect 2317 50263 2375 50269
rect 57701 50303 57759 50309
rect 57701 50269 57713 50303
rect 57747 50300 57759 50303
rect 58342 50300 58348 50312
rect 57747 50272 58348 50300
rect 57747 50269 57759 50272
rect 57701 50263 57759 50269
rect 58342 50260 58348 50272
rect 58400 50260 58406 50312
rect 1670 50164 1676 50176
rect 1631 50136 1676 50164
rect 1670 50124 1676 50136
rect 1728 50124 1734 50176
rect 58161 50167 58219 50173
rect 58161 50133 58173 50167
rect 58207 50164 58219 50167
rect 58434 50164 58440 50176
rect 58207 50136 58440 50164
rect 58207 50133 58219 50136
rect 58161 50127 58219 50133
rect 58434 50124 58440 50136
rect 58492 50124 58498 50176
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1857 49215 1915 49221
rect 1857 49181 1869 49215
rect 1903 49212 1915 49215
rect 2409 49215 2467 49221
rect 2409 49212 2421 49215
rect 1903 49184 2421 49212
rect 1903 49181 1915 49184
rect 1857 49175 1915 49181
rect 2409 49181 2421 49184
rect 2455 49212 2467 49215
rect 10778 49212 10784 49224
rect 2455 49184 10784 49212
rect 2455 49181 2467 49184
rect 2409 49175 2467 49181
rect 10778 49172 10784 49184
rect 10836 49172 10842 49224
rect 57701 49215 57759 49221
rect 57701 49181 57713 49215
rect 57747 49212 57759 49215
rect 58342 49212 58348 49224
rect 57747 49184 58348 49212
rect 57747 49181 57759 49184
rect 57701 49175 57759 49181
rect 58342 49172 58348 49184
rect 58400 49172 58406 49224
rect 1670 49076 1676 49088
rect 1631 49048 1676 49076
rect 1670 49036 1676 49048
rect 1728 49036 1734 49088
rect 57974 49036 57980 49088
rect 58032 49076 58038 49088
rect 58161 49079 58219 49085
rect 58161 49076 58173 49079
rect 58032 49048 58173 49076
rect 58032 49036 58038 49048
rect 58161 49045 58173 49048
rect 58207 49045 58219 49079
rect 58161 49039 58219 49045
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1857 48739 1915 48745
rect 1857 48705 1869 48739
rect 1903 48736 1915 48739
rect 2038 48736 2044 48748
rect 1903 48708 2044 48736
rect 1903 48705 1915 48708
rect 1857 48699 1915 48705
rect 2038 48696 2044 48708
rect 2096 48696 2102 48748
rect 57517 48739 57575 48745
rect 57517 48705 57529 48739
rect 57563 48736 57575 48739
rect 58342 48736 58348 48748
rect 57563 48708 58348 48736
rect 57563 48705 57575 48708
rect 57517 48699 57575 48705
rect 58342 48696 58348 48708
rect 58400 48696 58406 48748
rect 1670 48532 1676 48544
rect 1631 48504 1676 48532
rect 1670 48492 1676 48504
rect 1728 48492 1734 48544
rect 2038 48492 2044 48544
rect 2096 48532 2102 48544
rect 2317 48535 2375 48541
rect 2317 48532 2329 48535
rect 2096 48504 2329 48532
rect 2096 48492 2102 48504
rect 2317 48501 2329 48504
rect 2363 48501 2375 48535
rect 2317 48495 2375 48501
rect 57330 48492 57336 48544
rect 57388 48532 57394 48544
rect 58161 48535 58219 48541
rect 58161 48532 58173 48535
rect 57388 48504 58173 48532
rect 57388 48492 57394 48504
rect 58161 48501 58173 48504
rect 58207 48501 58219 48535
rect 58161 48495 58219 48501
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 58342 47988 58348 48000
rect 58303 47960 58348 47988
rect 58342 47948 58348 47960
rect 58400 47948 58406 48000
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1857 47651 1915 47657
rect 1857 47617 1869 47651
rect 1903 47648 1915 47651
rect 58342 47648 58348 47660
rect 1903 47620 2452 47648
rect 58303 47620 58348 47648
rect 1903 47617 1915 47620
rect 1857 47611 1915 47617
rect 1670 47512 1676 47524
rect 1631 47484 1676 47512
rect 1670 47472 1676 47484
rect 1728 47472 1734 47524
rect 2424 47453 2452 47620
rect 58342 47608 58348 47620
rect 58400 47608 58406 47660
rect 2866 47540 2872 47592
rect 2924 47580 2930 47592
rect 15194 47580 15200 47592
rect 2924 47552 15200 47580
rect 2924 47540 2930 47552
rect 15194 47540 15200 47552
rect 15252 47540 15258 47592
rect 2409 47447 2467 47453
rect 2409 47413 2421 47447
rect 2455 47444 2467 47447
rect 4706 47444 4712 47456
rect 2455 47416 4712 47444
rect 2455 47413 2467 47416
rect 2409 47407 2467 47413
rect 4706 47404 4712 47416
rect 4764 47404 4770 47456
rect 58161 47447 58219 47453
rect 58161 47413 58173 47447
rect 58207 47444 58219 47447
rect 58250 47444 58256 47456
rect 58207 47416 58256 47444
rect 58207 47413 58219 47416
rect 58161 47407 58219 47413
rect 58250 47404 58256 47416
rect 58308 47404 58314 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 58161 47175 58219 47181
rect 58161 47141 58173 47175
rect 58207 47172 58219 47175
rect 58618 47172 58624 47184
rect 58207 47144 58624 47172
rect 58207 47141 58219 47144
rect 58161 47135 58219 47141
rect 58618 47132 58624 47144
rect 58676 47132 58682 47184
rect 1857 47039 1915 47045
rect 1857 47005 1869 47039
rect 1903 47005 1915 47039
rect 1857 46999 1915 47005
rect 57701 47039 57759 47045
rect 57701 47005 57713 47039
rect 57747 47036 57759 47039
rect 58342 47036 58348 47048
rect 57747 47008 58348 47036
rect 57747 47005 57759 47008
rect 57701 46999 57759 47005
rect 1872 46968 1900 46999
rect 58342 46996 58348 47008
rect 58400 46996 58406 47048
rect 2130 46968 2136 46980
rect 1872 46940 2136 46968
rect 2130 46928 2136 46940
rect 2188 46968 2194 46980
rect 2317 46971 2375 46977
rect 2317 46968 2329 46971
rect 2188 46940 2329 46968
rect 2188 46928 2194 46940
rect 2317 46937 2329 46940
rect 2363 46937 2375 46971
rect 2317 46931 2375 46937
rect 1670 46900 1676 46912
rect 1631 46872 1676 46900
rect 1670 46860 1676 46872
rect 1728 46860 1734 46912
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 1857 45951 1915 45957
rect 1857 45917 1869 45951
rect 1903 45948 1915 45951
rect 57701 45951 57759 45957
rect 1903 45920 2452 45948
rect 1903 45917 1915 45920
rect 1857 45911 1915 45917
rect 1670 45812 1676 45824
rect 1631 45784 1676 45812
rect 1670 45772 1676 45784
rect 1728 45772 1734 45824
rect 2424 45821 2452 45920
rect 57701 45917 57713 45951
rect 57747 45948 57759 45951
rect 58342 45948 58348 45960
rect 57747 45920 58348 45948
rect 57747 45917 57759 45920
rect 57701 45911 57759 45917
rect 58342 45908 58348 45920
rect 58400 45908 58406 45960
rect 2409 45815 2467 45821
rect 2409 45781 2421 45815
rect 2455 45812 2467 45815
rect 3050 45812 3056 45824
rect 2455 45784 3056 45812
rect 2455 45781 2467 45784
rect 2409 45775 2467 45781
rect 3050 45772 3056 45784
rect 3108 45772 3114 45824
rect 58161 45815 58219 45821
rect 58161 45781 58173 45815
rect 58207 45812 58219 45815
rect 59630 45812 59636 45824
rect 58207 45784 59636 45812
rect 58207 45781 58219 45784
rect 58161 45775 58219 45781
rect 59630 45772 59636 45784
rect 59688 45772 59694 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1857 45475 1915 45481
rect 1857 45441 1869 45475
rect 1903 45472 1915 45475
rect 57517 45475 57575 45481
rect 1903 45444 2452 45472
rect 1903 45441 1915 45444
rect 1857 45435 1915 45441
rect 1670 45268 1676 45280
rect 1631 45240 1676 45268
rect 1670 45228 1676 45240
rect 1728 45228 1734 45280
rect 2424 45277 2452 45444
rect 57517 45441 57529 45475
rect 57563 45472 57575 45475
rect 58342 45472 58348 45484
rect 57563 45444 58348 45472
rect 57563 45441 57575 45444
rect 57517 45435 57575 45441
rect 58342 45432 58348 45444
rect 58400 45432 58406 45484
rect 2409 45271 2467 45277
rect 2409 45237 2421 45271
rect 2455 45268 2467 45271
rect 9582 45268 9588 45280
rect 2455 45240 9588 45268
rect 2455 45237 2467 45240
rect 2409 45231 2467 45237
rect 9582 45228 9588 45240
rect 9640 45228 9646 45280
rect 58161 45271 58219 45277
rect 58161 45237 58173 45271
rect 58207 45268 58219 45271
rect 59262 45268 59268 45280
rect 58207 45240 59268 45268
rect 58207 45237 58219 45240
rect 58161 45231 58219 45237
rect 59262 45228 59268 45240
rect 59320 45228 59326 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 2406 44820 2412 44872
rect 2464 44860 2470 44872
rect 17402 44860 17408 44872
rect 2464 44832 17408 44860
rect 2464 44820 2470 44832
rect 17402 44820 17408 44832
rect 17460 44820 17466 44872
rect 58342 44724 58348 44736
rect 58303 44696 58348 44724
rect 58342 44684 58348 44696
rect 58400 44684 58406 44736
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1857 44387 1915 44393
rect 1857 44353 1869 44387
rect 1903 44384 1915 44387
rect 58342 44384 58348 44396
rect 1903 44356 2452 44384
rect 58303 44356 58348 44384
rect 1903 44353 1915 44356
rect 1857 44347 1915 44353
rect 1670 44248 1676 44260
rect 1631 44220 1676 44248
rect 1670 44208 1676 44220
rect 1728 44208 1734 44260
rect 2424 44189 2452 44356
rect 58342 44344 58348 44356
rect 58400 44344 58406 44396
rect 2409 44183 2467 44189
rect 2409 44149 2421 44183
rect 2455 44180 2467 44183
rect 6178 44180 6184 44192
rect 2455 44152 6184 44180
rect 2455 44149 2467 44152
rect 2409 44143 2467 44149
rect 6178 44140 6184 44152
rect 6236 44140 6242 44192
rect 58161 44183 58219 44189
rect 58161 44149 58173 44183
rect 58207 44180 58219 44183
rect 59354 44180 59360 44192
rect 58207 44152 59360 44180
rect 58207 44149 58219 44152
rect 58161 44143 58219 44149
rect 59354 44140 59360 44152
rect 59412 44140 59418 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1857 43775 1915 43781
rect 1857 43741 1869 43775
rect 1903 43772 1915 43775
rect 57701 43775 57759 43781
rect 1903 43744 2452 43772
rect 1903 43741 1915 43744
rect 1857 43735 1915 43741
rect 1670 43636 1676 43648
rect 1631 43608 1676 43636
rect 1670 43596 1676 43608
rect 1728 43596 1734 43648
rect 2424 43645 2452 43744
rect 57701 43741 57713 43775
rect 57747 43772 57759 43775
rect 58342 43772 58348 43784
rect 57747 43744 58348 43772
rect 57747 43741 57759 43744
rect 57701 43735 57759 43741
rect 58342 43732 58348 43744
rect 58400 43732 58406 43784
rect 2409 43639 2467 43645
rect 2409 43605 2421 43639
rect 2455 43636 2467 43639
rect 3970 43636 3976 43648
rect 2455 43608 3976 43636
rect 2455 43605 2467 43608
rect 2409 43599 2467 43605
rect 3970 43596 3976 43608
rect 4028 43596 4034 43648
rect 56778 43596 56784 43648
rect 56836 43636 56842 43648
rect 58161 43639 58219 43645
rect 58161 43636 58173 43639
rect 56836 43608 58173 43636
rect 56836 43596 56842 43608
rect 58161 43605 58173 43608
rect 58207 43605 58219 43639
rect 58161 43599 58219 43605
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 1857 42687 1915 42693
rect 1857 42653 1869 42687
rect 1903 42684 1915 42687
rect 2409 42687 2467 42693
rect 2409 42684 2421 42687
rect 1903 42656 2421 42684
rect 1903 42653 1915 42656
rect 1857 42647 1915 42653
rect 2409 42653 2421 42656
rect 2455 42684 2467 42687
rect 15930 42684 15936 42696
rect 2455 42656 15936 42684
rect 2455 42653 2467 42656
rect 2409 42647 2467 42653
rect 15930 42644 15936 42656
rect 15988 42644 15994 42696
rect 57701 42687 57759 42693
rect 57701 42653 57713 42687
rect 57747 42684 57759 42687
rect 58342 42684 58348 42696
rect 57747 42656 58348 42684
rect 57747 42653 57759 42656
rect 57701 42647 57759 42653
rect 58342 42644 58348 42656
rect 58400 42644 58406 42696
rect 1670 42548 1676 42560
rect 1631 42520 1676 42548
rect 1670 42508 1676 42520
rect 1728 42508 1734 42560
rect 57790 42508 57796 42560
rect 57848 42548 57854 42560
rect 58161 42551 58219 42557
rect 58161 42548 58173 42551
rect 57848 42520 58173 42548
rect 57848 42508 57854 42520
rect 58161 42517 58173 42520
rect 58207 42517 58219 42551
rect 58161 42511 58219 42517
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 1857 42211 1915 42217
rect 1857 42177 1869 42211
rect 1903 42208 1915 42211
rect 2409 42211 2467 42217
rect 2409 42208 2421 42211
rect 1903 42180 2421 42208
rect 1903 42177 1915 42180
rect 1857 42171 1915 42177
rect 2409 42177 2421 42180
rect 2455 42208 2467 42211
rect 14458 42208 14464 42220
rect 2455 42180 14464 42208
rect 2455 42177 2467 42180
rect 2409 42171 2467 42177
rect 14458 42168 14464 42180
rect 14516 42168 14522 42220
rect 57517 42211 57575 42217
rect 57517 42177 57529 42211
rect 57563 42208 57575 42211
rect 58342 42208 58348 42220
rect 57563 42180 58348 42208
rect 57563 42177 57575 42180
rect 57517 42171 57575 42177
rect 58342 42168 58348 42180
rect 58400 42168 58406 42220
rect 1670 42004 1676 42016
rect 1631 41976 1676 42004
rect 1670 41964 1676 41976
rect 1728 41964 1734 42016
rect 58161 42007 58219 42013
rect 58161 41973 58173 42007
rect 58207 42004 58219 42007
rect 58986 42004 58992 42016
rect 58207 41976 58992 42004
rect 58207 41973 58219 41976
rect 58161 41967 58219 41973
rect 58986 41964 58992 41976
rect 59044 41964 59050 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 58342 41460 58348 41472
rect 58303 41432 58348 41460
rect 58342 41420 58348 41432
rect 58400 41420 58406 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1857 41123 1915 41129
rect 1857 41089 1869 41123
rect 1903 41120 1915 41123
rect 58342 41120 58348 41132
rect 1903 41092 2452 41120
rect 58303 41092 58348 41120
rect 1903 41089 1915 41092
rect 1857 41083 1915 41089
rect 1670 40984 1676 40996
rect 1631 40956 1676 40984
rect 1670 40944 1676 40956
rect 1728 40944 1734 40996
rect 2424 40925 2452 41092
rect 58342 41080 58348 41092
rect 58400 41080 58406 41132
rect 2409 40919 2467 40925
rect 2409 40885 2421 40919
rect 2455 40916 2467 40919
rect 7558 40916 7564 40928
rect 2455 40888 7564 40916
rect 2455 40885 2467 40888
rect 2409 40879 2467 40885
rect 7558 40876 7564 40888
rect 7616 40876 7622 40928
rect 57606 40876 57612 40928
rect 57664 40916 57670 40928
rect 58161 40919 58219 40925
rect 58161 40916 58173 40919
rect 57664 40888 58173 40916
rect 57664 40876 57670 40888
rect 58161 40885 58173 40888
rect 58207 40885 58219 40919
rect 58161 40879 58219 40885
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 1857 40511 1915 40517
rect 1857 40477 1869 40511
rect 1903 40508 1915 40511
rect 57701 40511 57759 40517
rect 1903 40480 2452 40508
rect 1903 40477 1915 40480
rect 1857 40471 1915 40477
rect 1670 40372 1676 40384
rect 1631 40344 1676 40372
rect 1670 40332 1676 40344
rect 1728 40332 1734 40384
rect 2424 40381 2452 40480
rect 57701 40477 57713 40511
rect 57747 40508 57759 40511
rect 58342 40508 58348 40520
rect 57747 40480 58348 40508
rect 57747 40477 57759 40480
rect 57701 40471 57759 40477
rect 58342 40468 58348 40480
rect 58400 40468 58406 40520
rect 2409 40375 2467 40381
rect 2409 40341 2421 40375
rect 2455 40372 2467 40375
rect 6270 40372 6276 40384
rect 2455 40344 6276 40372
rect 2455 40341 2467 40344
rect 2409 40335 2467 40341
rect 6270 40332 6276 40344
rect 6328 40332 6334 40384
rect 57054 40332 57060 40384
rect 57112 40372 57118 40384
rect 58161 40375 58219 40381
rect 58161 40372 58173 40375
rect 57112 40344 58173 40372
rect 57112 40332 57118 40344
rect 58161 40341 58173 40344
rect 58207 40341 58219 40375
rect 58161 40335 58219 40341
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 57238 40128 57244 40180
rect 57296 40168 57302 40180
rect 58161 40171 58219 40177
rect 58161 40168 58173 40171
rect 57296 40140 58173 40168
rect 57296 40128 57302 40140
rect 58161 40137 58173 40140
rect 58207 40137 58219 40171
rect 58161 40131 58219 40137
rect 57882 40100 57888 40112
rect 57532 40072 57888 40100
rect 57532 40041 57560 40072
rect 57882 40060 57888 40072
rect 57940 40100 57946 40112
rect 57940 40072 58388 40100
rect 57940 40060 57946 40072
rect 58360 40041 58388 40072
rect 57517 40035 57575 40041
rect 57517 40001 57529 40035
rect 57563 40001 57575 40035
rect 57517 39995 57575 40001
rect 58345 40035 58403 40041
rect 58345 40001 58357 40035
rect 58391 40001 58403 40035
rect 58345 39995 58403 40001
rect 56410 39828 56416 39840
rect 56371 39800 56416 39828
rect 56410 39788 56416 39800
rect 56468 39788 56474 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 56042 39448 56048 39500
rect 56100 39488 56106 39500
rect 56410 39488 56416 39500
rect 56100 39460 56416 39488
rect 56100 39448 56106 39460
rect 56410 39448 56416 39460
rect 56468 39488 56474 39500
rect 56468 39460 56994 39488
rect 56468 39448 56474 39460
rect 1857 39423 1915 39429
rect 1857 39389 1869 39423
rect 1903 39420 1915 39423
rect 57238 39420 57244 39432
rect 1903 39392 2452 39420
rect 57199 39392 57244 39420
rect 1903 39389 1915 39392
rect 1857 39383 1915 39389
rect 1670 39284 1676 39296
rect 1631 39256 1676 39284
rect 1670 39244 1676 39256
rect 1728 39244 1734 39296
rect 2424 39293 2452 39392
rect 57238 39380 57244 39392
rect 57296 39380 57302 39432
rect 57698 39420 57704 39432
rect 57659 39392 57704 39420
rect 57698 39380 57704 39392
rect 57756 39380 57762 39432
rect 57609 39355 57667 39361
rect 57609 39352 57621 39355
rect 56152 39324 57621 39352
rect 56152 39296 56180 39324
rect 57609 39321 57621 39324
rect 57655 39321 57667 39355
rect 57974 39352 57980 39364
rect 57935 39324 57980 39352
rect 57609 39315 57667 39321
rect 57974 39312 57980 39324
rect 58032 39312 58038 39364
rect 2409 39287 2467 39293
rect 2409 39253 2421 39287
rect 2455 39284 2467 39287
rect 7650 39284 7656 39296
rect 2455 39256 7656 39284
rect 2455 39253 2467 39256
rect 2409 39247 2467 39253
rect 7650 39244 7656 39256
rect 7708 39244 7714 39296
rect 56134 39284 56140 39296
rect 56095 39256 56140 39284
rect 56134 39244 56140 39256
rect 56192 39244 56198 39296
rect 56594 39244 56600 39296
rect 56652 39284 56658 39296
rect 56689 39287 56747 39293
rect 56689 39284 56701 39287
rect 56652 39256 56701 39284
rect 56652 39244 56658 39256
rect 56689 39253 56701 39256
rect 56735 39253 56747 39287
rect 56870 39284 56876 39296
rect 56831 39256 56876 39284
rect 56689 39247 56747 39253
rect 56870 39244 56876 39256
rect 56928 39244 56934 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 56137 39083 56195 39089
rect 56137 39049 56149 39083
rect 56183 39080 56195 39083
rect 57146 39080 57152 39092
rect 56183 39052 57152 39080
rect 56183 39049 56195 39052
rect 56137 39043 56195 39049
rect 57146 39040 57152 39052
rect 57204 39040 57210 39092
rect 57241 39083 57299 39089
rect 57241 39049 57253 39083
rect 57287 39080 57299 39083
rect 57330 39080 57336 39092
rect 57287 39052 57336 39080
rect 57287 39049 57299 39052
rect 57241 39043 57299 39049
rect 57330 39040 57336 39052
rect 57388 39040 57394 39092
rect 58161 39083 58219 39089
rect 58161 39049 58173 39083
rect 58207 39049 58219 39083
rect 58161 39043 58219 39049
rect 56505 39015 56563 39021
rect 56505 38981 56517 39015
rect 56551 39012 56563 39015
rect 58176 39012 58204 39043
rect 56551 38984 58204 39012
rect 56551 38981 56563 38984
rect 56505 38975 56563 38981
rect 1857 38947 1915 38953
rect 1857 38913 1869 38947
rect 1903 38944 1915 38947
rect 1903 38916 2452 38944
rect 1903 38913 1915 38916
rect 1857 38907 1915 38913
rect 1670 38740 1676 38752
rect 1631 38712 1676 38740
rect 1670 38700 1676 38712
rect 1728 38700 1734 38752
rect 2424 38749 2452 38916
rect 55398 38904 55404 38956
rect 55456 38944 55462 38956
rect 56134 38944 56140 38956
rect 55456 38916 56140 38944
rect 55456 38904 55462 38916
rect 56134 38904 56140 38916
rect 56192 38944 56198 38956
rect 56873 38947 56931 38953
rect 56873 38944 56885 38947
rect 56192 38916 56885 38944
rect 56192 38904 56198 38916
rect 56873 38913 56885 38916
rect 56919 38913 56931 38947
rect 56873 38907 56931 38913
rect 56965 38947 57023 38953
rect 56965 38913 56977 38947
rect 57011 38944 57023 38947
rect 58158 38944 58164 38956
rect 57011 38916 58164 38944
rect 57011 38913 57023 38916
rect 56965 38907 57023 38913
rect 58158 38904 58164 38916
rect 58216 38904 58222 38956
rect 58342 38944 58348 38956
rect 58303 38916 58348 38944
rect 58342 38904 58348 38916
rect 58400 38904 58406 38956
rect 56042 38836 56048 38888
rect 56100 38876 56106 38888
rect 56100 38848 56258 38876
rect 56100 38836 56106 38848
rect 2409 38743 2467 38749
rect 2409 38709 2421 38743
rect 2455 38740 2467 38743
rect 2774 38740 2780 38752
rect 2455 38712 2780 38740
rect 2455 38709 2467 38712
rect 2409 38703 2467 38709
rect 2774 38700 2780 38712
rect 2832 38700 2838 38752
rect 55398 38740 55404 38752
rect 55359 38712 55404 38740
rect 55398 38700 55404 38712
rect 55456 38700 55462 38752
rect 55950 38740 55956 38752
rect 55911 38712 55956 38740
rect 55950 38700 55956 38712
rect 56008 38700 56014 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 57054 38536 57060 38548
rect 57015 38508 57060 38536
rect 57054 38496 57060 38508
rect 57112 38496 57118 38548
rect 57609 38539 57667 38545
rect 57609 38505 57621 38539
rect 57655 38536 57667 38539
rect 58158 38536 58164 38548
rect 57655 38508 58164 38536
rect 57655 38505 57667 38508
rect 57609 38499 57667 38505
rect 58158 38496 58164 38508
rect 58216 38496 58222 38548
rect 55769 38199 55827 38205
rect 55769 38165 55781 38199
rect 55815 38196 55827 38199
rect 56042 38196 56048 38208
rect 55815 38168 56048 38196
rect 55815 38165 55827 38168
rect 55769 38159 55827 38165
rect 56042 38156 56048 38168
rect 56100 38156 56106 38208
rect 58342 38196 58348 38208
rect 58303 38168 58348 38196
rect 58342 38156 58348 38168
rect 58400 38156 58406 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 58161 37995 58219 38001
rect 58161 37992 58173 37995
rect 55186 37964 58173 37992
rect 54665 37927 54723 37933
rect 54665 37893 54677 37927
rect 54711 37924 54723 37927
rect 54846 37924 54852 37936
rect 54711 37896 54852 37924
rect 54711 37893 54723 37896
rect 54665 37887 54723 37893
rect 54846 37884 54852 37896
rect 54904 37884 54910 37936
rect 55033 37927 55091 37933
rect 55033 37893 55045 37927
rect 55079 37924 55091 37927
rect 55186 37924 55214 37964
rect 58161 37961 58173 37964
rect 58207 37961 58219 37995
rect 58161 37955 58219 37961
rect 55490 37924 55496 37936
rect 55079 37896 55214 37924
rect 55451 37896 55496 37924
rect 55079 37893 55091 37896
rect 55033 37887 55091 37893
rect 55490 37884 55496 37896
rect 55548 37884 55554 37936
rect 55769 37927 55827 37933
rect 55769 37893 55781 37927
rect 55815 37893 55827 37927
rect 55769 37887 55827 37893
rect 1857 37859 1915 37865
rect 1857 37825 1869 37859
rect 1903 37856 1915 37859
rect 53929 37859 53987 37865
rect 1903 37828 2452 37856
rect 1903 37825 1915 37828
rect 1857 37819 1915 37825
rect 1670 37720 1676 37732
rect 1631 37692 1676 37720
rect 1670 37680 1676 37692
rect 1728 37680 1734 37732
rect 2424 37664 2452 37828
rect 53929 37825 53941 37859
rect 53975 37856 53987 37859
rect 55398 37856 55404 37868
rect 53975 37828 55404 37856
rect 53975 37825 53987 37828
rect 53929 37819 53987 37825
rect 55398 37816 55404 37828
rect 55456 37816 55462 37868
rect 55784 37856 55812 37887
rect 55858 37884 55864 37936
rect 55916 37924 55922 37936
rect 56413 37927 56471 37933
rect 56413 37924 56425 37927
rect 55916 37896 56425 37924
rect 55916 37884 55922 37896
rect 56413 37893 56425 37896
rect 56459 37893 56471 37927
rect 58250 37924 58256 37936
rect 56413 37887 56471 37893
rect 56520 37896 58256 37924
rect 56520 37856 56548 37896
rect 58250 37884 58256 37896
rect 58308 37884 58314 37936
rect 58342 37856 58348 37868
rect 55784 37828 56548 37856
rect 58303 37828 58348 37856
rect 58342 37816 58348 37828
rect 58400 37816 58406 37868
rect 2774 37748 2780 37800
rect 2832 37788 2838 37800
rect 4614 37788 4620 37800
rect 2832 37760 4620 37788
rect 2832 37748 2838 37760
rect 4614 37748 4620 37760
rect 4672 37748 4678 37800
rect 56042 37788 56048 37800
rect 55955 37760 56048 37788
rect 56042 37748 56048 37760
rect 56100 37788 56106 37800
rect 56502 37788 56508 37800
rect 56100 37760 56508 37788
rect 56100 37748 56106 37760
rect 56502 37748 56508 37760
rect 56560 37748 56566 37800
rect 2406 37652 2412 37664
rect 2367 37624 2412 37652
rect 2406 37612 2412 37624
rect 2464 37612 2470 37664
rect 54481 37655 54539 37661
rect 54481 37621 54493 37655
rect 54527 37652 54539 37655
rect 54570 37652 54576 37664
rect 54527 37624 54576 37652
rect 54527 37621 54539 37624
rect 54481 37615 54539 37621
rect 54570 37612 54576 37624
rect 54628 37612 54634 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 2406 37408 2412 37460
rect 2464 37448 2470 37460
rect 13630 37448 13636 37460
rect 2464 37420 13636 37448
rect 2464 37408 2470 37420
rect 13630 37408 13636 37420
rect 13688 37408 13694 37460
rect 54297 37451 54355 37457
rect 54297 37417 54309 37451
rect 54343 37448 54355 37451
rect 56042 37448 56048 37460
rect 54343 37420 56048 37448
rect 54343 37417 54355 37420
rect 54297 37411 54355 37417
rect 56042 37408 56048 37420
rect 56100 37408 56106 37460
rect 57149 37315 57207 37321
rect 57149 37281 57161 37315
rect 57195 37281 57207 37315
rect 57149 37275 57207 37281
rect 57701 37315 57759 37321
rect 57701 37281 57713 37315
rect 57747 37312 57759 37315
rect 57882 37312 57888 37324
rect 57747 37284 57888 37312
rect 57747 37281 57759 37284
rect 57701 37275 57759 37281
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37244 1915 37247
rect 57164 37244 57192 37275
rect 57882 37272 57888 37284
rect 57940 37272 57946 37324
rect 58342 37244 58348 37256
rect 1903 37216 2452 37244
rect 57164 37216 58348 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 2424 37120 2452 37216
rect 58342 37204 58348 37216
rect 58400 37204 58406 37256
rect 1670 37108 1676 37120
rect 1631 37080 1676 37108
rect 1670 37068 1676 37080
rect 1728 37068 1734 37120
rect 2406 37108 2412 37120
rect 2367 37080 2412 37108
rect 2406 37068 2412 37080
rect 2464 37068 2470 37120
rect 57422 37068 57428 37120
rect 57480 37108 57486 37120
rect 58161 37111 58219 37117
rect 58161 37108 58173 37111
rect 57480 37080 58173 37108
rect 57480 37068 57486 37080
rect 58161 37077 58173 37080
rect 58207 37077 58219 37111
rect 58161 37071 58219 37077
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 2406 36864 2412 36916
rect 2464 36904 2470 36916
rect 16574 36904 16580 36916
rect 2464 36876 16580 36904
rect 2464 36864 2470 36876
rect 16574 36864 16580 36876
rect 16632 36864 16638 36916
rect 57517 36907 57575 36913
rect 57517 36873 57529 36907
rect 57563 36904 57575 36907
rect 57974 36904 57980 36916
rect 57563 36876 57980 36904
rect 57563 36873 57575 36876
rect 57517 36867 57575 36873
rect 57974 36864 57980 36876
rect 58032 36904 58038 36916
rect 59170 36904 59176 36916
rect 58032 36876 59176 36904
rect 58032 36864 58038 36876
rect 59170 36864 59176 36876
rect 59228 36864 59234 36916
rect 57882 36728 57888 36780
rect 57940 36768 57946 36780
rect 58345 36771 58403 36777
rect 58345 36768 58357 36771
rect 57940 36740 58357 36768
rect 57940 36728 57946 36740
rect 58345 36737 58357 36740
rect 58391 36737 58403 36771
rect 58345 36731 58403 36737
rect 56502 36524 56508 36576
rect 56560 36564 56566 36576
rect 56597 36567 56655 36573
rect 56597 36564 56609 36567
rect 56560 36536 56609 36564
rect 56560 36524 56566 36536
rect 56597 36533 56609 36536
rect 56643 36533 56655 36567
rect 56597 36527 56655 36533
rect 58066 36524 58072 36576
rect 58124 36564 58130 36576
rect 58161 36567 58219 36573
rect 58161 36564 58173 36567
rect 58124 36536 58173 36564
rect 58124 36524 58130 36536
rect 58161 36533 58173 36536
rect 58207 36533 58219 36567
rect 58161 36527 58219 36533
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 53098 36252 53104 36304
rect 53156 36292 53162 36304
rect 56873 36295 56931 36301
rect 56873 36292 56885 36295
rect 53156 36264 56885 36292
rect 53156 36252 53162 36264
rect 56873 36261 56885 36264
rect 56919 36261 56931 36295
rect 56873 36255 56931 36261
rect 56502 36184 56508 36236
rect 56560 36224 56566 36236
rect 56560 36196 57178 36224
rect 56560 36184 56566 36196
rect 1857 36159 1915 36165
rect 1857 36125 1869 36159
rect 1903 36156 1915 36159
rect 2409 36159 2467 36165
rect 2409 36156 2421 36159
rect 1903 36128 2421 36156
rect 1903 36125 1915 36128
rect 1857 36119 1915 36125
rect 2409 36125 2421 36128
rect 2455 36156 2467 36159
rect 8478 36156 8484 36168
rect 2455 36128 8484 36156
rect 2455 36125 2467 36128
rect 2409 36119 2467 36125
rect 8478 36116 8484 36128
rect 8536 36116 8542 36168
rect 57422 36156 57428 36168
rect 57383 36128 57428 36156
rect 57422 36116 57428 36128
rect 57480 36116 57486 36168
rect 57885 36159 57943 36165
rect 57885 36125 57897 36159
rect 57931 36156 57943 36159
rect 57974 36156 57980 36168
rect 57931 36128 57980 36156
rect 57931 36125 57943 36128
rect 57885 36119 57943 36125
rect 57974 36116 57980 36128
rect 58032 36116 58038 36168
rect 55398 36048 55404 36100
rect 55456 36088 55462 36100
rect 56318 36088 56324 36100
rect 55456 36060 56324 36088
rect 55456 36048 55462 36060
rect 56318 36048 56324 36060
rect 56376 36088 56382 36100
rect 57793 36091 57851 36097
rect 57793 36088 57805 36091
rect 56376 36060 57805 36088
rect 56376 36048 56382 36060
rect 57793 36057 57805 36060
rect 57839 36057 57851 36091
rect 59446 36088 59452 36100
rect 57793 36051 57851 36057
rect 58084 36060 59452 36088
rect 1670 36020 1676 36032
rect 1631 35992 1676 36020
rect 1670 35980 1676 35992
rect 1728 35980 1734 36032
rect 57057 36023 57115 36029
rect 57057 35989 57069 36023
rect 57103 36020 57115 36023
rect 58084 36020 58112 36060
rect 59446 36048 59452 36060
rect 59504 36048 59510 36100
rect 57103 35992 58112 36020
rect 58161 36023 58219 36029
rect 57103 35989 57115 35992
rect 57057 35983 57115 35989
rect 58161 35989 58173 36023
rect 58207 36020 58219 36023
rect 58618 36020 58624 36032
rect 58207 35992 58624 36020
rect 58207 35989 58219 35992
rect 58161 35983 58219 35989
rect 58618 35980 58624 35992
rect 58676 35980 58682 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 57517 35819 57575 35825
rect 57517 35785 57529 35819
rect 57563 35816 57575 35819
rect 57974 35816 57980 35828
rect 57563 35788 57980 35816
rect 57563 35785 57575 35788
rect 57517 35779 57575 35785
rect 57974 35776 57980 35788
rect 58032 35816 58038 35828
rect 59538 35816 59544 35828
rect 58032 35788 59544 35816
rect 58032 35776 58038 35788
rect 59538 35776 59544 35788
rect 59596 35776 59602 35828
rect 1857 35683 1915 35689
rect 1857 35649 1869 35683
rect 1903 35680 1915 35683
rect 2409 35683 2467 35689
rect 2409 35680 2421 35683
rect 1903 35652 2421 35680
rect 1903 35649 1915 35652
rect 1857 35643 1915 35649
rect 2409 35649 2421 35652
rect 2455 35680 2467 35683
rect 11698 35680 11704 35692
rect 2455 35652 11704 35680
rect 2455 35649 2467 35652
rect 2409 35643 2467 35649
rect 11698 35640 11704 35652
rect 11756 35640 11762 35692
rect 56965 35683 57023 35689
rect 56965 35649 56977 35683
rect 57011 35680 57023 35683
rect 58342 35680 58348 35692
rect 57011 35652 58348 35680
rect 57011 35649 57023 35652
rect 56965 35643 57023 35649
rect 58342 35640 58348 35652
rect 58400 35640 58406 35692
rect 1670 35476 1676 35488
rect 1631 35448 1676 35476
rect 1670 35436 1676 35448
rect 1728 35436 1734 35488
rect 56229 35479 56287 35485
rect 56229 35445 56241 35479
rect 56275 35476 56287 35479
rect 56410 35476 56416 35488
rect 56275 35448 56416 35476
rect 56275 35445 56287 35448
rect 56229 35439 56287 35445
rect 56410 35436 56416 35448
rect 56468 35476 56474 35488
rect 57514 35476 57520 35488
rect 56468 35448 57520 35476
rect 56468 35436 56474 35448
rect 57514 35436 57520 35448
rect 57572 35436 57578 35488
rect 58158 35476 58164 35488
rect 58119 35448 58164 35476
rect 58158 35436 58164 35448
rect 58216 35436 58222 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 57146 35232 57152 35284
rect 57204 35272 57210 35284
rect 59630 35272 59636 35284
rect 57204 35244 59636 35272
rect 57204 35232 57210 35244
rect 59630 35232 59636 35244
rect 59688 35232 59694 35284
rect 6270 35164 6276 35216
rect 6328 35204 6334 35216
rect 16022 35204 16028 35216
rect 6328 35176 16028 35204
rect 6328 35164 6334 35176
rect 16022 35164 16028 35176
rect 16080 35164 16086 35216
rect 57974 35204 57980 35216
rect 57440 35176 57980 35204
rect 55766 35096 55772 35148
rect 55824 35136 55830 35148
rect 56318 35136 56324 35148
rect 55824 35108 56324 35136
rect 55824 35096 55830 35108
rect 56318 35096 56324 35108
rect 56376 35136 56382 35148
rect 57146 35145 57152 35148
rect 56965 35139 57023 35145
rect 56965 35136 56977 35139
rect 56376 35108 56977 35136
rect 56376 35096 56382 35108
rect 56965 35105 56977 35108
rect 57011 35105 57023 35139
rect 56965 35099 57023 35105
rect 57124 35139 57152 35145
rect 57124 35105 57136 35139
rect 57124 35099 57152 35105
rect 57146 35096 57152 35099
rect 57204 35096 57210 35148
rect 57241 35139 57299 35145
rect 57241 35105 57253 35139
rect 57287 35136 57299 35139
rect 57440 35136 57468 35176
rect 57974 35164 57980 35176
rect 58032 35164 58038 35216
rect 57287 35108 57468 35136
rect 57287 35105 57299 35108
rect 57241 35099 57299 35105
rect 57514 35096 57520 35148
rect 57572 35136 57578 35148
rect 57572 35108 57617 35136
rect 57572 35096 57578 35108
rect 58066 35096 58072 35148
rect 58124 35136 58130 35148
rect 58161 35139 58219 35145
rect 58161 35136 58173 35139
rect 58124 35108 58173 35136
rect 58124 35096 58130 35108
rect 58161 35105 58173 35108
rect 58207 35105 58219 35139
rect 58161 35099 58219 35105
rect 57977 35071 58035 35077
rect 57977 35037 57989 35071
rect 58023 35037 58035 35071
rect 57977 35031 58035 35037
rect 52362 34960 52368 35012
rect 52420 35000 52426 35012
rect 56321 35003 56379 35009
rect 56321 35000 56333 35003
rect 52420 34972 56333 35000
rect 52420 34960 52426 34972
rect 56321 34969 56333 34972
rect 56367 34969 56379 35003
rect 57992 35000 58020 35031
rect 58066 35000 58072 35012
rect 57992 34972 58072 35000
rect 56321 34963 56379 34969
rect 58066 34960 58072 34972
rect 58124 34960 58130 35012
rect 55030 34892 55036 34944
rect 55088 34932 55094 34944
rect 55766 34932 55772 34944
rect 55088 34904 55772 34932
rect 55088 34892 55094 34904
rect 55766 34892 55772 34904
rect 55824 34892 55830 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 55306 34688 55312 34740
rect 55364 34728 55370 34740
rect 56686 34728 56692 34740
rect 55364 34700 56692 34728
rect 55364 34688 55370 34700
rect 56686 34688 56692 34700
rect 56744 34688 56750 34740
rect 58158 34660 58164 34672
rect 56244 34632 58164 34660
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34561 1915 34595
rect 52362 34592 52368 34604
rect 52323 34564 52368 34592
rect 1857 34555 1915 34561
rect 1872 34524 1900 34555
rect 52362 34552 52368 34564
rect 52420 34552 52426 34604
rect 55306 34592 55312 34604
rect 55267 34564 55312 34592
rect 55306 34552 55312 34564
rect 55364 34552 55370 34604
rect 56244 34601 56272 34632
rect 58158 34620 58164 34632
rect 58216 34620 58222 34672
rect 56229 34595 56287 34601
rect 56229 34561 56241 34595
rect 56275 34561 56287 34595
rect 56229 34555 56287 34561
rect 57517 34595 57575 34601
rect 57517 34561 57529 34595
rect 57563 34592 57575 34595
rect 58342 34592 58348 34604
rect 57563 34564 58348 34592
rect 57563 34561 57575 34564
rect 57517 34555 57575 34561
rect 58342 34552 58348 34564
rect 58400 34552 58406 34604
rect 2409 34527 2467 34533
rect 2409 34524 2421 34527
rect 1872 34496 2421 34524
rect 2409 34493 2421 34496
rect 2455 34524 2467 34527
rect 6914 34524 6920 34536
rect 2455 34496 6920 34524
rect 2455 34493 2467 34496
rect 2409 34487 2467 34493
rect 6914 34484 6920 34496
rect 6972 34484 6978 34536
rect 51442 34484 51448 34536
rect 51500 34524 51506 34536
rect 52089 34527 52147 34533
rect 52089 34524 52101 34527
rect 51500 34496 52101 34524
rect 51500 34484 51506 34496
rect 52089 34493 52101 34496
rect 52135 34493 52147 34527
rect 52089 34487 52147 34493
rect 53929 34527 53987 34533
rect 53929 34493 53941 34527
rect 53975 34524 53987 34527
rect 55030 34524 55036 34536
rect 53975 34496 55036 34524
rect 53975 34493 53987 34496
rect 53929 34487 53987 34493
rect 55030 34484 55036 34496
rect 55088 34484 55094 34536
rect 55192 34527 55250 34533
rect 55192 34493 55204 34527
rect 55238 34524 55250 34527
rect 55238 34496 55812 34524
rect 55238 34493 55250 34496
rect 55192 34487 55250 34493
rect 1670 34456 1676 34468
rect 1631 34428 1676 34456
rect 1670 34416 1676 34428
rect 1728 34416 1734 34468
rect 55582 34416 55588 34468
rect 55640 34456 55646 34468
rect 55784 34456 55812 34496
rect 55858 34484 55864 34536
rect 55916 34524 55922 34536
rect 56045 34527 56103 34533
rect 56045 34524 56057 34527
rect 55916 34496 56057 34524
rect 55916 34484 55922 34496
rect 56045 34493 56057 34496
rect 56091 34493 56103 34527
rect 59262 34524 59268 34536
rect 56045 34487 56103 34493
rect 56152 34496 59268 34524
rect 56152 34456 56180 34496
rect 59262 34484 59268 34496
rect 59320 34484 59326 34536
rect 55640 34428 55733 34456
rect 55784 34428 56180 34456
rect 55640 34416 55646 34428
rect 54386 34388 54392 34400
rect 54347 34360 54392 34388
rect 54386 34348 54392 34360
rect 54444 34348 54450 34400
rect 55692 34388 55720 34428
rect 56410 34388 56416 34400
rect 55692 34360 56416 34388
rect 56410 34348 56416 34360
rect 56468 34348 56474 34400
rect 58158 34388 58164 34400
rect 58119 34360 58164 34388
rect 58158 34348 58164 34360
rect 58216 34348 58222 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 54297 34187 54355 34193
rect 54297 34153 54309 34187
rect 54343 34184 54355 34187
rect 55582 34184 55588 34196
rect 54343 34156 55588 34184
rect 54343 34153 54355 34156
rect 54297 34147 54355 34153
rect 55582 34144 55588 34156
rect 55640 34144 55646 34196
rect 56962 34076 56968 34128
rect 57020 34116 57026 34128
rect 58161 34119 58219 34125
rect 58161 34116 58173 34119
rect 57020 34088 58173 34116
rect 57020 34076 57026 34088
rect 58161 34085 58173 34088
rect 58207 34085 58219 34119
rect 58161 34079 58219 34085
rect 1857 33983 1915 33989
rect 1857 33949 1869 33983
rect 1903 33980 1915 33983
rect 2317 33983 2375 33989
rect 2317 33980 2329 33983
rect 1903 33952 2329 33980
rect 1903 33949 1915 33952
rect 1857 33943 1915 33949
rect 2317 33949 2329 33952
rect 2363 33980 2375 33983
rect 2498 33980 2504 33992
rect 2363 33952 2504 33980
rect 2363 33949 2375 33952
rect 2317 33943 2375 33949
rect 2498 33940 2504 33952
rect 2556 33940 2562 33992
rect 57149 33983 57207 33989
rect 57149 33949 57161 33983
rect 57195 33980 57207 33983
rect 58342 33980 58348 33992
rect 57195 33952 58348 33980
rect 57195 33949 57207 33952
rect 57149 33943 57207 33949
rect 58342 33940 58348 33952
rect 58400 33940 58406 33992
rect 1670 33844 1676 33856
rect 1631 33816 1676 33844
rect 1670 33804 1676 33816
rect 1728 33804 1734 33856
rect 57701 33847 57759 33853
rect 57701 33813 57713 33847
rect 57747 33844 57759 33847
rect 57790 33844 57796 33856
rect 57747 33816 57796 33844
rect 57747 33813 57759 33816
rect 57701 33807 57759 33813
rect 57790 33804 57796 33816
rect 57848 33804 57854 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 57517 33643 57575 33649
rect 57517 33609 57529 33643
rect 57563 33640 57575 33643
rect 57974 33640 57980 33652
rect 57563 33612 57980 33640
rect 57563 33609 57575 33612
rect 57517 33603 57575 33609
rect 57974 33600 57980 33612
rect 58032 33640 58038 33652
rect 58526 33640 58532 33652
rect 58032 33612 58532 33640
rect 58032 33600 58038 33612
rect 58526 33600 58532 33612
rect 58584 33600 58590 33652
rect 54386 33464 54392 33516
rect 54444 33504 54450 33516
rect 55033 33507 55091 33513
rect 55033 33504 55045 33507
rect 54444 33476 55045 33504
rect 54444 33464 54450 33476
rect 55033 33473 55045 33476
rect 55079 33473 55091 33507
rect 55033 33467 55091 33473
rect 57790 33464 57796 33516
rect 57848 33504 57854 33516
rect 58345 33507 58403 33513
rect 58345 33504 58357 33507
rect 57848 33476 58357 33504
rect 57848 33464 57854 33476
rect 58345 33473 58357 33476
rect 58391 33473 58403 33507
rect 58345 33467 58403 33473
rect 54754 33436 54760 33448
rect 54715 33408 54760 33436
rect 54754 33396 54760 33408
rect 54812 33396 54818 33448
rect 56870 33260 56876 33312
rect 56928 33300 56934 33312
rect 58161 33303 58219 33309
rect 58161 33300 58173 33303
rect 56928 33272 58173 33300
rect 56928 33260 56934 33272
rect 58161 33269 58173 33272
rect 58207 33269 58219 33303
rect 58161 33263 58219 33269
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 48498 32988 48504 33040
rect 48556 33028 48562 33040
rect 56413 33031 56471 33037
rect 56413 33028 56425 33031
rect 48556 33000 56425 33028
rect 48556 32988 48562 33000
rect 56413 32997 56425 33000
rect 56459 32997 56471 33031
rect 56413 32991 56471 32997
rect 1857 32895 1915 32901
rect 1857 32861 1869 32895
rect 1903 32892 1915 32895
rect 1903 32864 2452 32892
rect 1903 32861 1915 32864
rect 1857 32855 1915 32861
rect 1670 32756 1676 32768
rect 1631 32728 1676 32756
rect 1670 32716 1676 32728
rect 1728 32716 1734 32768
rect 2424 32765 2452 32864
rect 56410 32852 56416 32904
rect 56468 32892 56474 32904
rect 56704 32892 56732 32946
rect 56962 32892 56968 32904
rect 56468 32864 56732 32892
rect 56923 32864 56968 32892
rect 56468 32852 56474 32864
rect 56962 32852 56968 32864
rect 57020 32852 57026 32904
rect 57425 32895 57483 32901
rect 57425 32861 57437 32895
rect 57471 32892 57483 32895
rect 57974 32892 57980 32904
rect 57471 32864 57980 32892
rect 57471 32861 57483 32864
rect 57425 32855 57483 32861
rect 57974 32852 57980 32864
rect 58032 32852 58038 32904
rect 56778 32784 56784 32836
rect 56836 32824 56842 32836
rect 57333 32827 57391 32833
rect 56836 32796 57284 32824
rect 56836 32784 56842 32796
rect 2409 32759 2467 32765
rect 2409 32725 2421 32759
rect 2455 32756 2467 32759
rect 2682 32756 2688 32768
rect 2455 32728 2688 32756
rect 2455 32725 2467 32728
rect 2409 32719 2467 32725
rect 2682 32716 2688 32728
rect 2740 32716 2746 32768
rect 55766 32756 55772 32768
rect 55727 32728 55772 32756
rect 55766 32716 55772 32728
rect 55824 32716 55830 32768
rect 56597 32759 56655 32765
rect 56597 32725 56609 32759
rect 56643 32756 56655 32759
rect 57054 32756 57060 32768
rect 56643 32728 57060 32756
rect 56643 32725 56655 32728
rect 56597 32719 56655 32725
rect 57054 32716 57060 32728
rect 57112 32716 57118 32768
rect 57256 32756 57284 32796
rect 57333 32793 57345 32827
rect 57379 32824 57391 32827
rect 57514 32824 57520 32836
rect 57379 32796 57520 32824
rect 57379 32793 57391 32796
rect 57333 32787 57391 32793
rect 57514 32784 57520 32796
rect 57572 32784 57578 32836
rect 57701 32759 57759 32765
rect 57701 32756 57713 32759
rect 57256 32728 57713 32756
rect 57701 32725 57713 32728
rect 57747 32725 57759 32759
rect 57701 32719 57759 32725
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 55766 32512 55772 32564
rect 55824 32552 55830 32564
rect 57514 32552 57520 32564
rect 55824 32524 57520 32552
rect 55824 32512 55830 32524
rect 57514 32512 57520 32524
rect 57572 32512 57578 32564
rect 1857 32419 1915 32425
rect 1857 32385 1869 32419
rect 1903 32416 1915 32419
rect 2409 32419 2467 32425
rect 2409 32416 2421 32419
rect 1903 32388 2421 32416
rect 1903 32385 1915 32388
rect 1857 32379 1915 32385
rect 2409 32385 2421 32388
rect 2455 32416 2467 32419
rect 12434 32416 12440 32428
rect 2455 32388 12440 32416
rect 2455 32385 2467 32388
rect 2409 32379 2467 32385
rect 12434 32376 12440 32388
rect 12492 32376 12498 32428
rect 57517 32419 57575 32425
rect 57517 32385 57529 32419
rect 57563 32416 57575 32419
rect 58342 32416 58348 32428
rect 57563 32388 58348 32416
rect 57563 32385 57575 32388
rect 57517 32379 57575 32385
rect 58342 32376 58348 32388
rect 58400 32376 58406 32428
rect 1670 32212 1676 32224
rect 1631 32184 1676 32212
rect 1670 32172 1676 32184
rect 1728 32172 1734 32224
rect 56229 32215 56287 32221
rect 56229 32181 56241 32215
rect 56275 32212 56287 32215
rect 56410 32212 56416 32224
rect 56275 32184 56416 32212
rect 56275 32181 56287 32184
rect 56229 32175 56287 32181
rect 56410 32172 56416 32184
rect 56468 32212 56474 32224
rect 57422 32212 57428 32224
rect 56468 32184 57428 32212
rect 56468 32172 56474 32184
rect 57422 32172 57428 32184
rect 57480 32172 57486 32224
rect 58161 32215 58219 32221
rect 58161 32181 58173 32215
rect 58207 32212 58219 32215
rect 58250 32212 58256 32224
rect 58207 32184 58256 32212
rect 58207 32181 58219 32184
rect 58161 32175 58219 32181
rect 58250 32172 58256 32184
rect 58308 32172 58314 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 56962 31968 56968 32020
rect 57020 32008 57026 32020
rect 59354 32008 59360 32020
rect 57020 31980 59360 32008
rect 57020 31968 57026 31980
rect 59354 31968 59360 31980
rect 59412 31968 59418 32020
rect 55766 31940 55772 31952
rect 55679 31912 55772 31940
rect 55766 31900 55772 31912
rect 55824 31940 55830 31952
rect 56226 31940 56232 31952
rect 55824 31912 56232 31940
rect 55824 31900 55830 31912
rect 56226 31900 56232 31912
rect 56284 31900 56290 31952
rect 57514 31940 57520 31952
rect 57348 31912 57520 31940
rect 56244 31872 56272 31900
rect 56873 31875 56931 31881
rect 56873 31872 56885 31875
rect 56244 31844 56885 31872
rect 56873 31841 56885 31844
rect 56919 31841 56931 31875
rect 56873 31835 56931 31841
rect 56962 31832 56968 31884
rect 57020 31881 57026 31884
rect 57020 31875 57069 31881
rect 57020 31841 57023 31875
rect 57057 31841 57069 31875
rect 57020 31835 57069 31841
rect 57149 31875 57207 31881
rect 57149 31841 57161 31875
rect 57195 31872 57207 31875
rect 57348 31872 57376 31912
rect 57514 31900 57520 31912
rect 57572 31940 57578 31952
rect 58894 31940 58900 31952
rect 57572 31912 58900 31940
rect 57572 31900 57578 31912
rect 58894 31900 58900 31912
rect 58952 31900 58958 31952
rect 57195 31844 57376 31872
rect 57195 31841 57207 31844
rect 57149 31835 57207 31841
rect 57020 31832 57026 31835
rect 57422 31832 57428 31884
rect 57480 31872 57486 31884
rect 58069 31875 58127 31881
rect 57480 31844 57525 31872
rect 57480 31832 57486 31844
rect 58069 31841 58081 31875
rect 58115 31872 58127 31875
rect 58158 31872 58164 31884
rect 58115 31844 58164 31872
rect 58115 31841 58127 31844
rect 58069 31835 58127 31841
rect 58158 31832 58164 31844
rect 58216 31832 58222 31884
rect 54478 31764 54484 31816
rect 54536 31804 54542 31816
rect 56229 31807 56287 31813
rect 56229 31804 56241 31807
rect 54536 31776 56241 31804
rect 54536 31764 54542 31776
rect 56229 31773 56241 31776
rect 56275 31773 56287 31807
rect 56229 31767 56287 31773
rect 57885 31807 57943 31813
rect 57885 31773 57897 31807
rect 57931 31804 57943 31807
rect 57974 31804 57980 31816
rect 57931 31776 57980 31804
rect 57931 31773 57943 31776
rect 57885 31767 57943 31773
rect 57974 31764 57980 31776
rect 58032 31764 58038 31816
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 57514 31464 57520 31476
rect 57475 31436 57520 31464
rect 57514 31424 57520 31436
rect 57572 31424 57578 31476
rect 56962 31356 56968 31408
rect 57020 31396 57026 31408
rect 59078 31396 59084 31408
rect 57020 31368 59084 31396
rect 57020 31356 57026 31368
rect 59078 31356 59084 31368
rect 59136 31356 59142 31408
rect 1857 31331 1915 31337
rect 1857 31297 1869 31331
rect 1903 31328 1915 31331
rect 2222 31328 2228 31340
rect 1903 31300 2228 31328
rect 1903 31297 1915 31300
rect 1857 31291 1915 31297
rect 2222 31288 2228 31300
rect 2280 31288 2286 31340
rect 53745 31331 53803 31337
rect 53745 31297 53757 31331
rect 53791 31328 53803 31331
rect 54478 31328 54484 31340
rect 53791 31300 54484 31328
rect 53791 31297 53803 31300
rect 53745 31291 53803 31297
rect 54478 31288 54484 31300
rect 54536 31288 54542 31340
rect 58158 31328 58164 31340
rect 58119 31300 58164 31328
rect 58158 31288 58164 31300
rect 58216 31288 58222 31340
rect 49050 31220 49056 31272
rect 49108 31260 49114 31272
rect 53469 31263 53527 31269
rect 53469 31260 53481 31263
rect 49108 31232 53481 31260
rect 49108 31220 49114 31232
rect 53469 31229 53481 31232
rect 53515 31229 53527 31263
rect 53469 31223 53527 31229
rect 1670 31192 1676 31204
rect 1631 31164 1676 31192
rect 1670 31152 1676 31164
rect 1728 31152 1734 31204
rect 2222 31084 2228 31136
rect 2280 31124 2286 31136
rect 2317 31127 2375 31133
rect 2317 31124 2329 31127
rect 2280 31096 2329 31124
rect 2280 31084 2286 31096
rect 2317 31093 2329 31096
rect 2363 31093 2375 31127
rect 2317 31087 2375 31093
rect 56137 31127 56195 31133
rect 56137 31093 56149 31127
rect 56183 31124 56195 31127
rect 56410 31124 56416 31136
rect 56183 31096 56416 31124
rect 56183 31093 56195 31096
rect 56137 31087 56195 31093
rect 56410 31084 56416 31096
rect 56468 31084 56474 31136
rect 58345 31127 58403 31133
rect 58345 31093 58357 31127
rect 58391 31124 58403 31127
rect 58526 31124 58532 31136
rect 58391 31096 58532 31124
rect 58391 31093 58403 31096
rect 58345 31087 58403 31093
rect 58526 31084 58532 31096
rect 58584 31084 58590 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 57701 30923 57759 30929
rect 57701 30889 57713 30923
rect 57747 30920 57759 30923
rect 58158 30920 58164 30932
rect 57747 30892 58164 30920
rect 57747 30889 57759 30892
rect 57701 30883 57759 30889
rect 58158 30880 58164 30892
rect 58216 30880 58222 30932
rect 57514 30812 57520 30864
rect 57572 30852 57578 30864
rect 58434 30852 58440 30864
rect 57572 30824 58440 30852
rect 57572 30812 57578 30824
rect 58434 30812 58440 30824
rect 58492 30812 58498 30864
rect 1857 30719 1915 30725
rect 1857 30685 1869 30719
rect 1903 30716 1915 30719
rect 58161 30719 58219 30725
rect 1903 30688 2452 30716
rect 1903 30685 1915 30688
rect 1857 30679 1915 30685
rect 2424 30592 2452 30688
rect 58161 30685 58173 30719
rect 58207 30716 58219 30719
rect 58434 30716 58440 30728
rect 58207 30688 58440 30716
rect 58207 30685 58219 30688
rect 58161 30679 58219 30685
rect 58434 30676 58440 30688
rect 58492 30676 58498 30728
rect 1670 30580 1676 30592
rect 1631 30552 1676 30580
rect 1670 30540 1676 30552
rect 1728 30540 1734 30592
rect 2406 30580 2412 30592
rect 2367 30552 2412 30580
rect 2406 30540 2412 30552
rect 2464 30540 2470 30592
rect 58342 30580 58348 30592
rect 58303 30552 58348 30580
rect 58342 30540 58348 30552
rect 58400 30540 58406 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 58345 30379 58403 30385
rect 58345 30345 58357 30379
rect 58391 30376 58403 30379
rect 58434 30376 58440 30388
rect 58391 30348 58440 30376
rect 58391 30345 58403 30348
rect 58345 30339 58403 30345
rect 58434 30336 58440 30348
rect 58492 30336 58498 30388
rect 12161 30311 12219 30317
rect 12161 30277 12173 30311
rect 12207 30308 12219 30311
rect 12434 30308 12440 30320
rect 12207 30280 12440 30308
rect 12207 30277 12219 30280
rect 12161 30271 12219 30277
rect 12434 30268 12440 30280
rect 12492 30308 12498 30320
rect 12618 30308 12624 30320
rect 12492 30280 12624 30308
rect 12492 30268 12498 30280
rect 12618 30268 12624 30280
rect 12676 30308 12682 30320
rect 12897 30311 12955 30317
rect 12897 30308 12909 30311
rect 12676 30280 12909 30308
rect 12676 30268 12682 30280
rect 12897 30277 12909 30280
rect 12943 30277 12955 30311
rect 12897 30271 12955 30277
rect 14458 30268 14464 30320
rect 14516 30308 14522 30320
rect 15654 30308 15660 30320
rect 14516 30280 15660 30308
rect 14516 30268 14522 30280
rect 15654 30268 15660 30280
rect 15712 30268 15718 30320
rect 56962 30308 56968 30320
rect 56923 30280 56968 30308
rect 56962 30268 56968 30280
rect 57020 30268 57026 30320
rect 11054 30200 11060 30252
rect 11112 30240 11118 30252
rect 12069 30243 12127 30249
rect 12069 30240 12081 30243
rect 11112 30212 12081 30240
rect 11112 30200 11118 30212
rect 12069 30209 12081 30212
rect 12115 30209 12127 30243
rect 12069 30203 12127 30209
rect 12342 30172 12348 30184
rect 12303 30144 12348 30172
rect 12342 30132 12348 30144
rect 12400 30132 12406 30184
rect 57146 30132 57152 30184
rect 57204 30172 57210 30184
rect 57606 30172 57612 30184
rect 57204 30144 57612 30172
rect 57204 30132 57210 30144
rect 57606 30132 57612 30144
rect 57664 30132 57670 30184
rect 11054 30036 11060 30048
rect 11015 30008 11060 30036
rect 11054 29996 11060 30008
rect 11112 29996 11118 30048
rect 11422 29996 11428 30048
rect 11480 30036 11486 30048
rect 11701 30039 11759 30045
rect 11701 30036 11713 30039
rect 11480 30008 11713 30036
rect 11480 29996 11486 30008
rect 11701 30005 11713 30008
rect 11747 30005 11759 30039
rect 11701 29999 11759 30005
rect 57146 29996 57152 30048
rect 57204 30036 57210 30048
rect 57422 30036 57428 30048
rect 57204 30008 57428 30036
rect 57204 29996 57210 30008
rect 57422 29996 57428 30008
rect 57480 29996 57486 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 57698 29724 57704 29776
rect 57756 29764 57762 29776
rect 57756 29736 57836 29764
rect 57756 29724 57762 29736
rect 9217 29699 9275 29705
rect 9217 29665 9229 29699
rect 9263 29696 9275 29699
rect 11146 29696 11152 29708
rect 9263 29668 11152 29696
rect 9263 29665 9275 29668
rect 9217 29659 9275 29665
rect 11146 29656 11152 29668
rect 11204 29656 11210 29708
rect 57808 29696 57836 29736
rect 58345 29699 58403 29705
rect 58345 29696 58357 29699
rect 57808 29682 58357 29696
rect 57822 29668 58357 29682
rect 58345 29665 58357 29668
rect 58391 29665 58403 29699
rect 58345 29659 58403 29665
rect 1857 29631 1915 29637
rect 1857 29597 1869 29631
rect 1903 29597 1915 29631
rect 11422 29628 11428 29640
rect 11383 29600 11428 29628
rect 1857 29591 1915 29597
rect 1872 29560 1900 29591
rect 11422 29588 11428 29600
rect 11480 29588 11486 29640
rect 56873 29631 56931 29637
rect 56873 29597 56885 29631
rect 56919 29628 56931 29631
rect 58250 29628 58256 29640
rect 56919 29600 58256 29628
rect 56919 29597 56931 29600
rect 56873 29591 56931 29597
rect 58250 29588 58256 29600
rect 58308 29588 58314 29640
rect 2409 29563 2467 29569
rect 2409 29560 2421 29563
rect 1872 29532 2421 29560
rect 2409 29529 2421 29532
rect 2455 29560 2467 29563
rect 9214 29560 9220 29572
rect 2455 29532 9220 29560
rect 2455 29529 2467 29532
rect 2409 29523 2467 29529
rect 9214 29520 9220 29532
rect 9272 29520 9278 29572
rect 9766 29560 9772 29572
rect 9679 29532 9772 29560
rect 9766 29520 9772 29532
rect 9824 29560 9830 29572
rect 9824 29532 12388 29560
rect 9824 29520 9830 29532
rect 12360 29504 12388 29532
rect 56134 29520 56140 29572
rect 56192 29560 56198 29572
rect 56505 29563 56563 29569
rect 56505 29560 56517 29563
rect 56192 29532 56517 29560
rect 56192 29520 56198 29532
rect 56505 29529 56517 29532
rect 56551 29529 56563 29563
rect 56505 29523 56563 29529
rect 57146 29520 57152 29572
rect 57204 29560 57210 29572
rect 57241 29563 57299 29569
rect 57241 29560 57253 29563
rect 57204 29532 57253 29560
rect 57204 29520 57210 29532
rect 57241 29529 57253 29532
rect 57287 29529 57299 29563
rect 57241 29523 57299 29529
rect 57333 29563 57391 29569
rect 57333 29529 57345 29563
rect 57379 29529 57391 29563
rect 57333 29523 57391 29529
rect 57609 29563 57667 29569
rect 57609 29529 57621 29563
rect 57655 29560 57667 29563
rect 58986 29560 58992 29572
rect 57655 29532 58992 29560
rect 57655 29529 57667 29532
rect 57609 29523 57667 29529
rect 1670 29492 1676 29504
rect 1631 29464 1676 29492
rect 1670 29452 1676 29464
rect 1728 29452 1734 29504
rect 11238 29492 11244 29504
rect 11199 29464 11244 29492
rect 11238 29452 11244 29464
rect 11296 29452 11302 29504
rect 12342 29452 12348 29504
rect 12400 29492 12406 29504
rect 12529 29495 12587 29501
rect 12529 29492 12541 29495
rect 12400 29464 12541 29492
rect 12400 29452 12406 29464
rect 12529 29461 12541 29464
rect 12575 29461 12587 29495
rect 12529 29455 12587 29461
rect 55582 29452 55588 29504
rect 55640 29492 55646 29504
rect 56321 29495 56379 29501
rect 56321 29492 56333 29495
rect 55640 29464 56333 29492
rect 55640 29452 55646 29464
rect 56321 29461 56333 29464
rect 56367 29461 56379 29495
rect 56321 29455 56379 29461
rect 56962 29452 56968 29504
rect 57020 29492 57026 29504
rect 57348 29492 57376 29523
rect 58986 29520 58992 29532
rect 59044 29520 59050 29572
rect 57020 29464 57376 29492
rect 57020 29452 57026 29464
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 8478 29288 8484 29300
rect 8439 29260 8484 29288
rect 8478 29248 8484 29260
rect 8536 29288 8542 29300
rect 9217 29291 9275 29297
rect 9217 29288 9229 29291
rect 8536 29260 9229 29288
rect 8536 29248 8542 29260
rect 9217 29257 9229 29260
rect 9263 29257 9275 29291
rect 9217 29251 9275 29257
rect 10689 29291 10747 29297
rect 10689 29257 10701 29291
rect 10735 29288 10747 29291
rect 10778 29288 10784 29300
rect 10735 29260 10784 29288
rect 10735 29257 10747 29260
rect 10689 29251 10747 29257
rect 10778 29248 10784 29260
rect 10836 29288 10842 29300
rect 11701 29291 11759 29297
rect 11701 29288 11713 29291
rect 10836 29260 11713 29288
rect 10836 29248 10842 29260
rect 11701 29257 11713 29260
rect 11747 29288 11759 29291
rect 11974 29288 11980 29300
rect 11747 29260 11980 29288
rect 11747 29257 11759 29260
rect 11701 29251 11759 29257
rect 11974 29248 11980 29260
rect 12032 29248 12038 29300
rect 57330 29288 57336 29300
rect 57291 29260 57336 29288
rect 57330 29248 57336 29260
rect 57388 29248 57394 29300
rect 57606 29248 57612 29300
rect 57664 29288 57670 29300
rect 58161 29291 58219 29297
rect 58161 29288 58173 29291
rect 57664 29260 58173 29288
rect 57664 29248 57670 29260
rect 58161 29257 58173 29260
rect 58207 29257 58219 29291
rect 58161 29251 58219 29257
rect 2409 29223 2467 29229
rect 2409 29220 2421 29223
rect 1872 29192 2421 29220
rect 1872 29161 1900 29192
rect 2409 29189 2421 29192
rect 2455 29220 2467 29223
rect 15010 29220 15016 29232
rect 2455 29192 15016 29220
rect 2455 29189 2467 29192
rect 2409 29183 2467 29189
rect 15010 29180 15016 29192
rect 15068 29180 15074 29232
rect 56321 29223 56379 29229
rect 56321 29189 56333 29223
rect 56367 29220 56379 29223
rect 56367 29192 58388 29220
rect 56367 29189 56379 29192
rect 56321 29183 56379 29189
rect 1857 29155 1915 29161
rect 1857 29121 1869 29155
rect 1903 29121 1915 29155
rect 1857 29115 1915 29121
rect 8389 29155 8447 29161
rect 8389 29121 8401 29155
rect 8435 29152 8447 29155
rect 10597 29155 10655 29161
rect 10597 29152 10609 29155
rect 8435 29124 10609 29152
rect 8435 29121 8447 29124
rect 8389 29115 8447 29121
rect 10597 29121 10609 29124
rect 10643 29152 10655 29155
rect 11146 29152 11152 29164
rect 10643 29124 11152 29152
rect 10643 29121 10655 29124
rect 10597 29115 10655 29121
rect 11146 29112 11152 29124
rect 11204 29112 11210 29164
rect 58360 29161 58388 29192
rect 57517 29155 57575 29161
rect 57517 29152 57529 29155
rect 57164 29124 57529 29152
rect 7469 29087 7527 29093
rect 7469 29084 7481 29087
rect 6886 29056 7481 29084
rect 1670 29016 1676 29028
rect 1631 28988 1676 29016
rect 1670 28976 1676 28988
rect 1728 28976 1734 29028
rect 5902 28976 5908 29028
rect 5960 29016 5966 29028
rect 6886 29016 6914 29056
rect 7469 29053 7481 29056
rect 7515 29084 7527 29087
rect 8665 29087 8723 29093
rect 8665 29084 8677 29087
rect 7515 29056 8677 29084
rect 7515 29053 7527 29056
rect 7469 29047 7527 29053
rect 8665 29053 8677 29056
rect 8711 29084 8723 29087
rect 9766 29084 9772 29096
rect 8711 29056 9772 29084
rect 8711 29053 8723 29056
rect 8665 29047 8723 29053
rect 9766 29044 9772 29056
rect 9824 29044 9830 29096
rect 10873 29087 10931 29093
rect 10873 29053 10885 29087
rect 10919 29053 10931 29087
rect 10873 29047 10931 29053
rect 5960 28988 6914 29016
rect 5960 28976 5966 28988
rect 9950 28976 9956 29028
rect 10008 29016 10014 29028
rect 10229 29019 10287 29025
rect 10229 29016 10241 29019
rect 10008 28988 10241 29016
rect 10008 28976 10014 28988
rect 10229 28985 10241 28988
rect 10275 28985 10287 29019
rect 10888 29016 10916 29047
rect 57164 29028 57192 29124
rect 57517 29121 57529 29124
rect 57563 29121 57575 29155
rect 57517 29115 57575 29121
rect 58345 29155 58403 29161
rect 58345 29121 58357 29155
rect 58391 29152 58403 29155
rect 58434 29152 58440 29164
rect 58391 29124 58440 29152
rect 58391 29121 58403 29124
rect 58345 29115 58403 29121
rect 58434 29112 58440 29124
rect 58492 29112 58498 29164
rect 10962 29016 10968 29028
rect 10888 28988 10968 29016
rect 10229 28979 10287 28985
rect 10962 28976 10968 28988
rect 11020 29016 11026 29028
rect 12253 29019 12311 29025
rect 12253 29016 12265 29019
rect 11020 28988 12265 29016
rect 11020 28976 11026 28988
rect 12253 28985 12265 28988
rect 12299 28985 12311 29019
rect 12253 28979 12311 28985
rect 56873 29019 56931 29025
rect 56873 28985 56885 29019
rect 56919 29016 56931 29019
rect 57146 29016 57152 29028
rect 56919 28988 57152 29016
rect 56919 28985 56931 28988
rect 56873 28979 56931 28985
rect 57146 28976 57152 28988
rect 57204 28976 57210 29028
rect 6822 28948 6828 28960
rect 6783 28920 6828 28948
rect 6822 28908 6828 28920
rect 6880 28908 6886 28960
rect 7650 28908 7656 28960
rect 7708 28948 7714 28960
rect 8021 28951 8079 28957
rect 8021 28948 8033 28951
rect 7708 28920 8033 28948
rect 7708 28908 7714 28920
rect 8021 28917 8033 28920
rect 8067 28917 8079 28951
rect 8021 28911 8079 28917
rect 56962 28908 56968 28960
rect 57020 28948 57026 28960
rect 57330 28948 57336 28960
rect 57020 28920 57336 28948
rect 57020 28908 57026 28920
rect 57330 28908 57336 28920
rect 57388 28908 57394 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 3786 28704 3792 28756
rect 3844 28744 3850 28756
rect 3844 28716 6914 28744
rect 3844 28704 3850 28716
rect 5902 28608 5908 28620
rect 5863 28580 5908 28608
rect 5902 28568 5908 28580
rect 5960 28568 5966 28620
rect 6886 28608 6914 28716
rect 7926 28704 7932 28756
rect 7984 28744 7990 28756
rect 8573 28747 8631 28753
rect 8573 28744 8585 28747
rect 7984 28716 8585 28744
rect 7984 28704 7990 28716
rect 8573 28713 8585 28716
rect 8619 28744 8631 28747
rect 8619 28716 9720 28744
rect 8619 28713 8631 28716
rect 8573 28707 8631 28713
rect 7837 28679 7895 28685
rect 7837 28645 7849 28679
rect 7883 28676 7895 28679
rect 8754 28676 8760 28688
rect 7883 28648 8760 28676
rect 7883 28645 7895 28648
rect 7837 28639 7895 28645
rect 8754 28636 8760 28648
rect 8812 28636 8818 28688
rect 9582 28608 9588 28620
rect 6886 28580 9444 28608
rect 9543 28580 9588 28608
rect 5994 28500 6000 28552
rect 6052 28540 6058 28552
rect 6181 28543 6239 28549
rect 6181 28540 6193 28543
rect 6052 28512 6193 28540
rect 6052 28500 6058 28512
rect 6181 28509 6193 28512
rect 6227 28540 6239 28543
rect 6822 28540 6828 28552
rect 6227 28512 6828 28540
rect 6227 28509 6239 28512
rect 6181 28503 6239 28509
rect 6822 28500 6828 28512
rect 6880 28500 6886 28552
rect 7650 28540 7656 28552
rect 7611 28512 7656 28540
rect 7650 28500 7656 28512
rect 7708 28500 7714 28552
rect 9416 28540 9444 28580
rect 9582 28568 9588 28580
rect 9640 28568 9646 28620
rect 9692 28617 9720 28716
rect 16574 28704 16580 28756
rect 16632 28744 16638 28756
rect 16632 28716 16677 28744
rect 16632 28704 16638 28716
rect 9766 28636 9772 28688
rect 9824 28676 9830 28688
rect 11793 28679 11851 28685
rect 11793 28676 11805 28679
rect 9824 28648 11805 28676
rect 9824 28636 9830 28648
rect 11793 28645 11805 28648
rect 11839 28645 11851 28679
rect 11793 28639 11851 28645
rect 9677 28611 9735 28617
rect 9677 28577 9689 28611
rect 9723 28608 9735 28611
rect 10962 28608 10968 28620
rect 9723 28580 10968 28608
rect 9723 28577 9735 28580
rect 9677 28571 9735 28577
rect 10962 28568 10968 28580
rect 11020 28568 11026 28620
rect 12342 28608 12348 28620
rect 12303 28580 12348 28608
rect 12342 28568 12348 28580
rect 12400 28568 12406 28620
rect 57698 28568 57704 28620
rect 57756 28568 57762 28620
rect 9490 28540 9496 28552
rect 9403 28512 9496 28540
rect 9490 28500 9496 28512
rect 9548 28500 9554 28552
rect 9600 28540 9628 28568
rect 10321 28543 10379 28549
rect 10321 28540 10333 28543
rect 9600 28512 10333 28540
rect 10321 28509 10333 28512
rect 10367 28540 10379 28543
rect 10502 28540 10508 28552
rect 10367 28512 10508 28540
rect 10367 28509 10379 28512
rect 10321 28503 10379 28509
rect 10502 28500 10508 28512
rect 10560 28500 10566 28552
rect 11698 28500 11704 28552
rect 11756 28540 11762 28552
rect 12253 28543 12311 28549
rect 12253 28540 12265 28543
rect 11756 28512 12265 28540
rect 11756 28500 11762 28512
rect 12253 28509 12265 28512
rect 12299 28509 12311 28543
rect 12253 28503 12311 28509
rect 56045 28543 56103 28549
rect 56045 28509 56057 28543
rect 56091 28540 56103 28543
rect 57149 28543 57207 28549
rect 56091 28512 57008 28540
rect 56091 28509 56103 28512
rect 56045 28503 56103 28509
rect 6089 28475 6147 28481
rect 6089 28441 6101 28475
rect 6135 28472 6147 28475
rect 6914 28472 6920 28484
rect 6135 28444 6920 28472
rect 6135 28441 6147 28444
rect 6089 28435 6147 28441
rect 6914 28432 6920 28444
rect 6972 28472 6978 28484
rect 7009 28475 7067 28481
rect 7009 28472 7021 28475
rect 6972 28444 7021 28472
rect 6972 28432 6978 28444
rect 7009 28441 7021 28444
rect 7055 28472 7067 28475
rect 7098 28472 7104 28484
rect 7055 28444 7104 28472
rect 7055 28441 7067 28444
rect 7009 28435 7067 28441
rect 7098 28432 7104 28444
rect 7156 28432 7162 28484
rect 12989 28475 13047 28481
rect 12989 28472 13001 28475
rect 12176 28444 13001 28472
rect 12176 28416 12204 28444
rect 12989 28441 13001 28444
rect 13035 28441 13047 28475
rect 56980 28472 57008 28512
rect 57149 28509 57161 28543
rect 57195 28540 57207 28543
rect 57330 28540 57336 28552
rect 57195 28512 57336 28540
rect 57195 28509 57207 28512
rect 57149 28503 57207 28509
rect 57330 28500 57336 28512
rect 57388 28500 57394 28552
rect 57422 28500 57428 28552
rect 57480 28540 57486 28552
rect 57517 28543 57575 28549
rect 57517 28540 57529 28543
rect 57480 28512 57529 28540
rect 57480 28500 57486 28512
rect 57517 28509 57529 28512
rect 57563 28509 57575 28543
rect 57517 28503 57575 28509
rect 57609 28543 57667 28549
rect 57609 28509 57621 28543
rect 57655 28540 57667 28543
rect 58710 28540 58716 28552
rect 57655 28512 58716 28540
rect 57655 28509 57667 28512
rect 57609 28503 57667 28509
rect 57624 28472 57652 28503
rect 58710 28500 58716 28512
rect 58768 28500 58774 28552
rect 57882 28472 57888 28484
rect 12989 28435 13047 28441
rect 56612 28444 56916 28472
rect 56980 28444 57652 28472
rect 57843 28444 57888 28472
rect 1946 28404 1952 28416
rect 1907 28376 1952 28404
rect 1946 28364 1952 28376
rect 2004 28364 2010 28416
rect 4062 28364 4068 28416
rect 4120 28404 4126 28416
rect 5261 28407 5319 28413
rect 5261 28404 5273 28407
rect 4120 28376 5273 28404
rect 4120 28364 4126 28376
rect 5261 28373 5273 28376
rect 5307 28373 5319 28407
rect 5261 28367 5319 28373
rect 6549 28407 6607 28413
rect 6549 28373 6561 28407
rect 6595 28404 6607 28407
rect 6822 28404 6828 28416
rect 6595 28376 6828 28404
rect 6595 28373 6607 28376
rect 6549 28367 6607 28373
rect 6822 28364 6828 28376
rect 6880 28364 6886 28416
rect 9122 28404 9128 28416
rect 9083 28376 9128 28404
rect 9122 28364 9128 28376
rect 9180 28364 9186 28416
rect 11146 28364 11152 28416
rect 11204 28404 11210 28416
rect 11241 28407 11299 28413
rect 11241 28404 11253 28407
rect 11204 28376 11253 28404
rect 11204 28364 11210 28376
rect 11241 28373 11253 28376
rect 11287 28373 11299 28407
rect 12158 28404 12164 28416
rect 12119 28376 12164 28404
rect 11241 28367 11299 28373
rect 12158 28364 12164 28376
rect 12216 28364 12222 28416
rect 56612 28413 56640 28444
rect 56597 28407 56655 28413
rect 56597 28373 56609 28407
rect 56643 28373 56655 28407
rect 56778 28404 56784 28416
rect 56739 28376 56784 28404
rect 56597 28367 56655 28373
rect 56778 28364 56784 28376
rect 56836 28364 56842 28416
rect 56888 28404 56916 28444
rect 57882 28432 57888 28444
rect 57940 28432 57946 28484
rect 57330 28404 57336 28416
rect 56888 28376 57336 28404
rect 57330 28364 57336 28376
rect 57388 28364 57394 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 4706 28200 4712 28212
rect 4667 28172 4712 28200
rect 4706 28160 4712 28172
rect 4764 28200 4770 28212
rect 5629 28203 5687 28209
rect 5629 28200 5641 28203
rect 4764 28172 5641 28200
rect 4764 28160 4770 28172
rect 5629 28169 5641 28172
rect 5675 28169 5687 28203
rect 5629 28163 5687 28169
rect 5644 28132 5672 28163
rect 6178 28160 6184 28212
rect 6236 28200 6242 28212
rect 8481 28203 8539 28209
rect 6236 28172 7972 28200
rect 6236 28160 6242 28172
rect 6454 28132 6460 28144
rect 5644 28104 6460 28132
rect 6454 28092 6460 28104
rect 6512 28092 6518 28144
rect 1857 28067 1915 28073
rect 1857 28033 1869 28067
rect 1903 28064 1915 28067
rect 4801 28067 4859 28073
rect 1903 28036 2452 28064
rect 1903 28033 1915 28036
rect 1857 28027 1915 28033
rect 1670 27928 1676 27940
rect 1631 27900 1676 27928
rect 1670 27888 1676 27900
rect 1728 27888 1734 27940
rect 2424 27937 2452 28036
rect 4801 28033 4813 28067
rect 4847 28064 4859 28067
rect 5994 28064 6000 28076
rect 4847 28036 6000 28064
rect 4847 28033 4859 28036
rect 4801 28027 4859 28033
rect 5994 28024 6000 28036
rect 6052 28024 6058 28076
rect 6822 28064 6828 28076
rect 6783 28036 6828 28064
rect 6822 28024 6828 28036
rect 6880 28024 6886 28076
rect 3418 27956 3424 28008
rect 3476 27996 3482 28008
rect 4062 27996 4068 28008
rect 3476 27968 4068 27996
rect 3476 27956 3482 27968
rect 4062 27956 4068 27968
rect 4120 27996 4126 28008
rect 4525 27999 4583 28005
rect 4525 27996 4537 27999
rect 4120 27968 4537 27996
rect 4120 27956 4126 27968
rect 4525 27965 4537 27968
rect 4571 27996 4583 27999
rect 7834 27996 7840 28008
rect 4571 27968 7840 27996
rect 4571 27965 4583 27968
rect 4525 27959 4583 27965
rect 7834 27956 7840 27968
rect 7892 27956 7898 28008
rect 7944 27996 7972 28172
rect 8481 28169 8493 28203
rect 8527 28169 8539 28203
rect 8481 28163 8539 28169
rect 9125 28203 9183 28209
rect 9125 28169 9137 28203
rect 9171 28200 9183 28203
rect 12066 28200 12072 28212
rect 9171 28172 12072 28200
rect 9171 28169 9183 28172
rect 9125 28163 9183 28169
rect 8110 28064 8116 28076
rect 8071 28036 8116 28064
rect 8110 28024 8116 28036
rect 8168 28024 8174 28076
rect 8496 28064 8524 28163
rect 12066 28160 12072 28172
rect 12124 28160 12130 28212
rect 12342 28160 12348 28212
rect 12400 28200 12406 28212
rect 12713 28203 12771 28209
rect 12713 28200 12725 28203
rect 12400 28172 12725 28200
rect 12400 28160 12406 28172
rect 12713 28169 12725 28172
rect 12759 28200 12771 28203
rect 56965 28203 57023 28209
rect 12759 28172 17540 28200
rect 12759 28169 12771 28172
rect 12713 28163 12771 28169
rect 9490 28092 9496 28144
rect 9548 28132 9554 28144
rect 10137 28135 10195 28141
rect 10137 28132 10149 28135
rect 9548 28104 10149 28132
rect 9548 28092 9554 28104
rect 10137 28101 10149 28104
rect 10183 28132 10195 28135
rect 11054 28132 11060 28144
rect 10183 28104 11060 28132
rect 10183 28101 10195 28104
rect 10137 28095 10195 28101
rect 11054 28092 11060 28104
rect 11112 28092 11118 28144
rect 11422 28092 11428 28144
rect 11480 28132 11486 28144
rect 11698 28132 11704 28144
rect 11480 28104 11704 28132
rect 11480 28092 11486 28104
rect 11698 28092 11704 28104
rect 11756 28092 11762 28144
rect 16574 28092 16580 28144
rect 16632 28132 16638 28144
rect 17313 28135 17371 28141
rect 17313 28132 17325 28135
rect 16632 28104 17325 28132
rect 16632 28092 16638 28104
rect 17313 28101 17325 28104
rect 17359 28101 17371 28135
rect 17313 28095 17371 28101
rect 8941 28067 8999 28073
rect 8941 28064 8953 28067
rect 8496 28036 8953 28064
rect 8941 28033 8953 28036
rect 8987 28033 8999 28067
rect 8941 28027 8999 28033
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28064 15991 28067
rect 17218 28064 17224 28076
rect 15979 28036 16574 28064
rect 17179 28036 17224 28064
rect 15979 28033 15991 28036
rect 15933 28027 15991 28033
rect 8021 27999 8079 28005
rect 8021 27996 8033 27999
rect 7944 27968 8033 27996
rect 8021 27965 8033 27968
rect 8067 27996 8079 27999
rect 8067 27968 9720 27996
rect 8067 27965 8079 27968
rect 8021 27959 8079 27965
rect 2409 27931 2467 27937
rect 2409 27897 2421 27931
rect 2455 27928 2467 27931
rect 5258 27928 5264 27940
rect 2455 27900 5264 27928
rect 2455 27897 2467 27900
rect 2409 27891 2467 27897
rect 5258 27888 5264 27900
rect 5316 27888 5322 27940
rect 9692 27872 9720 27968
rect 16546 27928 16574 28036
rect 17218 28024 17224 28036
rect 17276 28024 17282 28076
rect 17512 28005 17540 28172
rect 56965 28169 56977 28203
rect 57011 28200 57023 28203
rect 57146 28200 57152 28212
rect 57011 28172 57152 28200
rect 57011 28169 57023 28172
rect 56965 28163 57023 28169
rect 57146 28160 57152 28172
rect 57204 28200 57210 28212
rect 57422 28200 57428 28212
rect 57204 28172 57428 28200
rect 57204 28160 57210 28172
rect 57422 28160 57428 28172
rect 57480 28160 57486 28212
rect 57517 28203 57575 28209
rect 57517 28169 57529 28203
rect 57563 28200 57575 28203
rect 57698 28200 57704 28212
rect 57563 28172 57704 28200
rect 57563 28169 57575 28172
rect 57517 28163 57575 28169
rect 57698 28160 57704 28172
rect 57756 28160 57762 28212
rect 56778 28092 56784 28144
rect 56836 28132 56842 28144
rect 58710 28132 58716 28144
rect 56836 28104 58716 28132
rect 56836 28092 56842 28104
rect 58710 28092 58716 28104
rect 58768 28092 58774 28144
rect 56413 28067 56471 28073
rect 56413 28033 56425 28067
rect 56459 28064 56471 28067
rect 58345 28067 58403 28073
rect 58345 28064 58357 28067
rect 56459 28036 58357 28064
rect 56459 28033 56471 28036
rect 56413 28027 56471 28033
rect 58345 28033 58357 28036
rect 58391 28064 58403 28067
rect 58434 28064 58440 28076
rect 58391 28036 58440 28064
rect 58391 28033 58403 28036
rect 58345 28027 58403 28033
rect 58434 28024 58440 28036
rect 58492 28024 58498 28076
rect 17497 27999 17555 28005
rect 17497 27965 17509 27999
rect 17543 27996 17555 27999
rect 17543 27968 18184 27996
rect 17543 27965 17555 27968
rect 17497 27959 17555 27965
rect 16853 27931 16911 27937
rect 16853 27928 16865 27931
rect 16546 27900 16865 27928
rect 16853 27897 16865 27900
rect 16899 27897 16911 27931
rect 16853 27891 16911 27897
rect 2774 27820 2780 27872
rect 2832 27860 2838 27872
rect 3418 27860 3424 27872
rect 2832 27832 3424 27860
rect 2832 27820 2838 27832
rect 3418 27820 3424 27832
rect 3476 27820 3482 27872
rect 5166 27860 5172 27872
rect 5127 27832 5172 27860
rect 5166 27820 5172 27832
rect 5224 27820 5230 27872
rect 7009 27863 7067 27869
rect 7009 27829 7021 27863
rect 7055 27860 7067 27863
rect 8570 27860 8576 27872
rect 7055 27832 8576 27860
rect 7055 27829 7067 27832
rect 7009 27823 7067 27829
rect 8570 27820 8576 27832
rect 8628 27820 8634 27872
rect 9674 27860 9680 27872
rect 9635 27832 9680 27860
rect 9674 27820 9680 27832
rect 9732 27820 9738 27872
rect 10781 27863 10839 27869
rect 10781 27829 10793 27863
rect 10827 27860 10839 27863
rect 10962 27860 10968 27872
rect 10827 27832 10968 27860
rect 10827 27829 10839 27832
rect 10781 27823 10839 27829
rect 10962 27820 10968 27832
rect 11020 27820 11026 27872
rect 13538 27860 13544 27872
rect 13499 27832 13544 27860
rect 13538 27820 13544 27832
rect 13596 27820 13602 27872
rect 15746 27860 15752 27872
rect 15707 27832 15752 27860
rect 15746 27820 15752 27832
rect 15804 27820 15810 27872
rect 18156 27869 18184 27968
rect 54846 27888 54852 27940
rect 54904 27928 54910 27940
rect 58161 27931 58219 27937
rect 58161 27928 58173 27931
rect 54904 27900 58173 27928
rect 54904 27888 54910 27900
rect 58161 27897 58173 27900
rect 58207 27897 58219 27931
rect 58161 27891 58219 27897
rect 18141 27863 18199 27869
rect 18141 27829 18153 27863
rect 18187 27860 18199 27863
rect 19426 27860 19432 27872
rect 18187 27832 19432 27860
rect 18187 27829 18199 27832
rect 18141 27823 18199 27829
rect 19426 27820 19432 27832
rect 19484 27820 19490 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 5905 27659 5963 27665
rect 5905 27625 5917 27659
rect 5951 27656 5963 27659
rect 5994 27656 6000 27668
rect 5951 27628 6000 27656
rect 5951 27625 5963 27628
rect 5905 27619 5963 27625
rect 5994 27616 6000 27628
rect 6052 27616 6058 27668
rect 8110 27588 8116 27600
rect 6886 27560 8116 27588
rect 2774 27520 2780 27532
rect 2735 27492 2780 27520
rect 2774 27480 2780 27492
rect 2832 27480 2838 27532
rect 2869 27523 2927 27529
rect 2869 27489 2881 27523
rect 2915 27520 2927 27523
rect 3050 27520 3056 27532
rect 2915 27492 3056 27520
rect 2915 27489 2927 27492
rect 2869 27483 2927 27489
rect 3050 27480 3056 27492
rect 3108 27520 3114 27532
rect 3973 27523 4031 27529
rect 3973 27520 3985 27523
rect 3108 27492 3985 27520
rect 3108 27480 3114 27492
rect 3973 27489 3985 27492
rect 4019 27520 4031 27523
rect 4062 27520 4068 27532
rect 4019 27492 4068 27520
rect 4019 27489 4031 27492
rect 3973 27483 4031 27489
rect 4062 27480 4068 27492
rect 4120 27480 4126 27532
rect 6886 27520 6914 27560
rect 8110 27548 8116 27560
rect 8168 27588 8174 27600
rect 9125 27591 9183 27597
rect 9125 27588 9137 27591
rect 8168 27560 9137 27588
rect 8168 27548 8174 27560
rect 9125 27557 9137 27560
rect 9171 27557 9183 27591
rect 9125 27551 9183 27557
rect 10410 27548 10416 27600
rect 10468 27588 10474 27600
rect 13538 27588 13544 27600
rect 10468 27560 13544 27588
rect 10468 27548 10474 27560
rect 11149 27523 11207 27529
rect 11149 27520 11161 27523
rect 4172 27492 6914 27520
rect 10152 27492 11161 27520
rect 1857 27455 1915 27461
rect 1857 27421 1869 27455
rect 1903 27452 1915 27455
rect 1946 27452 1952 27464
rect 1903 27424 1952 27452
rect 1903 27421 1915 27424
rect 1857 27415 1915 27421
rect 1946 27412 1952 27424
rect 2004 27412 2010 27464
rect 2038 27412 2044 27464
rect 2096 27452 2102 27464
rect 2096 27424 3372 27452
rect 2096 27412 2102 27424
rect 2961 27387 3019 27393
rect 2961 27353 2973 27387
rect 3007 27384 3019 27387
rect 3234 27384 3240 27396
rect 3007 27356 3240 27384
rect 3007 27353 3019 27356
rect 2961 27347 3019 27353
rect 3234 27344 3240 27356
rect 3292 27344 3298 27396
rect 3344 27384 3372 27424
rect 3878 27412 3884 27464
rect 3936 27452 3942 27464
rect 4172 27452 4200 27492
rect 5166 27452 5172 27464
rect 3936 27424 4200 27452
rect 5127 27424 5172 27452
rect 3936 27412 3942 27424
rect 5166 27412 5172 27424
rect 5224 27412 5230 27464
rect 5350 27412 5356 27464
rect 5408 27452 5414 27464
rect 6365 27455 6423 27461
rect 6365 27452 6377 27455
rect 5408 27424 6377 27452
rect 5408 27412 5414 27424
rect 6365 27421 6377 27424
rect 6411 27421 6423 27455
rect 6365 27415 6423 27421
rect 8205 27455 8263 27461
rect 8205 27421 8217 27455
rect 8251 27452 8263 27455
rect 9122 27452 9128 27464
rect 8251 27424 9128 27452
rect 8251 27421 8263 27424
rect 8205 27415 8263 27421
rect 9122 27412 9128 27424
rect 9180 27412 9186 27464
rect 9858 27384 9864 27396
rect 3344 27356 9864 27384
rect 9858 27344 9864 27356
rect 9916 27384 9922 27396
rect 10152 27393 10180 27492
rect 11149 27489 11161 27492
rect 11195 27489 11207 27523
rect 11330 27520 11336 27532
rect 11291 27492 11336 27520
rect 11149 27483 11207 27489
rect 11330 27480 11336 27492
rect 11388 27480 11394 27532
rect 13280 27529 13308 27560
rect 13538 27548 13544 27560
rect 13596 27548 13602 27600
rect 57698 27588 57704 27600
rect 57659 27560 57704 27588
rect 57698 27548 57704 27560
rect 57756 27548 57762 27600
rect 13265 27523 13323 27529
rect 13265 27489 13277 27523
rect 13311 27489 13323 27523
rect 13556 27520 13584 27548
rect 14829 27523 14887 27529
rect 14829 27520 14841 27523
rect 13556 27492 14841 27520
rect 13265 27483 13323 27489
rect 14829 27489 14841 27492
rect 14875 27520 14887 27523
rect 15102 27520 15108 27532
rect 14875 27492 15108 27520
rect 14875 27489 14887 27492
rect 14829 27483 14887 27489
rect 15102 27480 15108 27492
rect 15160 27480 15166 27532
rect 57146 27520 57152 27532
rect 57107 27492 57152 27520
rect 57146 27480 57152 27492
rect 57204 27480 57210 27532
rect 57238 27480 57244 27532
rect 57296 27529 57302 27532
rect 57296 27523 57345 27529
rect 57296 27489 57299 27523
rect 57333 27489 57345 27523
rect 57296 27483 57345 27489
rect 57425 27523 57483 27529
rect 57425 27489 57437 27523
rect 57471 27520 57483 27523
rect 57606 27520 57612 27532
rect 57471 27492 57612 27520
rect 57471 27489 57483 27492
rect 57425 27483 57483 27489
rect 57296 27480 57302 27483
rect 57606 27480 57612 27492
rect 57664 27480 57670 27532
rect 58342 27520 58348 27532
rect 58303 27492 58348 27520
rect 58342 27480 58348 27492
rect 58400 27480 58406 27532
rect 11054 27412 11060 27464
rect 11112 27452 11118 27464
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 11112 27424 14657 27452
rect 11112 27412 11118 27424
rect 14645 27421 14657 27424
rect 14691 27452 14703 27455
rect 16025 27455 16083 27461
rect 16025 27452 16037 27455
rect 14691 27424 16037 27452
rect 14691 27421 14703 27424
rect 14645 27415 14703 27421
rect 16025 27421 16037 27424
rect 16071 27452 16083 27455
rect 58158 27452 58164 27464
rect 16071 27424 16574 27452
rect 58119 27424 58164 27452
rect 16071 27421 16083 27424
rect 16025 27415 16083 27421
rect 10137 27387 10195 27393
rect 10137 27384 10149 27387
rect 9916 27356 10149 27384
rect 9916 27344 9922 27356
rect 10137 27353 10149 27356
rect 10183 27353 10195 27387
rect 10137 27347 10195 27353
rect 10778 27344 10784 27396
rect 10836 27384 10842 27396
rect 12161 27387 12219 27393
rect 12161 27384 12173 27387
rect 10836 27356 12173 27384
rect 10836 27344 10842 27356
rect 12161 27353 12173 27356
rect 12207 27384 12219 27387
rect 13173 27387 13231 27393
rect 13173 27384 13185 27387
rect 12207 27356 13185 27384
rect 12207 27353 12219 27356
rect 12161 27347 12219 27353
rect 13173 27353 13185 27356
rect 13219 27353 13231 27387
rect 16546 27384 16574 27424
rect 58158 27412 58164 27424
rect 58216 27412 58222 27464
rect 16761 27387 16819 27393
rect 16761 27384 16773 27387
rect 16546 27356 16773 27384
rect 13173 27347 13231 27353
rect 16761 27353 16773 27356
rect 16807 27384 16819 27387
rect 17218 27384 17224 27396
rect 16807 27356 17224 27384
rect 16807 27353 16819 27356
rect 16761 27347 16819 27353
rect 17218 27344 17224 27356
rect 17276 27384 17282 27396
rect 19242 27384 19248 27396
rect 17276 27356 19248 27384
rect 17276 27344 17282 27356
rect 19242 27344 19248 27356
rect 19300 27344 19306 27396
rect 1670 27316 1676 27328
rect 1631 27288 1676 27316
rect 1670 27276 1676 27288
rect 1728 27276 1734 27328
rect 3326 27316 3332 27328
rect 3287 27288 3332 27316
rect 3326 27276 3332 27288
rect 3384 27276 3390 27328
rect 5353 27319 5411 27325
rect 5353 27285 5365 27319
rect 5399 27316 5411 27319
rect 5442 27316 5448 27328
rect 5399 27288 5448 27316
rect 5399 27285 5411 27288
rect 5353 27279 5411 27285
rect 5442 27276 5448 27288
rect 5500 27276 5506 27328
rect 8389 27319 8447 27325
rect 8389 27285 8401 27319
rect 8435 27316 8447 27319
rect 9030 27316 9036 27328
rect 8435 27288 9036 27316
rect 8435 27285 8447 27288
rect 8389 27279 8447 27285
rect 9030 27276 9036 27288
rect 9088 27276 9094 27328
rect 10689 27319 10747 27325
rect 10689 27285 10701 27319
rect 10735 27316 10747 27319
rect 10870 27316 10876 27328
rect 10735 27288 10876 27316
rect 10735 27285 10747 27288
rect 10689 27279 10747 27285
rect 10870 27276 10876 27288
rect 10928 27276 10934 27328
rect 11054 27316 11060 27328
rect 11015 27288 11060 27316
rect 11054 27276 11060 27288
rect 11112 27276 11118 27328
rect 12250 27276 12256 27328
rect 12308 27316 12314 27328
rect 12713 27319 12771 27325
rect 12713 27316 12725 27319
rect 12308 27288 12725 27316
rect 12308 27276 12314 27288
rect 12713 27285 12725 27288
rect 12759 27285 12771 27319
rect 12713 27279 12771 27285
rect 12986 27276 12992 27328
rect 13044 27316 13050 27328
rect 13081 27319 13139 27325
rect 13081 27316 13093 27319
rect 13044 27288 13093 27316
rect 13044 27276 13050 27288
rect 13081 27285 13093 27288
rect 13127 27285 13139 27319
rect 14274 27316 14280 27328
rect 14235 27288 14280 27316
rect 13081 27279 13139 27285
rect 14274 27276 14280 27288
rect 14332 27276 14338 27328
rect 14737 27319 14795 27325
rect 14737 27285 14749 27319
rect 14783 27316 14795 27319
rect 14918 27316 14924 27328
rect 14783 27288 14924 27316
rect 14783 27285 14795 27288
rect 14737 27279 14795 27285
rect 14918 27276 14924 27288
rect 14976 27316 14982 27328
rect 15473 27319 15531 27325
rect 15473 27316 15485 27319
rect 14976 27288 15485 27316
rect 14976 27276 14982 27288
rect 15473 27285 15485 27288
rect 15519 27285 15531 27319
rect 15473 27279 15531 27285
rect 17865 27319 17923 27325
rect 17865 27285 17877 27319
rect 17911 27316 17923 27319
rect 18046 27316 18052 27328
rect 17911 27288 18052 27316
rect 17911 27285 17923 27288
rect 17865 27279 17923 27285
rect 18046 27276 18052 27288
rect 18104 27276 18110 27328
rect 56502 27316 56508 27328
rect 56463 27288 56508 27316
rect 56502 27276 56508 27288
rect 56560 27276 56566 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 2314 27072 2320 27124
rect 2372 27112 2378 27124
rect 5537 27115 5595 27121
rect 5537 27112 5549 27115
rect 2372 27084 5549 27112
rect 2372 27072 2378 27084
rect 5537 27081 5549 27084
rect 5583 27112 5595 27115
rect 6549 27115 6607 27121
rect 6549 27112 6561 27115
rect 5583 27084 6561 27112
rect 5583 27081 5595 27084
rect 5537 27075 5595 27081
rect 6549 27081 6561 27084
rect 6595 27112 6607 27115
rect 6638 27112 6644 27124
rect 6595 27084 6644 27112
rect 6595 27081 6607 27084
rect 6549 27075 6607 27081
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 11054 27072 11060 27124
rect 11112 27112 11118 27124
rect 11701 27115 11759 27121
rect 11701 27112 11713 27115
rect 11112 27084 11713 27112
rect 11112 27072 11118 27084
rect 11701 27081 11713 27084
rect 11747 27081 11759 27115
rect 15102 27112 15108 27124
rect 15063 27084 15108 27112
rect 11701 27075 11759 27081
rect 15102 27072 15108 27084
rect 15160 27112 15166 27124
rect 18230 27112 18236 27124
rect 15160 27084 18236 27112
rect 15160 27072 15166 27084
rect 18230 27072 18236 27084
rect 18288 27072 18294 27124
rect 56965 27115 57023 27121
rect 56965 27081 56977 27115
rect 57011 27112 57023 27115
rect 57146 27112 57152 27124
rect 57011 27084 57152 27112
rect 57011 27081 57023 27084
rect 56965 27075 57023 27081
rect 57146 27072 57152 27084
rect 57204 27072 57210 27124
rect 57517 27115 57575 27121
rect 57517 27081 57529 27115
rect 57563 27112 57575 27115
rect 57698 27112 57704 27124
rect 57563 27084 57704 27112
rect 57563 27081 57575 27084
rect 57517 27075 57575 27081
rect 57698 27072 57704 27084
rect 57756 27072 57762 27124
rect 58161 27115 58219 27121
rect 58161 27081 58173 27115
rect 58207 27112 58219 27115
rect 59446 27112 59452 27124
rect 58207 27084 59452 27112
rect 58207 27081 58219 27084
rect 58161 27075 58219 27081
rect 59446 27072 59452 27084
rect 59504 27072 59510 27124
rect 1673 27047 1731 27053
rect 1673 27013 1685 27047
rect 1719 27044 1731 27047
rect 5810 27044 5816 27056
rect 1719 27016 5816 27044
rect 1719 27013 1731 27016
rect 1673 27007 1731 27013
rect 2240 26976 2268 27016
rect 5810 27004 5816 27016
rect 5868 27004 5874 27056
rect 10962 27004 10968 27056
rect 11020 27044 11026 27056
rect 11149 27047 11207 27053
rect 11149 27044 11161 27047
rect 11020 27016 11161 27044
rect 11020 27004 11026 27016
rect 11149 27013 11161 27016
rect 11195 27044 11207 27047
rect 11330 27044 11336 27056
rect 11195 27016 11336 27044
rect 11195 27013 11207 27016
rect 11149 27007 11207 27013
rect 11330 27004 11336 27016
rect 11388 27044 11394 27056
rect 18046 27044 18052 27056
rect 11388 27016 18052 27044
rect 11388 27004 11394 27016
rect 18046 27004 18052 27016
rect 18104 27004 18110 27056
rect 2314 26976 2320 26988
rect 2240 26948 2320 26976
rect 2240 26917 2268 26948
rect 2314 26936 2320 26948
rect 2372 26936 2378 26988
rect 2501 26979 2559 26985
rect 2501 26945 2513 26979
rect 2547 26976 2559 26979
rect 3234 26976 3240 26988
rect 2547 26948 3240 26976
rect 2547 26945 2559 26948
rect 2501 26939 2559 26945
rect 3234 26936 3240 26948
rect 3292 26936 3298 26988
rect 3326 26936 3332 26988
rect 3384 26976 3390 26988
rect 4157 26979 4215 26985
rect 4157 26976 4169 26979
rect 3384 26948 4169 26976
rect 3384 26936 3390 26948
rect 4157 26945 4169 26948
rect 4203 26945 4215 26979
rect 4157 26939 4215 26945
rect 4798 26936 4804 26988
rect 4856 26976 4862 26988
rect 5629 26979 5687 26985
rect 5629 26976 5641 26979
rect 4856 26948 5641 26976
rect 4856 26936 4862 26948
rect 5629 26945 5641 26948
rect 5675 26976 5687 26979
rect 7101 26979 7159 26985
rect 7101 26976 7113 26979
rect 5675 26948 7113 26976
rect 5675 26945 5687 26948
rect 5629 26939 5687 26945
rect 7101 26945 7113 26948
rect 7147 26945 7159 26979
rect 7101 26939 7159 26945
rect 8757 26979 8815 26985
rect 8757 26945 8769 26979
rect 8803 26976 8815 26979
rect 9766 26976 9772 26988
rect 8803 26948 9772 26976
rect 8803 26945 8815 26948
rect 8757 26939 8815 26945
rect 9766 26936 9772 26948
rect 9824 26936 9830 26988
rect 9950 26976 9956 26988
rect 9911 26948 9956 26976
rect 9950 26936 9956 26948
rect 10008 26936 10014 26988
rect 12250 26976 12256 26988
rect 12211 26948 12256 26976
rect 12250 26936 12256 26948
rect 12308 26936 12314 26988
rect 13081 26979 13139 26985
rect 13081 26945 13093 26979
rect 13127 26976 13139 26979
rect 14274 26976 14280 26988
rect 13127 26948 14280 26976
rect 13127 26945 13139 26948
rect 13081 26939 13139 26945
rect 14274 26936 14280 26948
rect 14332 26936 14338 26988
rect 17313 26979 17371 26985
rect 17313 26945 17325 26979
rect 17359 26976 17371 26979
rect 58342 26976 58348 26988
rect 17359 26948 18276 26976
rect 58303 26948 58348 26976
rect 17359 26945 17371 26948
rect 17313 26939 17371 26945
rect 2225 26911 2283 26917
rect 2225 26877 2237 26911
rect 2271 26877 2283 26911
rect 2225 26871 2283 26877
rect 2409 26911 2467 26917
rect 2409 26877 2421 26911
rect 2455 26908 2467 26911
rect 2682 26908 2688 26920
rect 2455 26880 2688 26908
rect 2455 26877 2467 26880
rect 2409 26871 2467 26877
rect 2682 26868 2688 26880
rect 2740 26868 2746 26920
rect 5350 26908 5356 26920
rect 5311 26880 5356 26908
rect 5350 26868 5356 26880
rect 5408 26868 5414 26920
rect 7650 26868 7656 26920
rect 7708 26908 7714 26920
rect 12158 26908 12164 26920
rect 7708 26880 12164 26908
rect 7708 26868 7714 26880
rect 12158 26868 12164 26880
rect 12216 26908 12222 26920
rect 12986 26908 12992 26920
rect 12216 26880 12992 26908
rect 12216 26868 12222 26880
rect 12986 26868 12992 26880
rect 13044 26908 13050 26920
rect 13725 26911 13783 26917
rect 13725 26908 13737 26911
rect 13044 26880 13737 26908
rect 13044 26868 13050 26880
rect 13725 26877 13737 26880
rect 13771 26877 13783 26911
rect 13725 26871 13783 26877
rect 16206 26868 16212 26920
rect 16264 26908 16270 26920
rect 16301 26911 16359 26917
rect 16301 26908 16313 26911
rect 16264 26880 16313 26908
rect 16264 26868 16270 26880
rect 16301 26877 16313 26880
rect 16347 26908 16359 26911
rect 17405 26911 17463 26917
rect 17405 26908 17417 26911
rect 16347 26880 17417 26908
rect 16347 26877 16359 26880
rect 16301 26871 16359 26877
rect 17405 26877 17417 26880
rect 17451 26877 17463 26911
rect 17405 26871 17463 26877
rect 17589 26911 17647 26917
rect 17589 26877 17601 26911
rect 17635 26908 17647 26911
rect 18046 26908 18052 26920
rect 17635 26880 18052 26908
rect 17635 26877 17647 26880
rect 17589 26871 17647 26877
rect 18046 26868 18052 26880
rect 18104 26868 18110 26920
rect 12437 26843 12495 26849
rect 12437 26809 12449 26843
rect 12483 26840 12495 26843
rect 13354 26840 13360 26852
rect 12483 26812 13360 26840
rect 12483 26809 12495 26812
rect 12437 26803 12495 26809
rect 13354 26800 13360 26812
rect 13412 26800 13418 26852
rect 2866 26772 2872 26784
rect 2827 26744 2872 26772
rect 2866 26732 2872 26744
rect 2924 26732 2930 26784
rect 3326 26732 3332 26784
rect 3384 26772 3390 26784
rect 3605 26775 3663 26781
rect 3605 26772 3617 26775
rect 3384 26744 3617 26772
rect 3384 26732 3390 26744
rect 3605 26741 3617 26744
rect 3651 26741 3663 26775
rect 3605 26735 3663 26741
rect 4341 26775 4399 26781
rect 4341 26741 4353 26775
rect 4387 26772 4399 26775
rect 4706 26772 4712 26784
rect 4387 26744 4712 26772
rect 4387 26741 4399 26744
rect 4341 26735 4399 26741
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 5994 26772 6000 26784
rect 5955 26744 6000 26772
rect 5994 26732 6000 26744
rect 6052 26732 6058 26784
rect 8941 26775 8999 26781
rect 8941 26741 8953 26775
rect 8987 26772 8999 26775
rect 9122 26772 9128 26784
rect 8987 26744 9128 26772
rect 8987 26741 8999 26744
rect 8941 26735 8999 26741
rect 9122 26732 9128 26744
rect 9180 26732 9186 26784
rect 10137 26775 10195 26781
rect 10137 26741 10149 26775
rect 10183 26772 10195 26775
rect 10686 26772 10692 26784
rect 10183 26744 10692 26772
rect 10183 26741 10195 26744
rect 10137 26735 10195 26741
rect 10686 26732 10692 26744
rect 10744 26732 10750 26784
rect 12897 26775 12955 26781
rect 12897 26741 12909 26775
rect 12943 26772 12955 26775
rect 13446 26772 13452 26784
rect 12943 26744 13452 26772
rect 12943 26741 12955 26744
rect 12897 26735 12955 26741
rect 13446 26732 13452 26744
rect 13504 26732 13510 26784
rect 16945 26775 17003 26781
rect 16945 26741 16957 26775
rect 16991 26772 17003 26775
rect 17034 26772 17040 26784
rect 16991 26744 17040 26772
rect 16991 26741 17003 26744
rect 16945 26735 17003 26741
rect 17034 26732 17040 26744
rect 17092 26732 17098 26784
rect 18248 26781 18276 26948
rect 58342 26936 58348 26948
rect 58400 26936 58406 26988
rect 18233 26775 18291 26781
rect 18233 26741 18245 26775
rect 18279 26772 18291 26775
rect 18506 26772 18512 26784
rect 18279 26744 18512 26772
rect 18279 26741 18291 26744
rect 18233 26735 18291 26741
rect 18506 26732 18512 26744
rect 18564 26732 18570 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 2130 26528 2136 26580
rect 2188 26568 2194 26580
rect 8386 26568 8392 26580
rect 2188 26540 8392 26568
rect 2188 26528 2194 26540
rect 4525 26503 4583 26509
rect 4525 26500 4537 26503
rect 2516 26472 4537 26500
rect 2516 26444 2544 26472
rect 4525 26469 4537 26472
rect 4571 26500 4583 26503
rect 5626 26500 5632 26512
rect 4571 26472 5632 26500
rect 4571 26469 4583 26472
rect 4525 26463 4583 26469
rect 5626 26460 5632 26472
rect 5684 26460 5690 26512
rect 2314 26432 2320 26444
rect 2275 26404 2320 26432
rect 2314 26392 2320 26404
rect 2372 26392 2378 26444
rect 2498 26432 2504 26444
rect 2459 26404 2504 26432
rect 2498 26392 2504 26404
rect 2556 26392 2562 26444
rect 2774 26392 2780 26444
rect 2832 26432 2838 26444
rect 5350 26432 5356 26444
rect 2832 26404 5356 26432
rect 2832 26392 2838 26404
rect 5350 26392 5356 26404
rect 5408 26432 5414 26444
rect 5736 26441 5764 26540
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 10413 26571 10471 26577
rect 10413 26537 10425 26571
rect 10459 26568 10471 26571
rect 12342 26568 12348 26580
rect 10459 26540 12348 26568
rect 10459 26537 10471 26540
rect 10413 26531 10471 26537
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 57149 26571 57207 26577
rect 57149 26537 57161 26571
rect 57195 26568 57207 26571
rect 58342 26568 58348 26580
rect 57195 26540 58348 26568
rect 57195 26537 57207 26540
rect 57149 26531 57207 26537
rect 58342 26528 58348 26540
rect 58400 26528 58406 26580
rect 6181 26503 6239 26509
rect 6181 26469 6193 26503
rect 6227 26469 6239 26503
rect 6181 26463 6239 26469
rect 5537 26435 5595 26441
rect 5537 26432 5549 26435
rect 5408 26404 5549 26432
rect 5408 26392 5414 26404
rect 5537 26401 5549 26404
rect 5583 26401 5595 26435
rect 5537 26395 5595 26401
rect 5721 26435 5779 26441
rect 5721 26401 5733 26435
rect 5767 26401 5779 26435
rect 5721 26395 5779 26401
rect 2682 26324 2688 26376
rect 2740 26364 2746 26376
rect 4065 26367 4123 26373
rect 4065 26364 4077 26367
rect 2740 26336 4077 26364
rect 2740 26324 2746 26336
rect 4065 26333 4077 26336
rect 4111 26364 4123 26367
rect 6196 26364 6224 26463
rect 6362 26460 6368 26512
rect 6420 26500 6426 26512
rect 7650 26500 7656 26512
rect 6420 26472 7656 26500
rect 6420 26460 6426 26472
rect 7650 26460 7656 26472
rect 7708 26460 7714 26512
rect 11057 26503 11115 26509
rect 11057 26469 11069 26503
rect 11103 26500 11115 26503
rect 11422 26500 11428 26512
rect 11103 26472 11428 26500
rect 11103 26469 11115 26472
rect 11057 26463 11115 26469
rect 11422 26460 11428 26472
rect 11480 26460 11486 26512
rect 17037 26503 17095 26509
rect 17037 26500 17049 26503
rect 16546 26472 17049 26500
rect 9861 26435 9919 26441
rect 9861 26401 9873 26435
rect 9907 26432 9919 26435
rect 10410 26432 10416 26444
rect 9907 26404 10416 26432
rect 9907 26401 9919 26404
rect 9861 26395 9919 26401
rect 10410 26392 10416 26404
rect 10468 26392 10474 26444
rect 7009 26367 7067 26373
rect 7009 26364 7021 26367
rect 4111 26336 5580 26364
rect 6196 26336 7021 26364
rect 4111 26333 4123 26336
rect 4065 26327 4123 26333
rect 5552 26308 5580 26336
rect 7009 26333 7021 26336
rect 7055 26333 7067 26367
rect 10870 26364 10876 26376
rect 7009 26327 7067 26333
rect 7208 26336 9812 26364
rect 10831 26336 10876 26364
rect 5534 26256 5540 26308
rect 5592 26256 5598 26308
rect 5813 26299 5871 26305
rect 5813 26265 5825 26299
rect 5859 26296 5871 26299
rect 6362 26296 6368 26308
rect 5859 26268 6368 26296
rect 5859 26265 5871 26268
rect 5813 26259 5871 26265
rect 6362 26256 6368 26268
rect 6420 26256 6426 26308
rect 2593 26231 2651 26237
rect 2593 26197 2605 26231
rect 2639 26228 2651 26231
rect 2682 26228 2688 26240
rect 2639 26200 2688 26228
rect 2639 26197 2651 26200
rect 2593 26191 2651 26197
rect 2682 26188 2688 26200
rect 2740 26188 2746 26240
rect 2958 26188 2964 26240
rect 3016 26228 3022 26240
rect 7208 26237 7236 26336
rect 9784 26308 9812 26336
rect 10870 26324 10876 26336
rect 10928 26324 10934 26376
rect 16393 26367 16451 26373
rect 16393 26333 16405 26367
rect 16439 26364 16451 26367
rect 16546 26364 16574 26472
rect 17037 26469 17049 26472
rect 17083 26469 17095 26503
rect 17037 26463 17095 26469
rect 43714 26460 43720 26512
rect 43772 26500 43778 26512
rect 44085 26503 44143 26509
rect 44085 26500 44097 26503
rect 43772 26472 44097 26500
rect 43772 26460 43778 26472
rect 44085 26469 44097 26472
rect 44131 26469 44143 26503
rect 57606 26500 57612 26512
rect 57567 26472 57612 26500
rect 44085 26463 44143 26469
rect 57606 26460 57612 26472
rect 57664 26460 57670 26512
rect 58066 26460 58072 26512
rect 58124 26500 58130 26512
rect 58161 26503 58219 26509
rect 58161 26500 58173 26503
rect 58124 26472 58173 26500
rect 58124 26460 58130 26472
rect 58161 26469 58173 26472
rect 58207 26469 58219 26503
rect 58161 26463 58219 26469
rect 17681 26435 17739 26441
rect 17681 26401 17693 26435
rect 17727 26432 17739 26435
rect 18230 26432 18236 26444
rect 17727 26404 18236 26432
rect 17727 26401 17739 26404
rect 17681 26395 17739 26401
rect 18230 26392 18236 26404
rect 18288 26392 18294 26444
rect 16439 26336 16574 26364
rect 17405 26367 17463 26373
rect 16439 26333 16451 26336
rect 16393 26327 16451 26333
rect 17405 26333 17417 26367
rect 17451 26364 17463 26367
rect 18506 26364 18512 26376
rect 17451 26336 18512 26364
rect 17451 26333 17463 26336
rect 17405 26327 17463 26333
rect 18506 26324 18512 26336
rect 18564 26324 18570 26376
rect 44269 26367 44327 26373
rect 44269 26333 44281 26367
rect 44315 26364 44327 26367
rect 56502 26364 56508 26376
rect 44315 26336 56508 26364
rect 44315 26333 44327 26336
rect 44269 26327 44327 26333
rect 56502 26324 56508 26336
rect 56560 26324 56566 26376
rect 57514 26324 57520 26376
rect 57572 26364 57578 26376
rect 58342 26364 58348 26376
rect 57572 26336 58348 26364
rect 57572 26324 57578 26336
rect 58342 26324 58348 26336
rect 58400 26324 58406 26376
rect 7745 26299 7803 26305
rect 7745 26265 7757 26299
rect 7791 26296 7803 26299
rect 8386 26296 8392 26308
rect 7791 26268 8392 26296
rect 7791 26265 7803 26268
rect 7745 26259 7803 26265
rect 8386 26256 8392 26268
rect 8444 26256 8450 26308
rect 9766 26256 9772 26308
rect 9824 26256 9830 26308
rect 9950 26296 9956 26308
rect 9911 26268 9956 26296
rect 9950 26256 9956 26268
rect 10008 26256 10014 26308
rect 10045 26299 10103 26305
rect 10045 26265 10057 26299
rect 10091 26296 10103 26299
rect 11146 26296 11152 26308
rect 10091 26268 11152 26296
rect 10091 26265 10103 26268
rect 10045 26259 10103 26265
rect 11146 26256 11152 26268
rect 11204 26296 11210 26308
rect 11609 26299 11667 26305
rect 11609 26296 11621 26299
rect 11204 26268 11621 26296
rect 11204 26256 11210 26268
rect 11609 26265 11621 26268
rect 11655 26296 11667 26299
rect 12158 26296 12164 26308
rect 11655 26268 12164 26296
rect 11655 26265 11667 26268
rect 11609 26259 11667 26265
rect 12158 26256 12164 26268
rect 12216 26256 12222 26308
rect 17497 26299 17555 26305
rect 17497 26265 17509 26299
rect 17543 26296 17555 26299
rect 17954 26296 17960 26308
rect 17543 26268 17960 26296
rect 17543 26265 17555 26268
rect 17497 26259 17555 26265
rect 17954 26256 17960 26268
rect 18012 26296 18018 26308
rect 18233 26299 18291 26305
rect 18233 26296 18245 26299
rect 18012 26268 18245 26296
rect 18012 26256 18018 26268
rect 18233 26265 18245 26268
rect 18279 26265 18291 26299
rect 18233 26259 18291 26265
rect 7193 26231 7251 26237
rect 3016 26200 3061 26228
rect 3016 26188 3022 26200
rect 7193 26197 7205 26231
rect 7239 26228 7251 26231
rect 7239 26200 7273 26228
rect 7239 26197 7251 26200
rect 7193 26191 7251 26197
rect 16574 26188 16580 26240
rect 16632 26228 16638 26240
rect 16632 26200 16677 26228
rect 16632 26188 16638 26200
rect 18506 26188 18512 26240
rect 18564 26228 18570 26240
rect 18785 26231 18843 26237
rect 18785 26228 18797 26231
rect 18564 26200 18797 26228
rect 18564 26188 18570 26200
rect 18785 26197 18797 26200
rect 18831 26197 18843 26231
rect 18785 26191 18843 26197
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1670 26024 1676 26036
rect 1631 25996 1676 26024
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 2130 25984 2136 26036
rect 2188 26024 2194 26036
rect 2314 26024 2320 26036
rect 2188 25996 2320 26024
rect 2188 25984 2194 25996
rect 2314 25984 2320 25996
rect 2372 25984 2378 26036
rect 2682 25984 2688 26036
rect 2740 26024 2746 26036
rect 3234 26024 3240 26036
rect 2740 25996 3240 26024
rect 2740 25984 2746 25996
rect 3234 25984 3240 25996
rect 3292 25984 3298 26036
rect 3326 25984 3332 26036
rect 3384 26024 3390 26036
rect 3513 26027 3571 26033
rect 3513 26024 3525 26027
rect 3384 25996 3525 26024
rect 3384 25984 3390 25996
rect 3513 25993 3525 25996
rect 3559 25993 3571 26027
rect 3513 25987 3571 25993
rect 5350 25984 5356 26036
rect 5408 26024 5414 26036
rect 5905 26027 5963 26033
rect 5905 26024 5917 26027
rect 5408 25996 5917 26024
rect 5408 25984 5414 25996
rect 5905 25993 5917 25996
rect 5951 25993 5963 26027
rect 57514 26024 57520 26036
rect 57475 25996 57520 26024
rect 5905 25987 5963 25993
rect 57514 25984 57520 25996
rect 57572 25984 57578 26036
rect 18506 25916 18512 25968
rect 18564 25956 18570 25968
rect 19337 25959 19395 25965
rect 19337 25956 19349 25959
rect 18564 25928 19349 25956
rect 18564 25916 18570 25928
rect 19337 25925 19349 25928
rect 19383 25925 19395 25959
rect 19337 25919 19395 25925
rect 1857 25891 1915 25897
rect 1857 25857 1869 25891
rect 1903 25888 1915 25891
rect 2038 25888 2044 25900
rect 1903 25860 2044 25888
rect 1903 25857 1915 25860
rect 1857 25851 1915 25857
rect 2038 25848 2044 25860
rect 2096 25848 2102 25900
rect 2866 25888 2872 25900
rect 2827 25860 2872 25888
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 5994 25848 6000 25900
rect 6052 25888 6058 25900
rect 6549 25891 6607 25897
rect 6549 25888 6561 25891
rect 6052 25860 6561 25888
rect 6052 25848 6058 25860
rect 6549 25857 6561 25860
rect 6595 25857 6607 25891
rect 6549 25851 6607 25857
rect 12342 25848 12348 25900
rect 12400 25888 12406 25900
rect 12713 25891 12771 25897
rect 12713 25888 12725 25891
rect 12400 25860 12725 25888
rect 12400 25848 12406 25860
rect 12713 25857 12725 25860
rect 12759 25857 12771 25891
rect 17034 25888 17040 25900
rect 16995 25860 17040 25888
rect 12713 25851 12771 25857
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 18322 25848 18328 25900
rect 18380 25888 18386 25900
rect 19245 25891 19303 25897
rect 19245 25888 19257 25891
rect 18380 25860 19257 25888
rect 18380 25848 18386 25860
rect 19245 25857 19257 25860
rect 19291 25857 19303 25891
rect 19245 25851 19303 25857
rect 56965 25891 57023 25897
rect 56965 25857 56977 25891
rect 57011 25888 57023 25891
rect 58342 25888 58348 25900
rect 57011 25860 58348 25888
rect 57011 25857 57023 25860
rect 56965 25851 57023 25857
rect 58342 25848 58348 25860
rect 58400 25848 58406 25900
rect 19153 25823 19211 25829
rect 19153 25789 19165 25823
rect 19199 25820 19211 25823
rect 19426 25820 19432 25832
rect 19199 25792 19432 25820
rect 19199 25789 19211 25792
rect 19153 25783 19211 25789
rect 19426 25780 19432 25792
rect 19484 25820 19490 25832
rect 19484 25792 20300 25820
rect 19484 25780 19490 25792
rect 6362 25712 6368 25764
rect 6420 25752 6426 25764
rect 7193 25755 7251 25761
rect 7193 25752 7205 25755
rect 6420 25724 7205 25752
rect 6420 25712 6426 25724
rect 7193 25721 7205 25724
rect 7239 25721 7251 25755
rect 7193 25715 7251 25721
rect 9214 25712 9220 25764
rect 9272 25752 9278 25764
rect 14090 25752 14096 25764
rect 9272 25724 14096 25752
rect 9272 25712 9278 25724
rect 14090 25712 14096 25724
rect 14148 25712 14154 25764
rect 3050 25684 3056 25696
rect 3011 25656 3056 25684
rect 3050 25644 3056 25656
rect 3108 25644 3114 25696
rect 3234 25644 3240 25696
rect 3292 25684 3298 25696
rect 4157 25687 4215 25693
rect 4157 25684 4169 25687
rect 3292 25656 4169 25684
rect 3292 25644 3298 25656
rect 4157 25653 4169 25656
rect 4203 25684 4215 25687
rect 4798 25684 4804 25696
rect 4203 25656 4804 25684
rect 4203 25653 4215 25656
rect 4157 25647 4215 25653
rect 4798 25644 4804 25656
rect 4856 25644 4862 25696
rect 6733 25687 6791 25693
rect 6733 25653 6745 25687
rect 6779 25684 6791 25687
rect 6822 25684 6828 25696
rect 6779 25656 6828 25684
rect 6779 25653 6791 25656
rect 6733 25647 6791 25653
rect 6822 25644 6828 25656
rect 6880 25644 6886 25696
rect 10410 25644 10416 25696
rect 10468 25684 10474 25696
rect 10505 25687 10563 25693
rect 10505 25684 10517 25687
rect 10468 25656 10517 25684
rect 10468 25644 10474 25656
rect 10505 25653 10517 25656
rect 10551 25653 10563 25687
rect 10505 25647 10563 25653
rect 12897 25687 12955 25693
rect 12897 25653 12909 25687
rect 12943 25684 12955 25687
rect 14182 25684 14188 25696
rect 12943 25656 14188 25684
rect 12943 25653 12955 25656
rect 12897 25647 12955 25653
rect 14182 25644 14188 25656
rect 14240 25644 14246 25696
rect 16850 25684 16856 25696
rect 16811 25656 16856 25684
rect 16850 25644 16856 25656
rect 16908 25644 16914 25696
rect 17957 25687 18015 25693
rect 17957 25653 17969 25687
rect 18003 25684 18015 25687
rect 18230 25684 18236 25696
rect 18003 25656 18236 25684
rect 18003 25653 18015 25656
rect 17957 25647 18015 25653
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 18506 25684 18512 25696
rect 18467 25656 18512 25684
rect 18506 25644 18512 25656
rect 18564 25644 18570 25696
rect 19610 25644 19616 25696
rect 19668 25684 19674 25696
rect 20272 25693 20300 25792
rect 55858 25712 55864 25764
rect 55916 25752 55922 25764
rect 58161 25755 58219 25761
rect 58161 25752 58173 25755
rect 55916 25724 58173 25752
rect 55916 25712 55922 25724
rect 58161 25721 58173 25724
rect 58207 25721 58219 25755
rect 58161 25715 58219 25721
rect 19705 25687 19763 25693
rect 19705 25684 19717 25687
rect 19668 25656 19717 25684
rect 19668 25644 19674 25656
rect 19705 25653 19717 25656
rect 19751 25653 19763 25687
rect 19705 25647 19763 25653
rect 20257 25687 20315 25693
rect 20257 25653 20269 25687
rect 20303 25684 20315 25687
rect 20346 25684 20352 25696
rect 20303 25656 20352 25684
rect 20303 25653 20315 25656
rect 20257 25647 20315 25653
rect 20346 25644 20352 25656
rect 20404 25644 20410 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1670 25480 1676 25492
rect 1631 25452 1676 25480
rect 1670 25440 1676 25452
rect 1728 25440 1734 25492
rect 3145 25483 3203 25489
rect 3145 25449 3157 25483
rect 3191 25480 3203 25483
rect 8294 25480 8300 25492
rect 3191 25452 8300 25480
rect 3191 25449 3203 25452
rect 3145 25443 3203 25449
rect 8294 25440 8300 25452
rect 8352 25440 8358 25492
rect 9674 25440 9680 25492
rect 9732 25480 9738 25492
rect 10873 25483 10931 25489
rect 10873 25480 10885 25483
rect 9732 25452 10885 25480
rect 9732 25440 9738 25452
rect 10873 25449 10885 25452
rect 10919 25449 10931 25483
rect 10873 25443 10931 25449
rect 57422 25440 57428 25492
rect 57480 25480 57486 25492
rect 58802 25480 58808 25492
rect 57480 25452 58808 25480
rect 57480 25440 57486 25452
rect 58802 25440 58808 25452
rect 58860 25440 58866 25492
rect 2590 25372 2596 25424
rect 2648 25412 2654 25424
rect 5905 25415 5963 25421
rect 5905 25412 5917 25415
rect 2648 25384 5917 25412
rect 2648 25372 2654 25384
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25276 1915 25279
rect 2406 25276 2412 25288
rect 1903 25248 2412 25276
rect 1903 25245 1915 25248
rect 1857 25239 1915 25245
rect 2406 25236 2412 25248
rect 2464 25236 2470 25288
rect 2958 25276 2964 25288
rect 2919 25248 2964 25276
rect 2958 25236 2964 25248
rect 3016 25236 3022 25288
rect 5644 25276 5672 25384
rect 5905 25381 5917 25384
rect 5951 25381 5963 25415
rect 57790 25412 57796 25424
rect 5905 25375 5963 25381
rect 57624 25384 57796 25412
rect 5718 25304 5724 25356
rect 5776 25344 5782 25356
rect 7653 25347 7711 25353
rect 7653 25344 7665 25347
rect 5776 25316 7665 25344
rect 5776 25304 5782 25316
rect 7653 25313 7665 25316
rect 7699 25313 7711 25347
rect 16850 25344 16856 25356
rect 7653 25307 7711 25313
rect 11072 25316 16856 25344
rect 5644 25248 6132 25276
rect 2038 25168 2044 25220
rect 2096 25208 2102 25220
rect 2317 25211 2375 25217
rect 2317 25208 2329 25211
rect 2096 25180 2329 25208
rect 2096 25168 2102 25180
rect 2317 25177 2329 25180
rect 2363 25208 2375 25211
rect 5994 25208 6000 25220
rect 2363 25180 6000 25208
rect 2363 25177 2375 25180
rect 2317 25171 2375 25177
rect 5994 25168 6000 25180
rect 6052 25168 6058 25220
rect 6104 25140 6132 25248
rect 6914 25168 6920 25220
rect 6972 25168 6978 25220
rect 7377 25211 7435 25217
rect 7377 25177 7389 25211
rect 7423 25208 7435 25211
rect 11072 25208 11100 25316
rect 16850 25304 16856 25316
rect 16908 25304 16914 25356
rect 57308 25347 57366 25353
rect 57308 25313 57320 25347
rect 57354 25344 57366 25347
rect 57624 25344 57652 25384
rect 57790 25372 57796 25384
rect 57848 25372 57854 25424
rect 57354 25316 57652 25344
rect 57354 25313 57366 25316
rect 57308 25307 57366 25313
rect 57698 25304 57704 25356
rect 57756 25344 57762 25356
rect 58345 25347 58403 25353
rect 57756 25316 57801 25344
rect 57756 25304 57762 25316
rect 58345 25313 58357 25347
rect 58391 25344 58403 25347
rect 58526 25344 58532 25356
rect 58391 25316 58532 25344
rect 58391 25313 58403 25316
rect 58345 25307 58403 25313
rect 58526 25304 58532 25316
rect 58584 25304 58590 25356
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25276 12679 25279
rect 15378 25276 15384 25288
rect 12667 25248 15384 25276
rect 12667 25245 12679 25248
rect 12621 25239 12679 25245
rect 15378 25236 15384 25248
rect 15436 25236 15442 25288
rect 19610 25276 19616 25288
rect 19571 25248 19616 25276
rect 19610 25236 19616 25248
rect 19668 25236 19674 25288
rect 57146 25236 57152 25288
rect 57204 25276 57210 25288
rect 57422 25276 57428 25288
rect 57204 25248 57249 25276
rect 57383 25248 57428 25276
rect 57204 25236 57210 25248
rect 57422 25236 57428 25248
rect 57480 25236 57486 25288
rect 58158 25276 58164 25288
rect 58119 25248 58164 25276
rect 58158 25236 58164 25248
rect 58216 25236 58222 25288
rect 7423 25180 11100 25208
rect 7423 25177 7435 25180
rect 7377 25171 7435 25177
rect 11790 25168 11796 25220
rect 11848 25168 11854 25220
rect 12066 25168 12072 25220
rect 12124 25208 12130 25220
rect 12345 25211 12403 25217
rect 12345 25208 12357 25211
rect 12124 25180 12357 25208
rect 12124 25168 12130 25180
rect 12345 25177 12357 25180
rect 12391 25177 12403 25211
rect 12345 25171 12403 25177
rect 16206 25140 16212 25152
rect 6104 25112 16212 25140
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 18322 25100 18328 25152
rect 18380 25140 18386 25152
rect 18601 25143 18659 25149
rect 18601 25140 18613 25143
rect 18380 25112 18613 25140
rect 18380 25100 18386 25112
rect 18601 25109 18613 25112
rect 18647 25109 18659 25143
rect 18601 25103 18659 25109
rect 18690 25100 18696 25152
rect 18748 25140 18754 25152
rect 19429 25143 19487 25149
rect 19429 25140 19441 25143
rect 18748 25112 19441 25140
rect 18748 25100 18754 25112
rect 19429 25109 19441 25112
rect 19475 25109 19487 25143
rect 56502 25140 56508 25152
rect 56463 25112 56508 25140
rect 19429 25103 19487 25109
rect 56502 25100 56508 25112
rect 56560 25100 56566 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 4982 24828 4988 24880
rect 5040 24828 5046 24880
rect 14826 24868 14832 24880
rect 14674 24840 14832 24868
rect 14826 24828 14832 24840
rect 14884 24828 14890 24880
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 2961 24803 3019 24809
rect 2961 24800 2973 24803
rect 1903 24772 2973 24800
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 2961 24769 2973 24772
rect 3007 24800 3019 24803
rect 3694 24800 3700 24812
rect 3007 24772 3700 24800
rect 3007 24769 3019 24772
rect 2961 24763 3019 24769
rect 3694 24760 3700 24772
rect 3752 24760 3758 24812
rect 5718 24760 5724 24812
rect 5776 24800 5782 24812
rect 5776 24772 5821 24800
rect 5776 24760 5782 24772
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 8202 24800 8208 24812
rect 6972 24772 8208 24800
rect 6972 24760 6978 24772
rect 8202 24760 8208 24772
rect 8260 24800 8266 24812
rect 8260 24772 8694 24800
rect 8260 24760 8266 24772
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 19153 24803 19211 24809
rect 15436 24772 15481 24800
rect 15436 24760 15442 24772
rect 19153 24769 19165 24803
rect 19199 24800 19211 24803
rect 19610 24800 19616 24812
rect 19199 24772 19616 24800
rect 19199 24769 19211 24772
rect 19153 24763 19211 24769
rect 19610 24760 19616 24772
rect 19668 24760 19674 24812
rect 58342 24800 58348 24812
rect 58303 24772 58348 24800
rect 58342 24760 58348 24772
rect 58400 24760 58406 24812
rect 2498 24692 2504 24744
rect 2556 24732 2562 24744
rect 5445 24735 5503 24741
rect 5445 24732 5457 24735
rect 2556 24704 5457 24732
rect 2556 24692 2562 24704
rect 5445 24701 5457 24704
rect 5491 24701 5503 24735
rect 5445 24695 5503 24701
rect 8297 24735 8355 24741
rect 8297 24701 8309 24735
rect 8343 24732 8355 24735
rect 8386 24732 8392 24744
rect 8343 24704 8392 24732
rect 8343 24701 8355 24704
rect 8297 24695 8355 24701
rect 8386 24692 8392 24704
rect 8444 24692 8450 24744
rect 9766 24732 9772 24744
rect 9727 24704 9772 24732
rect 9766 24692 9772 24704
rect 9824 24692 9830 24744
rect 10042 24732 10048 24744
rect 10003 24704 10048 24732
rect 10042 24692 10048 24704
rect 10100 24692 10106 24744
rect 15105 24735 15163 24741
rect 15105 24701 15117 24735
rect 15151 24732 15163 24735
rect 18690 24732 18696 24744
rect 15151 24704 18696 24732
rect 15151 24701 15163 24704
rect 15105 24695 15163 24701
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 1670 24664 1676 24676
rect 1631 24636 1676 24664
rect 1670 24624 1676 24636
rect 1728 24624 1734 24676
rect 1854 24624 1860 24676
rect 1912 24664 1918 24676
rect 3973 24667 4031 24673
rect 3973 24664 3985 24667
rect 1912 24636 3985 24664
rect 1912 24624 1918 24636
rect 3973 24633 3985 24636
rect 4019 24633 4031 24667
rect 3973 24627 4031 24633
rect 17218 24624 17224 24676
rect 17276 24664 17282 24676
rect 18969 24667 19027 24673
rect 18969 24664 18981 24667
rect 17276 24636 18981 24664
rect 17276 24624 17282 24636
rect 18969 24633 18981 24636
rect 19015 24633 19027 24667
rect 18969 24627 19027 24633
rect 58066 24624 58072 24676
rect 58124 24664 58130 24676
rect 58161 24667 58219 24673
rect 58161 24664 58173 24667
rect 58124 24636 58173 24664
rect 58124 24624 58130 24636
rect 58161 24633 58173 24636
rect 58207 24633 58219 24667
rect 58161 24627 58219 24633
rect 2406 24596 2412 24608
rect 2367 24568 2412 24596
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 3510 24596 3516 24608
rect 3471 24568 3516 24596
rect 3510 24556 3516 24568
rect 3568 24556 3574 24608
rect 4062 24556 4068 24608
rect 4120 24596 4126 24608
rect 9214 24596 9220 24608
rect 4120 24568 9220 24596
rect 4120 24556 4126 24568
rect 9214 24556 9220 24568
rect 9272 24556 9278 24608
rect 13630 24596 13636 24608
rect 13543 24568 13636 24596
rect 13630 24556 13636 24568
rect 13688 24596 13694 24608
rect 18322 24596 18328 24608
rect 13688 24568 18328 24596
rect 13688 24556 13694 24568
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 18509 24599 18567 24605
rect 18509 24565 18521 24599
rect 18555 24596 18567 24599
rect 18782 24596 18788 24608
rect 18555 24568 18788 24596
rect 18555 24565 18567 24568
rect 18509 24559 18567 24565
rect 18782 24556 18788 24568
rect 18840 24556 18846 24608
rect 19334 24556 19340 24608
rect 19392 24596 19398 24608
rect 19613 24599 19671 24605
rect 19613 24596 19625 24599
rect 19392 24568 19625 24596
rect 19392 24556 19398 24568
rect 19613 24565 19625 24568
rect 19659 24565 19671 24599
rect 19613 24559 19671 24565
rect 56965 24599 57023 24605
rect 56965 24565 56977 24599
rect 57011 24596 57023 24599
rect 57146 24596 57152 24608
rect 57011 24568 57152 24596
rect 57011 24565 57023 24568
rect 56965 24559 57023 24565
rect 57146 24556 57152 24568
rect 57204 24556 57210 24608
rect 57238 24556 57244 24608
rect 57296 24596 57302 24608
rect 57425 24599 57483 24605
rect 57425 24596 57437 24599
rect 57296 24568 57437 24596
rect 57296 24556 57302 24568
rect 57425 24565 57437 24568
rect 57471 24596 57483 24599
rect 57698 24596 57704 24608
rect 57471 24568 57704 24596
rect 57471 24565 57483 24568
rect 57425 24559 57483 24565
rect 57698 24556 57704 24568
rect 57756 24556 57762 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 3510 24352 3516 24404
rect 3568 24392 3574 24404
rect 3568 24364 11928 24392
rect 3568 24352 3574 24364
rect 2774 24256 2780 24268
rect 2735 24228 2780 24256
rect 2774 24216 2780 24228
rect 2832 24216 2838 24268
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24256 3019 24259
rect 3418 24256 3424 24268
rect 3007 24228 3424 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 3418 24216 3424 24228
rect 3476 24216 3482 24268
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24188 1915 24191
rect 3528 24188 3556 24352
rect 3694 24284 3700 24336
rect 3752 24324 3758 24336
rect 6086 24324 6092 24336
rect 3752 24296 6092 24324
rect 3752 24284 3758 24296
rect 6086 24284 6092 24296
rect 6144 24284 6150 24336
rect 11900 24324 11928 24364
rect 11974 24352 11980 24404
rect 12032 24392 12038 24404
rect 12161 24395 12219 24401
rect 12161 24392 12173 24395
rect 12032 24364 12173 24392
rect 12032 24352 12038 24364
rect 12161 24361 12173 24364
rect 12207 24361 12219 24395
rect 12161 24355 12219 24361
rect 18046 24352 18052 24404
rect 18104 24392 18110 24404
rect 18509 24395 18567 24401
rect 18509 24392 18521 24395
rect 18104 24364 18521 24392
rect 18104 24352 18110 24364
rect 18509 24361 18521 24364
rect 18555 24361 18567 24395
rect 19610 24392 19616 24404
rect 19571 24364 19616 24392
rect 18509 24355 18567 24361
rect 19610 24352 19616 24364
rect 19668 24352 19674 24404
rect 57701 24395 57759 24401
rect 57701 24361 57713 24395
rect 57747 24392 57759 24395
rect 58342 24392 58348 24404
rect 57747 24364 58348 24392
rect 57747 24361 57759 24364
rect 57701 24355 57759 24361
rect 58342 24352 58348 24364
rect 58400 24352 58406 24404
rect 14918 24324 14924 24336
rect 11900 24296 14924 24324
rect 14918 24284 14924 24296
rect 14976 24284 14982 24336
rect 57054 24284 57060 24336
rect 57112 24324 57118 24336
rect 58161 24327 58219 24333
rect 58161 24324 58173 24327
rect 57112 24296 58173 24324
rect 57112 24284 57118 24296
rect 58161 24293 58173 24296
rect 58207 24293 58219 24327
rect 58161 24287 58219 24293
rect 10042 24216 10048 24268
rect 10100 24256 10106 24268
rect 10413 24259 10471 24265
rect 10413 24256 10425 24259
rect 10100 24228 10425 24256
rect 10100 24216 10106 24228
rect 10413 24225 10425 24228
rect 10459 24225 10471 24259
rect 10686 24256 10692 24268
rect 10647 24228 10692 24256
rect 10413 24219 10471 24225
rect 10686 24216 10692 24228
rect 10744 24216 10750 24268
rect 20254 24256 20260 24268
rect 20215 24228 20260 24256
rect 20254 24216 20260 24228
rect 20312 24216 20318 24268
rect 1903 24160 3556 24188
rect 1903 24157 1915 24160
rect 1857 24151 1915 24157
rect 11790 24148 11796 24200
rect 11848 24188 11854 24200
rect 13906 24188 13912 24200
rect 11848 24160 13912 24188
rect 11848 24148 11854 24160
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 18782 24188 18788 24200
rect 18695 24160 18788 24188
rect 18782 24148 18788 24160
rect 18840 24188 18846 24200
rect 20272 24188 20300 24216
rect 18840 24160 20300 24188
rect 57149 24191 57207 24197
rect 18840 24148 18846 24160
rect 57149 24157 57161 24191
rect 57195 24188 57207 24191
rect 58342 24188 58348 24200
rect 57195 24160 58348 24188
rect 57195 24157 57207 24160
rect 57149 24151 57207 24157
rect 58342 24148 58348 24160
rect 58400 24148 58406 24200
rect 3053 24123 3111 24129
rect 3053 24089 3065 24123
rect 3099 24120 3111 24123
rect 3694 24120 3700 24132
rect 3099 24092 3700 24120
rect 3099 24089 3111 24092
rect 3053 24083 3111 24089
rect 3694 24080 3700 24092
rect 3752 24120 3758 24132
rect 4525 24123 4583 24129
rect 4525 24120 4537 24123
rect 3752 24092 4537 24120
rect 3752 24080 3758 24092
rect 4525 24089 4537 24092
rect 4571 24089 4583 24123
rect 4525 24083 4583 24089
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 20073 24123 20131 24129
rect 20073 24120 20085 24123
rect 19392 24092 20085 24120
rect 19392 24080 19398 24092
rect 20073 24089 20085 24092
rect 20119 24089 20131 24123
rect 20073 24083 20131 24089
rect 1670 24052 1676 24064
rect 1631 24024 1676 24052
rect 1670 24012 1676 24024
rect 1728 24012 1734 24064
rect 3418 24052 3424 24064
rect 3379 24024 3424 24052
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 3510 24012 3516 24064
rect 3568 24052 3574 24064
rect 3970 24052 3976 24064
rect 3568 24024 3976 24052
rect 3568 24012 3574 24024
rect 3970 24012 3976 24024
rect 4028 24052 4034 24064
rect 4065 24055 4123 24061
rect 4065 24052 4077 24055
rect 4028 24024 4077 24052
rect 4028 24012 4034 24024
rect 4065 24021 4077 24024
rect 4111 24052 4123 24055
rect 5166 24052 5172 24064
rect 4111 24024 5172 24052
rect 4111 24021 4123 24024
rect 4065 24015 4123 24021
rect 5166 24012 5172 24024
rect 5224 24012 5230 24064
rect 19978 24052 19984 24064
rect 19939 24024 19984 24052
rect 19978 24012 19984 24024
rect 20036 24012 20042 24064
rect 20254 24012 20260 24064
rect 20312 24052 20318 24064
rect 20809 24055 20867 24061
rect 20809 24052 20821 24055
rect 20312 24024 20821 24052
rect 20312 24012 20318 24024
rect 20809 24021 20821 24024
rect 20855 24021 20867 24055
rect 20809 24015 20867 24021
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 2774 23808 2780 23860
rect 2832 23848 2838 23860
rect 3513 23851 3571 23857
rect 3513 23848 3525 23851
rect 2832 23820 3525 23848
rect 2832 23808 2838 23820
rect 3513 23817 3525 23820
rect 3559 23817 3571 23851
rect 3513 23811 3571 23817
rect 19521 23851 19579 23857
rect 19521 23817 19533 23851
rect 19567 23848 19579 23851
rect 19978 23848 19984 23860
rect 19567 23820 19984 23848
rect 19567 23817 19579 23820
rect 19521 23811 19579 23817
rect 19978 23808 19984 23820
rect 20036 23808 20042 23860
rect 58345 23851 58403 23857
rect 58345 23817 58357 23851
rect 58391 23848 58403 23851
rect 58802 23848 58808 23860
rect 58391 23820 58808 23848
rect 58391 23817 58403 23820
rect 58345 23811 58403 23817
rect 58802 23808 58808 23820
rect 58860 23808 58866 23860
rect 2038 23740 2044 23792
rect 2096 23780 2102 23792
rect 2225 23783 2283 23789
rect 2225 23780 2237 23783
rect 2096 23752 2237 23780
rect 2096 23740 2102 23752
rect 2225 23749 2237 23752
rect 2271 23749 2283 23783
rect 2225 23743 2283 23749
rect 2406 23740 2412 23792
rect 2464 23780 2470 23792
rect 14274 23780 14280 23792
rect 2464 23752 14280 23780
rect 2464 23740 2470 23752
rect 14274 23740 14280 23752
rect 14332 23740 14338 23792
rect 2317 23715 2375 23721
rect 2317 23681 2329 23715
rect 2363 23712 2375 23715
rect 2774 23712 2780 23724
rect 2363 23684 2780 23712
rect 2363 23681 2375 23684
rect 2317 23675 2375 23681
rect 2774 23672 2780 23684
rect 2832 23672 2838 23724
rect 4890 23672 4896 23724
rect 4948 23712 4954 23724
rect 6178 23712 6184 23724
rect 4948 23684 6184 23712
rect 4948 23672 4954 23684
rect 6178 23672 6184 23684
rect 6236 23672 6242 23724
rect 18601 23715 18659 23721
rect 18601 23681 18613 23715
rect 18647 23712 18659 23715
rect 19426 23712 19432 23724
rect 18647 23684 19432 23712
rect 18647 23681 18659 23684
rect 18601 23675 18659 23681
rect 19426 23672 19432 23684
rect 19484 23672 19490 23724
rect 2133 23647 2191 23653
rect 2133 23613 2145 23647
rect 2179 23613 2191 23647
rect 2133 23607 2191 23613
rect 2148 23576 2176 23607
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 5902 23644 5908 23656
rect 4028 23616 5908 23644
rect 4028 23604 4034 23616
rect 5902 23604 5908 23616
rect 5960 23604 5966 23656
rect 6086 23604 6092 23656
rect 6144 23644 6150 23656
rect 6144 23616 6914 23644
rect 6144 23604 6150 23616
rect 2406 23576 2412 23588
rect 2148 23548 2412 23576
rect 2406 23536 2412 23548
rect 2464 23576 2470 23588
rect 4157 23579 4215 23585
rect 4157 23576 4169 23579
rect 2464 23548 4169 23576
rect 2464 23536 2470 23548
rect 4157 23545 4169 23548
rect 4203 23576 4215 23579
rect 6886 23576 6914 23616
rect 17954 23576 17960 23588
rect 4203 23548 5948 23576
rect 6886 23548 17960 23576
rect 4203 23545 4215 23548
rect 4157 23539 4215 23545
rect 2314 23468 2320 23520
rect 2372 23508 2378 23520
rect 2685 23511 2743 23517
rect 2685 23508 2697 23511
rect 2372 23480 2697 23508
rect 2372 23468 2378 23480
rect 2685 23477 2697 23480
rect 2731 23477 2743 23511
rect 5920 23508 5948 23548
rect 17954 23536 17960 23548
rect 18012 23576 18018 23588
rect 18598 23576 18604 23588
rect 18012 23548 18604 23576
rect 18012 23536 18018 23548
rect 18598 23536 18604 23548
rect 18656 23536 18662 23588
rect 10410 23508 10416 23520
rect 5920 23480 10416 23508
rect 2685 23471 2743 23477
rect 10410 23468 10416 23480
rect 10468 23468 10474 23520
rect 18414 23508 18420 23520
rect 18375 23480 18420 23508
rect 18414 23468 18420 23480
rect 18472 23468 18478 23520
rect 20070 23468 20076 23520
rect 20128 23508 20134 23520
rect 20257 23511 20315 23517
rect 20257 23508 20269 23511
rect 20128 23480 20269 23508
rect 20128 23468 20134 23480
rect 20257 23477 20269 23480
rect 20303 23477 20315 23511
rect 20257 23471 20315 23477
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 16022 23304 16028 23316
rect 15983 23276 16028 23304
rect 16022 23264 16028 23276
rect 16080 23304 16086 23316
rect 18785 23307 18843 23313
rect 18785 23304 18797 23307
rect 16080 23276 18797 23304
rect 16080 23264 16086 23276
rect 18785 23273 18797 23276
rect 18831 23273 18843 23307
rect 19426 23304 19432 23316
rect 19387 23276 19432 23304
rect 18785 23267 18843 23273
rect 2501 23239 2559 23245
rect 2501 23205 2513 23239
rect 2547 23236 2559 23239
rect 4890 23236 4896 23248
rect 2547 23208 4896 23236
rect 2547 23205 2559 23208
rect 2501 23199 2559 23205
rect 4890 23196 4896 23208
rect 4948 23196 4954 23248
rect 16482 23128 16488 23180
rect 16540 23168 16546 23180
rect 17773 23171 17831 23177
rect 17773 23168 17785 23171
rect 16540 23140 17785 23168
rect 16540 23128 16546 23140
rect 17773 23137 17785 23140
rect 17819 23137 17831 23171
rect 18800 23168 18828 23267
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 58161 23307 58219 23313
rect 58161 23273 58173 23307
rect 58207 23304 58219 23307
rect 58710 23304 58716 23316
rect 58207 23276 58716 23304
rect 58207 23273 58219 23276
rect 58161 23267 58219 23273
rect 58710 23264 58716 23276
rect 58768 23264 58774 23316
rect 19889 23171 19947 23177
rect 19889 23168 19901 23171
rect 18800 23140 19901 23168
rect 17773 23131 17831 23137
rect 19889 23137 19901 23140
rect 19935 23137 19947 23171
rect 20070 23168 20076 23180
rect 20031 23140 20076 23168
rect 19889 23131 19947 23137
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 1857 23103 1915 23109
rect 1857 23069 1869 23103
rect 1903 23069 1915 23103
rect 2314 23100 2320 23112
rect 2275 23072 2320 23100
rect 1857 23063 1915 23069
rect 1872 23032 1900 23063
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 3973 23103 4031 23109
rect 3973 23100 3985 23103
rect 3476 23072 3985 23100
rect 3476 23060 3482 23072
rect 3973 23069 3985 23072
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 57701 23103 57759 23109
rect 57701 23069 57713 23103
rect 57747 23100 57759 23103
rect 58342 23100 58348 23112
rect 57747 23072 58348 23100
rect 57747 23069 57759 23072
rect 57701 23063 57759 23069
rect 58342 23060 58348 23072
rect 58400 23060 58406 23112
rect 9950 23032 9956 23044
rect 1872 23004 9956 23032
rect 9950 22992 9956 23004
rect 10008 23032 10014 23044
rect 10870 23032 10876 23044
rect 10008 23004 10876 23032
rect 10008 22992 10014 23004
rect 10870 22992 10876 23004
rect 10928 22992 10934 23044
rect 14826 22992 14832 23044
rect 14884 23032 14890 23044
rect 17497 23035 17555 23041
rect 14884 23004 16330 23032
rect 14884 22992 14890 23004
rect 17497 23001 17509 23035
rect 17543 23032 17555 23035
rect 18414 23032 18420 23044
rect 17543 23004 18420 23032
rect 17543 23001 17555 23004
rect 17497 22995 17555 23001
rect 18414 22992 18420 23004
rect 18472 22992 18478 23044
rect 1670 22964 1676 22976
rect 1631 22936 1676 22964
rect 1670 22924 1676 22936
rect 1728 22924 1734 22976
rect 2774 22924 2780 22976
rect 2832 22964 2838 22976
rect 3053 22967 3111 22973
rect 3053 22964 3065 22967
rect 2832 22936 3065 22964
rect 2832 22924 2838 22936
rect 3053 22933 3065 22936
rect 3099 22964 3111 22967
rect 3970 22964 3976 22976
rect 3099 22936 3976 22964
rect 3099 22933 3111 22936
rect 3053 22927 3111 22933
rect 3970 22924 3976 22936
rect 4028 22924 4034 22976
rect 4157 22967 4215 22973
rect 4157 22933 4169 22967
rect 4203 22964 4215 22967
rect 4798 22964 4804 22976
rect 4203 22936 4804 22964
rect 4203 22933 4215 22936
rect 4157 22927 4215 22933
rect 4798 22924 4804 22936
rect 4856 22924 4862 22976
rect 19797 22967 19855 22973
rect 19797 22933 19809 22967
rect 19843 22964 19855 22967
rect 19978 22964 19984 22976
rect 19843 22936 19984 22964
rect 19843 22933 19855 22936
rect 19797 22927 19855 22933
rect 19978 22924 19984 22936
rect 20036 22964 20042 22976
rect 20625 22967 20683 22973
rect 20625 22964 20637 22967
rect 20036 22936 20637 22964
rect 20036 22924 20042 22936
rect 20625 22933 20637 22936
rect 20671 22933 20683 22967
rect 20625 22927 20683 22933
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 2317 22763 2375 22769
rect 2317 22729 2329 22763
rect 2363 22760 2375 22763
rect 2774 22760 2780 22772
rect 2363 22732 2780 22760
rect 2363 22729 2375 22732
rect 2317 22723 2375 22729
rect 2774 22720 2780 22732
rect 2832 22760 2838 22772
rect 3694 22760 3700 22772
rect 2832 22732 3700 22760
rect 2832 22720 2838 22732
rect 3694 22720 3700 22732
rect 3752 22720 3758 22772
rect 8297 22763 8355 22769
rect 8297 22729 8309 22763
rect 8343 22760 8355 22763
rect 8478 22760 8484 22772
rect 8343 22732 8484 22760
rect 8343 22729 8355 22732
rect 8297 22723 8355 22729
rect 8478 22720 8484 22732
rect 8536 22720 8542 22772
rect 18598 22760 18604 22772
rect 18559 22732 18604 22760
rect 18598 22720 18604 22732
rect 18656 22720 18662 22772
rect 56134 22720 56140 22772
rect 56192 22760 56198 22772
rect 58161 22763 58219 22769
rect 58161 22760 58173 22763
rect 56192 22732 58173 22760
rect 56192 22720 56198 22732
rect 58161 22729 58173 22732
rect 58207 22729 58219 22763
rect 58161 22723 58219 22729
rect 2225 22695 2283 22701
rect 2225 22661 2237 22695
rect 2271 22692 2283 22695
rect 2590 22692 2596 22704
rect 2271 22664 2596 22692
rect 2271 22661 2283 22664
rect 2225 22655 2283 22661
rect 2590 22652 2596 22664
rect 2648 22692 2654 22704
rect 3145 22695 3203 22701
rect 3145 22692 3157 22695
rect 2648 22664 3157 22692
rect 2648 22652 2654 22664
rect 3145 22661 3157 22664
rect 3191 22692 3203 22695
rect 3191 22664 6914 22692
rect 3191 22661 3203 22664
rect 3145 22655 3203 22661
rect 2130 22556 2136 22568
rect 2091 22528 2136 22556
rect 2130 22516 2136 22528
rect 2188 22516 2194 22568
rect 2590 22380 2596 22432
rect 2648 22420 2654 22432
rect 2685 22423 2743 22429
rect 2685 22420 2697 22423
rect 2648 22392 2697 22420
rect 2648 22380 2654 22392
rect 2685 22389 2697 22392
rect 2731 22389 2743 22423
rect 6886 22420 6914 22664
rect 8386 22652 8392 22704
rect 8444 22692 8450 22704
rect 8444 22664 8602 22692
rect 8444 22652 8450 22664
rect 13906 22652 13912 22704
rect 13964 22692 13970 22704
rect 13964 22664 17618 22692
rect 13964 22652 13970 22664
rect 10042 22584 10048 22636
rect 10100 22624 10106 22636
rect 57517 22627 57575 22633
rect 10100 22596 10145 22624
rect 10100 22584 10106 22596
rect 57517 22593 57529 22627
rect 57563 22624 57575 22627
rect 58342 22624 58348 22636
rect 57563 22596 58348 22624
rect 57563 22593 57575 22596
rect 57517 22587 57575 22593
rect 58342 22584 58348 22596
rect 58400 22584 58406 22636
rect 8754 22516 8760 22568
rect 8812 22556 8818 22568
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 8812 22528 9781 22556
rect 8812 22516 8818 22528
rect 9769 22525 9781 22528
rect 9815 22525 9827 22559
rect 9769 22519 9827 22525
rect 15378 22516 15384 22568
rect 15436 22556 15442 22568
rect 16482 22556 16488 22568
rect 15436 22528 16488 22556
rect 15436 22516 15442 22528
rect 16482 22516 16488 22528
rect 16540 22556 16546 22568
rect 16853 22559 16911 22565
rect 16853 22556 16865 22559
rect 16540 22528 16865 22556
rect 16540 22516 16546 22528
rect 16853 22525 16865 22528
rect 16899 22525 16911 22559
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 16853 22519 16911 22525
rect 16960 22528 17141 22556
rect 16574 22448 16580 22500
rect 16632 22488 16638 22500
rect 16960 22488 16988 22528
rect 17129 22525 17141 22528
rect 17175 22525 17187 22559
rect 17129 22519 17187 22525
rect 19245 22559 19303 22565
rect 19245 22525 19257 22559
rect 19291 22556 19303 22559
rect 19426 22556 19432 22568
rect 19291 22528 19432 22556
rect 19291 22525 19303 22528
rect 19245 22519 19303 22525
rect 19426 22516 19432 22528
rect 19484 22516 19490 22568
rect 19521 22559 19579 22565
rect 19521 22525 19533 22559
rect 19567 22525 19579 22559
rect 19521 22519 19579 22525
rect 16632 22460 16988 22488
rect 16632 22448 16638 22460
rect 18138 22448 18144 22500
rect 18196 22488 18202 22500
rect 19536 22488 19564 22519
rect 18196 22460 19564 22488
rect 18196 22448 18202 22460
rect 10410 22420 10416 22432
rect 6886 22392 10416 22420
rect 2685 22383 2743 22389
rect 10410 22380 10416 22392
rect 10468 22380 10474 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1670 22216 1676 22228
rect 1631 22188 1676 22216
rect 1670 22176 1676 22188
rect 1728 22176 1734 22228
rect 8570 22176 8576 22228
rect 8628 22216 8634 22228
rect 13001 22219 13059 22225
rect 13001 22216 13013 22219
rect 8628 22188 13013 22216
rect 8628 22176 8634 22188
rect 13001 22185 13013 22188
rect 13047 22185 13059 22219
rect 13001 22179 13059 22185
rect 16298 22176 16304 22228
rect 16356 22216 16362 22228
rect 18138 22216 18144 22228
rect 16356 22188 18144 22216
rect 16356 22176 16362 22188
rect 18138 22176 18144 22188
rect 18196 22176 18202 22228
rect 19426 22176 19432 22228
rect 19484 22216 19490 22228
rect 19613 22219 19671 22225
rect 19613 22216 19625 22219
rect 19484 22188 19625 22216
rect 19484 22176 19490 22188
rect 19613 22185 19625 22188
rect 19659 22185 19671 22219
rect 19613 22179 19671 22185
rect 2130 22040 2136 22092
rect 2188 22080 2194 22092
rect 2682 22080 2688 22092
rect 2188 22052 2688 22080
rect 2188 22040 2194 22052
rect 2682 22040 2688 22052
rect 2740 22080 2746 22092
rect 2777 22083 2835 22089
rect 2777 22080 2789 22083
rect 2740 22052 2789 22080
rect 2740 22040 2746 22052
rect 2777 22049 2789 22052
rect 2823 22049 2835 22083
rect 2777 22043 2835 22049
rect 7098 22040 7104 22092
rect 7156 22080 7162 22092
rect 11517 22083 11575 22089
rect 11517 22080 11529 22083
rect 7156 22052 11529 22080
rect 7156 22040 7162 22052
rect 11517 22049 11529 22052
rect 11563 22049 11575 22083
rect 11517 22043 11575 22049
rect 13265 22083 13323 22089
rect 13265 22049 13277 22083
rect 13311 22080 13323 22083
rect 15378 22080 15384 22092
rect 13311 22052 15384 22080
rect 13311 22049 13323 22052
rect 13265 22043 13323 22049
rect 15378 22040 15384 22052
rect 15436 22040 15442 22092
rect 20070 22040 20076 22092
rect 20128 22080 20134 22092
rect 20257 22083 20315 22089
rect 20257 22080 20269 22083
rect 20128 22052 20269 22080
rect 20128 22040 20134 22052
rect 20257 22049 20269 22052
rect 20303 22080 20315 22083
rect 20622 22080 20628 22092
rect 20303 22052 20628 22080
rect 20303 22049 20315 22052
rect 20257 22043 20315 22049
rect 20622 22040 20628 22052
rect 20680 22040 20686 22092
rect 56502 22040 56508 22092
rect 56560 22080 56566 22092
rect 58253 22083 58311 22089
rect 58253 22080 58265 22083
rect 56560 22052 58265 22080
rect 56560 22040 56566 22052
rect 58253 22049 58265 22052
rect 58299 22049 58311 22083
rect 58253 22043 58311 22049
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 21981 1915 22015
rect 1857 21975 1915 21981
rect 18877 22015 18935 22021
rect 18877 21981 18889 22015
rect 18923 22012 18935 22015
rect 19150 22012 19156 22024
rect 18923 21984 19156 22012
rect 18923 21981 18935 21984
rect 18877 21975 18935 21981
rect 1872 21944 1900 21975
rect 19150 21972 19156 21984
rect 19208 22012 19214 22024
rect 19981 22015 20039 22021
rect 19981 22012 19993 22015
rect 19208 21984 19993 22012
rect 19208 21972 19214 21984
rect 19981 21981 19993 21984
rect 20027 22012 20039 22015
rect 20162 22012 20168 22024
rect 20027 21984 20168 22012
rect 20027 21981 20039 21984
rect 19981 21975 20039 21981
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 57974 22012 57980 22024
rect 57935 21984 57980 22012
rect 57974 21972 57980 21984
rect 58032 21972 58038 22024
rect 3421 21947 3479 21953
rect 3421 21944 3433 21947
rect 1872 21916 3433 21944
rect 3421 21913 3433 21916
rect 3467 21944 3479 21947
rect 10686 21944 10692 21956
rect 3467 21916 10692 21944
rect 3467 21913 3479 21916
rect 3421 21907 3479 21913
rect 10686 21904 10692 21916
rect 10744 21904 10750 21956
rect 12558 21916 12940 21944
rect 12342 21836 12348 21888
rect 12400 21876 12406 21888
rect 12636 21876 12664 21916
rect 12400 21848 12664 21876
rect 12912 21876 12940 21916
rect 16206 21904 16212 21956
rect 16264 21944 16270 21956
rect 18325 21947 18383 21953
rect 18325 21944 18337 21947
rect 16264 21916 18337 21944
rect 16264 21904 16270 21916
rect 18325 21913 18337 21916
rect 18371 21944 18383 21947
rect 20073 21947 20131 21953
rect 20073 21944 20085 21947
rect 18371 21916 20085 21944
rect 18371 21913 18383 21916
rect 18325 21907 18383 21913
rect 20073 21913 20085 21916
rect 20119 21913 20131 21947
rect 20073 21907 20131 21913
rect 14826 21876 14832 21888
rect 12912 21848 14832 21876
rect 12400 21836 12406 21848
rect 14826 21836 14832 21848
rect 14884 21836 14890 21888
rect 20622 21836 20628 21888
rect 20680 21876 20686 21888
rect 20809 21879 20867 21885
rect 20809 21876 20821 21879
rect 20680 21848 20821 21876
rect 20680 21836 20686 21848
rect 20809 21845 20821 21848
rect 20855 21845 20867 21879
rect 20809 21839 20867 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 19058 21632 19064 21684
rect 19116 21672 19122 21684
rect 19429 21675 19487 21681
rect 19429 21672 19441 21675
rect 19116 21644 19441 21672
rect 19116 21632 19122 21644
rect 19429 21641 19441 21644
rect 19475 21641 19487 21675
rect 58158 21672 58164 21684
rect 58119 21644 58164 21672
rect 19429 21635 19487 21641
rect 58158 21632 58164 21644
rect 58216 21632 58222 21684
rect 2406 21604 2412 21616
rect 2056 21576 2412 21604
rect 2056 21477 2084 21576
rect 2406 21564 2412 21576
rect 2464 21564 2470 21616
rect 14737 21607 14795 21613
rect 14737 21573 14749 21607
rect 14783 21604 14795 21607
rect 15378 21604 15384 21616
rect 14783 21576 15384 21604
rect 14783 21573 14795 21576
rect 14737 21567 14795 21573
rect 15378 21564 15384 21576
rect 15436 21564 15442 21616
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21536 2375 21539
rect 3234 21536 3240 21548
rect 2363 21508 3240 21536
rect 2363 21505 2375 21508
rect 2317 21499 2375 21505
rect 3234 21496 3240 21508
rect 3292 21496 3298 21548
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 12492 21508 13001 21536
rect 12492 21496 12498 21508
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 18690 21496 18696 21548
rect 18748 21536 18754 21548
rect 19337 21539 19395 21545
rect 19337 21536 19349 21539
rect 18748 21508 19349 21536
rect 18748 21496 18754 21508
rect 19337 21505 19349 21508
rect 19383 21505 19395 21539
rect 19337 21499 19395 21505
rect 57517 21539 57575 21545
rect 57517 21505 57529 21539
rect 57563 21536 57575 21539
rect 58342 21536 58348 21548
rect 57563 21508 58348 21536
rect 57563 21505 57575 21508
rect 57517 21499 57575 21505
rect 58342 21496 58348 21508
rect 58400 21496 58406 21548
rect 2041 21471 2099 21477
rect 2041 21437 2053 21471
rect 2087 21437 2099 21471
rect 2222 21468 2228 21480
rect 2183 21440 2228 21468
rect 2041 21431 2099 21437
rect 2222 21428 2228 21440
rect 2280 21428 2286 21480
rect 19613 21471 19671 21477
rect 19613 21437 19625 21471
rect 19659 21468 19671 21471
rect 19659 21440 20300 21468
rect 19659 21437 19671 21440
rect 19613 21431 19671 21437
rect 1946 21360 1952 21412
rect 2004 21400 2010 21412
rect 14366 21400 14372 21412
rect 2004 21372 14372 21400
rect 2004 21360 2010 21372
rect 14366 21360 14372 21372
rect 14424 21360 14430 21412
rect 20272 21344 20300 21440
rect 2314 21292 2320 21344
rect 2372 21332 2378 21344
rect 2685 21335 2743 21341
rect 2685 21332 2697 21335
rect 2372 21304 2697 21332
rect 2372 21292 2378 21304
rect 2685 21301 2697 21304
rect 2731 21301 2743 21335
rect 3234 21332 3240 21344
rect 3195 21304 3240 21332
rect 2685 21295 2743 21301
rect 3234 21292 3240 21304
rect 3292 21292 3298 21344
rect 12434 21332 12440 21344
rect 12395 21304 12440 21332
rect 12434 21292 12440 21304
rect 12492 21292 12498 21344
rect 18509 21335 18567 21341
rect 18509 21301 18521 21335
rect 18555 21332 18567 21335
rect 18690 21332 18696 21344
rect 18555 21304 18696 21332
rect 18555 21301 18567 21304
rect 18509 21295 18567 21301
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 18966 21332 18972 21344
rect 18927 21304 18972 21332
rect 18966 21292 18972 21304
rect 19024 21292 19030 21344
rect 20254 21332 20260 21344
rect 20215 21304 20260 21332
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1670 21128 1676 21140
rect 1631 21100 1676 21128
rect 1670 21088 1676 21100
rect 1728 21088 1734 21140
rect 2222 21088 2228 21140
rect 2280 21128 2286 21140
rect 3973 21131 4031 21137
rect 3973 21128 3985 21131
rect 2280 21100 3985 21128
rect 2280 21088 2286 21100
rect 3973 21097 3985 21100
rect 4019 21097 4031 21131
rect 3973 21091 4031 21097
rect 5810 21088 5816 21140
rect 5868 21128 5874 21140
rect 6825 21131 6883 21137
rect 6825 21128 6837 21131
rect 5868 21100 6837 21128
rect 5868 21088 5874 21100
rect 6825 21097 6837 21100
rect 6871 21097 6883 21131
rect 6825 21091 6883 21097
rect 8294 21088 8300 21140
rect 8352 21137 8358 21140
rect 8352 21131 8367 21137
rect 8355 21097 8367 21131
rect 14366 21128 14372 21140
rect 14327 21100 14372 21128
rect 8352 21091 8367 21097
rect 8352 21088 8358 21091
rect 14366 21088 14372 21100
rect 14424 21088 14430 21140
rect 18693 21131 18751 21137
rect 18693 21097 18705 21131
rect 18739 21128 18751 21131
rect 18874 21128 18880 21140
rect 18739 21100 18880 21128
rect 18739 21097 18751 21100
rect 18693 21091 18751 21097
rect 18874 21088 18880 21100
rect 18932 21128 18938 21140
rect 19058 21128 19064 21140
rect 18932 21100 19064 21128
rect 18932 21088 18938 21100
rect 19058 21088 19064 21100
rect 19116 21088 19122 21140
rect 58161 21131 58219 21137
rect 58161 21097 58173 21131
rect 58207 21128 58219 21131
rect 58250 21128 58256 21140
rect 58207 21100 58256 21128
rect 58207 21097 58219 21100
rect 58161 21091 58219 21097
rect 58250 21088 58256 21100
rect 58308 21088 58314 21140
rect 2501 21063 2559 21069
rect 2501 21029 2513 21063
rect 2547 21029 2559 21063
rect 2501 21023 2559 21029
rect 2516 20992 2544 21023
rect 5445 20995 5503 21001
rect 5445 20992 5457 20995
rect 2516 20964 5457 20992
rect 5445 20961 5457 20964
rect 5491 20961 5503 20995
rect 5718 20992 5724 21004
rect 5679 20964 5724 20992
rect 5445 20955 5503 20961
rect 5718 20952 5724 20964
rect 5776 20992 5782 21004
rect 8294 20992 8300 21004
rect 5776 20964 8300 20992
rect 5776 20952 5782 20964
rect 8294 20952 8300 20964
rect 8352 20992 8358 21004
rect 8573 20995 8631 21001
rect 8573 20992 8585 20995
rect 8352 20964 8585 20992
rect 8352 20952 8358 20964
rect 8573 20961 8585 20964
rect 8619 20992 8631 20995
rect 10042 20992 10048 21004
rect 8619 20964 10048 20992
rect 8619 20961 8631 20964
rect 8573 20955 8631 20961
rect 10042 20952 10048 20964
rect 10100 20952 10106 21004
rect 15378 20952 15384 21004
rect 15436 20992 15442 21004
rect 16114 20992 16120 21004
rect 15436 20964 16120 20992
rect 15436 20952 15442 20964
rect 16114 20952 16120 20964
rect 16172 20952 16178 21004
rect 1857 20927 1915 20933
rect 1857 20893 1869 20927
rect 1903 20924 1915 20927
rect 2038 20924 2044 20936
rect 1903 20896 2044 20924
rect 1903 20893 1915 20896
rect 1857 20887 1915 20893
rect 2038 20884 2044 20896
rect 2096 20884 2102 20936
rect 2314 20924 2320 20936
rect 2275 20896 2320 20924
rect 2314 20884 2320 20896
rect 2372 20884 2378 20936
rect 2406 20884 2412 20936
rect 2464 20924 2470 20936
rect 2961 20927 3019 20933
rect 2961 20924 2973 20927
rect 2464 20896 2973 20924
rect 2464 20884 2470 20896
rect 2961 20893 2973 20896
rect 3007 20893 3019 20927
rect 2961 20887 3019 20893
rect 57701 20927 57759 20933
rect 57701 20893 57713 20927
rect 57747 20924 57759 20927
rect 58342 20924 58348 20936
rect 57747 20896 58348 20924
rect 57747 20893 57759 20896
rect 57701 20887 57759 20893
rect 58342 20884 58348 20896
rect 58400 20884 58406 20936
rect 1946 20816 1952 20868
rect 2004 20856 2010 20868
rect 2424 20856 2452 20884
rect 2004 20828 2452 20856
rect 2004 20816 2010 20828
rect 4982 20816 4988 20868
rect 5040 20856 5046 20868
rect 5040 20828 6914 20856
rect 7866 20828 7972 20856
rect 5040 20816 5046 20828
rect 6886 20788 6914 20828
rect 7944 20788 7972 20828
rect 14826 20816 14832 20868
rect 14884 20816 14890 20868
rect 15841 20859 15899 20865
rect 15841 20825 15853 20859
rect 15887 20856 15899 20859
rect 16942 20856 16948 20868
rect 15887 20828 16948 20856
rect 15887 20825 15899 20828
rect 15841 20819 15899 20825
rect 16942 20816 16948 20828
rect 17000 20816 17006 20868
rect 8386 20788 8392 20800
rect 6886 20760 8392 20788
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 11882 20788 11888 20800
rect 11843 20760 11888 20788
rect 11882 20748 11888 20760
rect 11940 20748 11946 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 1670 20584 1676 20596
rect 1631 20556 1676 20584
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 2682 20544 2688 20596
rect 2740 20584 2746 20596
rect 2777 20587 2835 20593
rect 2777 20584 2789 20587
rect 2740 20556 2789 20584
rect 2740 20544 2746 20556
rect 2777 20553 2789 20556
rect 2823 20553 2835 20587
rect 8294 20584 8300 20596
rect 8255 20556 8300 20584
rect 2777 20547 2835 20553
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 14274 20584 14280 20596
rect 14235 20556 14280 20584
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 4982 20516 4988 20528
rect 4943 20488 4988 20516
rect 4982 20476 4988 20488
rect 5040 20476 5046 20528
rect 11882 20516 11888 20528
rect 6886 20488 11888 20516
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20448 1915 20451
rect 2222 20448 2228 20460
rect 1903 20420 2228 20448
rect 1903 20417 1915 20420
rect 1857 20411 1915 20417
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 5169 20451 5227 20457
rect 5169 20417 5181 20451
rect 5215 20448 5227 20451
rect 5810 20448 5816 20460
rect 5215 20420 5816 20448
rect 5215 20417 5227 20420
rect 5169 20411 5227 20417
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 5810 20244 5816 20256
rect 5771 20216 5816 20244
rect 5810 20204 5816 20216
rect 5868 20244 5874 20256
rect 6886 20244 6914 20488
rect 11882 20476 11888 20488
rect 11940 20516 11946 20528
rect 12161 20519 12219 20525
rect 12161 20516 12173 20519
rect 11940 20488 12173 20516
rect 11940 20476 11946 20488
rect 12161 20485 12173 20488
rect 12207 20485 12219 20519
rect 12342 20516 12348 20528
rect 12303 20488 12348 20516
rect 12161 20479 12219 20485
rect 12342 20476 12348 20488
rect 12400 20476 12406 20528
rect 13906 20476 13912 20528
rect 13964 20516 13970 20528
rect 13964 20488 14582 20516
rect 13964 20476 13970 20488
rect 18690 20476 18696 20528
rect 18748 20516 18754 20528
rect 19153 20519 19211 20525
rect 19153 20516 19165 20519
rect 18748 20488 19165 20516
rect 18748 20476 18754 20488
rect 19153 20485 19165 20488
rect 19199 20485 19211 20519
rect 20346 20516 20352 20528
rect 20307 20488 20352 20516
rect 19153 20479 19211 20485
rect 20346 20476 20352 20488
rect 20404 20476 20410 20528
rect 9585 20451 9643 20457
rect 9585 20417 9597 20451
rect 9631 20448 9643 20451
rect 16025 20451 16083 20457
rect 9631 20420 10180 20448
rect 9631 20417 9643 20420
rect 9585 20411 9643 20417
rect 10152 20321 10180 20420
rect 16025 20417 16037 20451
rect 16071 20448 16083 20451
rect 16114 20448 16120 20460
rect 16071 20420 16120 20448
rect 16071 20417 16083 20420
rect 16025 20411 16083 20417
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20448 18383 20451
rect 18966 20448 18972 20460
rect 18371 20420 18972 20448
rect 18371 20417 18383 20420
rect 18325 20411 18383 20417
rect 18966 20408 18972 20420
rect 19024 20408 19030 20460
rect 20622 20448 20628 20460
rect 19444 20420 20628 20448
rect 19444 20392 19472 20420
rect 20622 20408 20628 20420
rect 20680 20448 20686 20460
rect 21085 20451 21143 20457
rect 21085 20448 21097 20451
rect 20680 20420 21097 20448
rect 20680 20408 20686 20420
rect 21085 20417 21097 20420
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 15749 20383 15807 20389
rect 15749 20349 15761 20383
rect 15795 20380 15807 20383
rect 17310 20380 17316 20392
rect 15795 20352 17316 20380
rect 15795 20349 15807 20352
rect 15749 20343 15807 20349
rect 17310 20340 17316 20352
rect 17368 20340 17374 20392
rect 19245 20383 19303 20389
rect 19245 20380 19257 20383
rect 17604 20352 19257 20380
rect 10137 20315 10195 20321
rect 10137 20281 10149 20315
rect 10183 20312 10195 20315
rect 12434 20312 12440 20324
rect 10183 20284 12440 20312
rect 10183 20281 10195 20284
rect 10137 20275 10195 20281
rect 12434 20272 12440 20284
rect 12492 20272 12498 20324
rect 17604 20256 17632 20352
rect 19245 20349 19257 20352
rect 19291 20349 19303 20383
rect 19426 20380 19432 20392
rect 19387 20352 19432 20380
rect 19245 20343 19303 20349
rect 19426 20340 19432 20352
rect 19484 20340 19490 20392
rect 5868 20216 6914 20244
rect 5868 20204 5874 20216
rect 14366 20204 14372 20256
rect 14424 20244 14430 20256
rect 17218 20244 17224 20256
rect 14424 20216 17224 20244
rect 14424 20204 14430 20216
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 17586 20244 17592 20256
rect 17547 20216 17592 20244
rect 17586 20204 17592 20216
rect 17644 20204 17650 20256
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 18141 20247 18199 20253
rect 18141 20244 18153 20247
rect 18104 20216 18153 20244
rect 18104 20204 18110 20216
rect 18141 20213 18153 20216
rect 18187 20213 18199 20247
rect 18782 20244 18788 20256
rect 18743 20216 18788 20244
rect 18141 20207 18199 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 6196 20012 16574 20040
rect 6196 19984 6224 20012
rect 6178 19972 6184 19984
rect 5552 19944 6184 19972
rect 2133 19907 2191 19913
rect 2133 19873 2145 19907
rect 2179 19904 2191 19907
rect 2682 19904 2688 19916
rect 2179 19876 2688 19904
rect 2179 19873 2191 19876
rect 2133 19867 2191 19873
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 5552 19913 5580 19944
rect 6178 19932 6184 19944
rect 6236 19932 6242 19984
rect 12618 19972 12624 19984
rect 12579 19944 12624 19972
rect 12618 19932 12624 19944
rect 12676 19932 12682 19984
rect 5537 19907 5595 19913
rect 5537 19873 5549 19907
rect 5583 19873 5595 19907
rect 5537 19867 5595 19873
rect 7561 19907 7619 19913
rect 7561 19873 7573 19907
rect 7607 19904 7619 19907
rect 8294 19904 8300 19916
rect 7607 19876 8300 19904
rect 7607 19873 7619 19876
rect 7561 19867 7619 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 10042 19864 10048 19916
rect 10100 19904 10106 19916
rect 10873 19907 10931 19913
rect 10873 19904 10885 19907
rect 10100 19876 10885 19904
rect 10100 19864 10106 19876
rect 10873 19873 10885 19876
rect 10919 19873 10931 19907
rect 10873 19867 10931 19873
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19904 11207 19907
rect 11238 19904 11244 19916
rect 11195 19876 11244 19904
rect 11195 19873 11207 19876
rect 11149 19867 11207 19873
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 12342 19864 12348 19916
rect 12400 19864 12406 19916
rect 16546 19904 16574 20012
rect 19334 19904 19340 19916
rect 16546 19876 19340 19904
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 2317 19839 2375 19845
rect 2317 19805 2329 19839
rect 2363 19836 2375 19839
rect 3878 19836 3884 19848
rect 2363 19808 3884 19836
rect 2363 19805 2375 19808
rect 2317 19799 2375 19805
rect 3878 19796 3884 19808
rect 3936 19796 3942 19848
rect 4982 19796 4988 19848
rect 5040 19836 5046 19848
rect 12360 19836 12388 19864
rect 5040 19808 6210 19836
rect 12282 19808 12388 19836
rect 57701 19839 57759 19845
rect 5040 19796 5046 19808
rect 57701 19805 57713 19839
rect 57747 19836 57759 19839
rect 58342 19836 58348 19848
rect 57747 19808 58348 19836
rect 57747 19805 57759 19808
rect 57701 19799 57759 19805
rect 58342 19796 58348 19808
rect 58400 19796 58406 19848
rect 2130 19728 2136 19780
rect 2188 19768 2194 19780
rect 2225 19771 2283 19777
rect 2225 19768 2237 19771
rect 2188 19740 2237 19768
rect 2188 19728 2194 19740
rect 2225 19737 2237 19740
rect 2271 19768 2283 19771
rect 3145 19771 3203 19777
rect 3145 19768 3157 19771
rect 2271 19740 3157 19768
rect 2271 19737 2283 19740
rect 2225 19731 2283 19737
rect 3145 19737 3157 19740
rect 3191 19737 3203 19771
rect 3145 19731 3203 19737
rect 7285 19771 7343 19777
rect 7285 19737 7297 19771
rect 7331 19737 7343 19771
rect 7285 19731 7343 19737
rect 2406 19660 2412 19712
rect 2464 19700 2470 19712
rect 2685 19703 2743 19709
rect 2685 19700 2697 19703
rect 2464 19672 2697 19700
rect 2464 19660 2470 19672
rect 2685 19669 2697 19672
rect 2731 19669 2743 19703
rect 3160 19700 3188 19731
rect 4982 19700 4988 19712
rect 3160 19672 4988 19700
rect 2685 19663 2743 19669
rect 4982 19660 4988 19672
rect 5040 19660 5046 19712
rect 7300 19700 7328 19731
rect 14366 19700 14372 19712
rect 7300 19672 14372 19700
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 18690 19700 18696 19712
rect 18651 19672 18696 19700
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 19705 19703 19763 19709
rect 19705 19700 19717 19703
rect 19484 19672 19717 19700
rect 19484 19660 19490 19672
rect 19705 19669 19717 19672
rect 19751 19700 19763 19703
rect 20162 19700 20168 19712
rect 19751 19672 20168 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 58161 19703 58219 19709
rect 58161 19669 58173 19703
rect 58207 19700 58219 19703
rect 58618 19700 58624 19712
rect 58207 19672 58624 19700
rect 58207 19669 58219 19672
rect 58161 19663 58219 19669
rect 58618 19660 58624 19672
rect 58676 19660 58682 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 1670 19496 1676 19508
rect 1631 19468 1676 19496
rect 1670 19456 1676 19468
rect 1728 19456 1734 19508
rect 10502 19496 10508 19508
rect 10463 19468 10508 19496
rect 10502 19456 10508 19468
rect 10560 19456 10566 19508
rect 10870 19456 10876 19508
rect 10928 19496 10934 19508
rect 12713 19499 12771 19505
rect 12713 19496 12725 19499
rect 10928 19468 12725 19496
rect 10928 19456 10934 19468
rect 12713 19465 12725 19468
rect 12759 19465 12771 19499
rect 12713 19459 12771 19465
rect 13814 19456 13820 19508
rect 13872 19496 13878 19508
rect 17405 19499 17463 19505
rect 17405 19496 17417 19499
rect 13872 19468 17417 19496
rect 13872 19456 13878 19468
rect 17405 19465 17417 19468
rect 17451 19465 17463 19499
rect 17405 19459 17463 19465
rect 18601 19499 18659 19505
rect 18601 19465 18613 19499
rect 18647 19465 18659 19499
rect 18601 19459 18659 19465
rect 58161 19499 58219 19505
rect 58161 19465 58173 19499
rect 58207 19496 58219 19499
rect 58434 19496 58440 19508
rect 58207 19468 58440 19496
rect 58207 19465 58219 19468
rect 58161 19459 58219 19465
rect 8202 19388 8208 19440
rect 8260 19428 8266 19440
rect 13906 19428 13912 19440
rect 8260 19400 9522 19428
rect 13754 19400 13912 19428
rect 8260 19388 8266 19400
rect 13906 19388 13912 19400
rect 13964 19388 13970 19440
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 3053 19295 3111 19301
rect 3053 19261 3065 19295
rect 3099 19292 3111 19295
rect 3142 19292 3148 19304
rect 3099 19264 3148 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 3142 19252 3148 19264
rect 3200 19292 3206 19304
rect 3878 19292 3884 19304
rect 3200 19264 3884 19292
rect 3200 19252 3206 19264
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 7650 19252 7656 19304
rect 7708 19292 7714 19304
rect 8220 19292 8248 19388
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 8757 19363 8815 19369
rect 8757 19360 8769 19363
rect 8352 19332 8769 19360
rect 8352 19320 8358 19332
rect 8757 19329 8769 19332
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 15378 19360 15384 19372
rect 14507 19332 15384 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19360 17647 19363
rect 18616 19360 18644 19459
rect 58434 19456 58440 19468
rect 58492 19456 58498 19508
rect 17635 19332 18644 19360
rect 18969 19363 19027 19369
rect 17635 19329 17647 19332
rect 17589 19323 17647 19329
rect 18969 19329 18981 19363
rect 19015 19360 19027 19363
rect 19334 19360 19340 19372
rect 19015 19332 19340 19360
rect 19015 19329 19027 19332
rect 18969 19323 19027 19329
rect 19334 19320 19340 19332
rect 19392 19360 19398 19372
rect 58342 19360 58348 19372
rect 19392 19332 19932 19360
rect 58303 19332 58348 19360
rect 19392 19320 19398 19332
rect 9030 19292 9036 19304
rect 7708 19264 8248 19292
rect 8991 19264 9036 19292
rect 7708 19252 7714 19264
rect 9030 19252 9036 19264
rect 9088 19252 9094 19304
rect 14182 19292 14188 19304
rect 14143 19264 14188 19292
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 19904 19301 19932 19332
rect 58342 19320 58348 19332
rect 58400 19320 58406 19372
rect 19061 19295 19119 19301
rect 19061 19261 19073 19295
rect 19107 19261 19119 19295
rect 19061 19255 19119 19261
rect 19245 19295 19303 19301
rect 19245 19261 19257 19295
rect 19291 19261 19303 19295
rect 19245 19255 19303 19261
rect 19889 19295 19947 19301
rect 19889 19261 19901 19295
rect 19935 19292 19947 19295
rect 19978 19292 19984 19304
rect 19935 19264 19984 19292
rect 19935 19261 19947 19264
rect 19889 19255 19947 19261
rect 18138 19156 18144 19168
rect 18099 19128 18144 19156
rect 18138 19116 18144 19128
rect 18196 19156 18202 19168
rect 19076 19156 19104 19255
rect 19260 19224 19288 19255
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20254 19224 20260 19236
rect 19260 19196 20260 19224
rect 20254 19184 20260 19196
rect 20312 19224 20318 19236
rect 20312 19196 20484 19224
rect 20312 19184 20318 19196
rect 20456 19165 20484 19196
rect 18196 19128 19104 19156
rect 20441 19159 20499 19165
rect 18196 19116 18202 19128
rect 20441 19125 20453 19159
rect 20487 19156 20499 19159
rect 20622 19156 20628 19168
rect 20487 19128 20628 19156
rect 20487 19125 20499 19128
rect 20441 19119 20499 19125
rect 20622 19116 20628 19128
rect 20680 19116 20686 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1670 18952 1676 18964
rect 1631 18924 1676 18952
rect 1670 18912 1676 18924
rect 1728 18912 1734 18964
rect 2498 18952 2504 18964
rect 2459 18924 2504 18952
rect 2498 18912 2504 18924
rect 2556 18912 2562 18964
rect 3053 18955 3111 18961
rect 3053 18921 3065 18955
rect 3099 18952 3111 18955
rect 3326 18952 3332 18964
rect 3099 18924 3332 18952
rect 3099 18921 3111 18924
rect 3053 18915 3111 18921
rect 3326 18912 3332 18924
rect 3384 18912 3390 18964
rect 16942 18952 16948 18964
rect 16903 18924 16948 18952
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 58342 18952 58348 18964
rect 58303 18924 58348 18952
rect 58342 18912 58348 18924
rect 58400 18912 58406 18964
rect 3602 18776 3608 18828
rect 3660 18816 3666 18828
rect 18138 18816 18144 18828
rect 3660 18788 18144 18816
rect 3660 18776 3666 18788
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 18230 18776 18236 18828
rect 18288 18816 18294 18828
rect 18601 18819 18659 18825
rect 18601 18816 18613 18819
rect 18288 18788 18613 18816
rect 18288 18776 18294 18788
rect 18601 18785 18613 18788
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 20073 18819 20131 18825
rect 20073 18785 20085 18819
rect 20119 18816 20131 18819
rect 20530 18816 20536 18828
rect 20119 18788 20536 18816
rect 20119 18785 20131 18788
rect 20073 18779 20131 18785
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18748 1915 18751
rect 2222 18748 2228 18760
rect 1903 18720 2228 18748
rect 1903 18717 1915 18720
rect 1857 18711 1915 18717
rect 2222 18708 2228 18720
rect 2280 18708 2286 18760
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18748 2375 18751
rect 2406 18748 2412 18760
rect 2363 18720 2412 18748
rect 2363 18717 2375 18720
rect 2317 18711 2375 18717
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 5258 18708 5264 18760
rect 5316 18748 5322 18760
rect 15838 18748 15844 18760
rect 5316 18720 15844 18748
rect 5316 18708 5322 18720
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 17126 18748 17132 18760
rect 17087 18720 17132 18748
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18748 18015 18751
rect 18782 18748 18788 18760
rect 18003 18720 18788 18748
rect 18003 18717 18015 18720
rect 17957 18711 18015 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 18877 18751 18935 18757
rect 18877 18717 18889 18751
rect 18923 18748 18935 18751
rect 20088 18748 20116 18779
rect 20530 18776 20536 18788
rect 20588 18776 20594 18828
rect 18923 18720 20116 18748
rect 18923 18717 18935 18720
rect 18877 18711 18935 18717
rect 5994 18640 6000 18692
rect 6052 18680 6058 18692
rect 11514 18680 11520 18692
rect 6052 18652 11520 18680
rect 6052 18640 6058 18652
rect 11514 18640 11520 18652
rect 11572 18640 11578 18692
rect 18690 18640 18696 18692
rect 18748 18680 18754 18692
rect 19797 18683 19855 18689
rect 19797 18680 19809 18683
rect 18748 18652 19809 18680
rect 18748 18640 18754 18652
rect 19797 18649 19809 18652
rect 19843 18680 19855 18683
rect 20254 18680 20260 18692
rect 19843 18652 20260 18680
rect 19843 18649 19855 18652
rect 19797 18643 19855 18649
rect 20254 18640 20260 18652
rect 20312 18640 20318 18692
rect 6822 18572 6828 18624
rect 6880 18612 6886 18624
rect 8110 18612 8116 18624
rect 6880 18584 8116 18612
rect 6880 18572 6886 18584
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 17773 18615 17831 18621
rect 17773 18612 17785 18615
rect 17092 18584 17785 18612
rect 17092 18572 17098 18584
rect 17773 18581 17785 18584
rect 17819 18581 17831 18615
rect 19426 18612 19432 18624
rect 19387 18584 19432 18612
rect 17773 18575 17831 18581
rect 19426 18572 19432 18584
rect 19484 18572 19490 18624
rect 19889 18615 19947 18621
rect 19889 18581 19901 18615
rect 19935 18612 19947 18615
rect 19978 18612 19984 18624
rect 19935 18584 19984 18612
rect 19935 18581 19947 18584
rect 19889 18575 19947 18581
rect 19978 18572 19984 18584
rect 20036 18612 20042 18624
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 20036 18584 20637 18612
rect 20036 18572 20042 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 1949 18411 2007 18417
rect 1949 18408 1961 18411
rect 1912 18380 1961 18408
rect 1912 18368 1918 18380
rect 1949 18377 1961 18380
rect 1995 18377 2007 18411
rect 2406 18408 2412 18420
rect 2367 18380 2412 18408
rect 1949 18371 2007 18377
rect 2406 18368 2412 18380
rect 2464 18368 2470 18420
rect 6638 18408 6644 18420
rect 6599 18380 6644 18408
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 6730 18368 6736 18420
rect 6788 18408 6794 18420
rect 13814 18408 13820 18420
rect 6788 18380 13820 18408
rect 6788 18368 6794 18380
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 17126 18368 17132 18420
rect 17184 18408 17190 18420
rect 18325 18411 18383 18417
rect 18325 18408 18337 18411
rect 17184 18380 18337 18408
rect 17184 18368 17190 18380
rect 18325 18377 18337 18380
rect 18371 18377 18383 18411
rect 18325 18371 18383 18377
rect 18693 18411 18751 18417
rect 18693 18377 18705 18411
rect 18739 18408 18751 18411
rect 19334 18408 19340 18420
rect 18739 18380 19340 18408
rect 18739 18377 18751 18380
rect 18693 18371 18751 18377
rect 19334 18368 19340 18380
rect 19392 18408 19398 18420
rect 19518 18408 19524 18420
rect 19392 18380 19524 18408
rect 19392 18368 19398 18380
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 2041 18343 2099 18349
rect 2041 18309 2053 18343
rect 2087 18340 2099 18343
rect 3326 18340 3332 18352
rect 2087 18312 3332 18340
rect 2087 18309 2099 18312
rect 2041 18303 2099 18309
rect 3326 18300 3332 18312
rect 3384 18300 3390 18352
rect 4186 18312 5304 18340
rect 5276 18272 5304 18312
rect 7650 18300 7656 18352
rect 7708 18300 7714 18352
rect 8110 18340 8116 18352
rect 8071 18312 8116 18340
rect 8110 18300 8116 18312
rect 8168 18300 8174 18352
rect 14458 18300 14464 18352
rect 14516 18340 14522 18352
rect 18785 18343 18843 18349
rect 18785 18340 18797 18343
rect 14516 18312 18797 18340
rect 14516 18300 14522 18312
rect 18785 18309 18797 18312
rect 18831 18340 18843 18343
rect 20073 18343 20131 18349
rect 20073 18340 20085 18343
rect 18831 18312 20085 18340
rect 18831 18309 18843 18312
rect 18785 18303 18843 18309
rect 20073 18309 20085 18312
rect 20119 18309 20131 18343
rect 20073 18303 20131 18309
rect 5534 18272 5540 18284
rect 5276 18244 5540 18272
rect 5534 18232 5540 18244
rect 5592 18272 5598 18284
rect 7098 18272 7104 18284
rect 5592 18244 7104 18272
rect 5592 18232 5598 18244
rect 7098 18232 7104 18244
rect 7156 18232 7162 18284
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 18138 18272 18144 18284
rect 17543 18244 18144 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 18138 18232 18144 18244
rect 18196 18232 18202 18284
rect 57517 18275 57575 18281
rect 57517 18241 57529 18275
rect 57563 18272 57575 18275
rect 58342 18272 58348 18284
rect 57563 18244 58348 18272
rect 57563 18241 57575 18244
rect 57517 18235 57575 18241
rect 58342 18232 58348 18244
rect 58400 18232 58406 18284
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18204 1915 18207
rect 1946 18204 1952 18216
rect 1903 18176 1952 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 3602 18204 3608 18216
rect 2915 18176 3608 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 3602 18164 3608 18176
rect 3660 18164 3666 18216
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 4893 18207 4951 18213
rect 4663 18176 4844 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 4816 18136 4844 18176
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 5902 18204 5908 18216
rect 4939 18176 5908 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 5902 18164 5908 18176
rect 5960 18204 5966 18216
rect 8389 18207 8447 18213
rect 8389 18204 8401 18207
rect 5960 18176 8401 18204
rect 5960 18164 5966 18176
rect 8389 18173 8401 18176
rect 8435 18204 8447 18207
rect 8662 18204 8668 18216
rect 8435 18176 8668 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 8662 18164 8668 18176
rect 8720 18164 8726 18216
rect 18969 18207 19027 18213
rect 18969 18173 18981 18207
rect 19015 18204 19027 18207
rect 19334 18204 19340 18216
rect 19015 18176 19340 18204
rect 19015 18173 19027 18176
rect 18969 18167 19027 18173
rect 19334 18164 19340 18176
rect 19392 18204 19398 18216
rect 20530 18204 20536 18216
rect 19392 18176 20536 18204
rect 19392 18164 19398 18176
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 6730 18136 6736 18148
rect 4816 18108 6736 18136
rect 6730 18096 6736 18108
rect 6788 18096 6794 18148
rect 17310 18136 17316 18148
rect 17271 18108 17316 18136
rect 17310 18096 17316 18108
rect 17368 18096 17374 18148
rect 7098 18028 7104 18080
rect 7156 18068 7162 18080
rect 7650 18068 7656 18080
rect 7156 18040 7656 18068
rect 7156 18028 7162 18040
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 19613 18071 19671 18077
rect 19613 18037 19625 18071
rect 19659 18068 19671 18071
rect 20254 18068 20260 18080
rect 19659 18040 20260 18068
rect 19659 18037 19671 18040
rect 19613 18031 19671 18037
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 58161 18071 58219 18077
rect 58161 18037 58173 18071
rect 58207 18068 58219 18071
rect 58802 18068 58808 18080
rect 58207 18040 58808 18068
rect 58207 18037 58219 18040
rect 58161 18031 58219 18037
rect 58802 18028 58808 18040
rect 58860 18028 58866 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1670 17864 1676 17876
rect 1631 17836 1676 17864
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 1946 17824 1952 17876
rect 2004 17864 2010 17876
rect 3053 17867 3111 17873
rect 3053 17864 3065 17867
rect 2004 17836 3065 17864
rect 2004 17824 2010 17836
rect 3053 17833 3065 17836
rect 3099 17833 3111 17867
rect 3053 17827 3111 17833
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 10045 17867 10103 17873
rect 10045 17864 10057 17867
rect 9916 17836 10057 17864
rect 9916 17824 9922 17836
rect 10045 17833 10057 17836
rect 10091 17833 10103 17867
rect 10045 17827 10103 17833
rect 11974 17824 11980 17876
rect 12032 17864 12038 17876
rect 17586 17864 17592 17876
rect 12032 17836 17592 17864
rect 12032 17824 12038 17836
rect 17586 17824 17592 17836
rect 17644 17824 17650 17876
rect 18138 17864 18144 17876
rect 18099 17836 18144 17864
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 19518 17864 19524 17876
rect 19479 17836 19524 17864
rect 19518 17824 19524 17836
rect 19576 17864 19582 17876
rect 20438 17864 20444 17876
rect 19576 17836 20444 17864
rect 19576 17824 19582 17836
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 11422 17688 11428 17740
rect 11480 17728 11486 17740
rect 11517 17731 11575 17737
rect 11517 17728 11529 17731
rect 11480 17700 11529 17728
rect 11480 17688 11486 17700
rect 11517 17697 11529 17700
rect 11563 17697 11575 17731
rect 15194 17728 15200 17740
rect 15155 17700 15200 17728
rect 11517 17691 11575 17697
rect 15194 17688 15200 17700
rect 15252 17728 15258 17740
rect 18506 17728 18512 17740
rect 15252 17700 18512 17728
rect 15252 17688 15258 17700
rect 18506 17688 18512 17700
rect 18564 17688 18570 17740
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 19334 17728 19340 17740
rect 18831 17700 19340 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 19334 17688 19340 17700
rect 19392 17688 19398 17740
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17660 1915 17663
rect 2498 17660 2504 17672
rect 1903 17632 2504 17660
rect 1903 17629 1915 17632
rect 1857 17623 1915 17629
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17660 2651 17663
rect 2682 17660 2688 17672
rect 2639 17632 2688 17660
rect 2639 17629 2651 17632
rect 2593 17623 2651 17629
rect 2682 17620 2688 17632
rect 2740 17620 2746 17672
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17660 11851 17663
rect 13814 17660 13820 17672
rect 11839 17632 13820 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 19150 17660 19156 17672
rect 17276 17632 17321 17660
rect 18524 17632 19156 17660
rect 17276 17620 17282 17632
rect 7650 17552 7656 17604
rect 7708 17592 7714 17604
rect 9674 17592 9680 17604
rect 7708 17564 9680 17592
rect 7708 17552 7714 17564
rect 9674 17552 9680 17564
rect 9732 17592 9738 17604
rect 9732 17564 10350 17592
rect 9732 17552 9738 17564
rect 13906 17552 13912 17604
rect 13964 17592 13970 17604
rect 15010 17592 15016 17604
rect 13964 17564 15016 17592
rect 13964 17552 13970 17564
rect 15010 17552 15016 17564
rect 15068 17592 15074 17604
rect 16945 17595 17003 17601
rect 15068 17564 15778 17592
rect 15068 17552 15074 17564
rect 16945 17561 16957 17595
rect 16991 17592 17003 17595
rect 17770 17592 17776 17604
rect 16991 17564 17776 17592
rect 16991 17561 17003 17564
rect 16945 17555 17003 17561
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 2406 17524 2412 17536
rect 2367 17496 2412 17524
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 14274 17484 14280 17536
rect 14332 17524 14338 17536
rect 17586 17524 17592 17536
rect 14332 17496 17592 17524
rect 14332 17484 14338 17496
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 18524 17533 18552 17632
rect 19150 17620 19156 17632
rect 19208 17620 19214 17672
rect 57701 17663 57759 17669
rect 57701 17629 57713 17663
rect 57747 17660 57759 17663
rect 58342 17660 58348 17672
rect 57747 17632 58348 17660
rect 57747 17629 57759 17632
rect 57701 17623 57759 17629
rect 58342 17620 58348 17632
rect 58400 17620 58406 17672
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17493 18567 17527
rect 18509 17487 18567 17493
rect 18598 17484 18604 17536
rect 18656 17524 18662 17536
rect 58161 17527 58219 17533
rect 18656 17496 18701 17524
rect 18656 17484 18662 17496
rect 58161 17493 58173 17527
rect 58207 17524 58219 17527
rect 58250 17524 58256 17536
rect 58207 17496 58256 17524
rect 58207 17493 58219 17496
rect 58161 17487 58219 17493
rect 58250 17484 58256 17496
rect 58308 17484 58314 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 2317 17323 2375 17329
rect 2317 17289 2329 17323
rect 2363 17320 2375 17323
rect 2774 17320 2780 17332
rect 2363 17292 2780 17320
rect 2363 17289 2375 17292
rect 2317 17283 2375 17289
rect 2774 17280 2780 17292
rect 2832 17320 2838 17332
rect 3789 17323 3847 17329
rect 3789 17320 3801 17323
rect 2832 17292 3801 17320
rect 2832 17280 2838 17292
rect 3789 17289 3801 17292
rect 3835 17289 3847 17323
rect 3789 17283 3847 17289
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 11974 17320 11980 17332
rect 7800 17292 11980 17320
rect 7800 17280 7806 17292
rect 11974 17280 11980 17292
rect 12032 17280 12038 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 17218 17320 17224 17332
rect 13872 17292 17224 17320
rect 13872 17280 13878 17292
rect 2225 17255 2283 17261
rect 2225 17221 2237 17255
rect 2271 17252 2283 17255
rect 2682 17252 2688 17264
rect 2271 17224 2688 17252
rect 2271 17221 2283 17224
rect 2225 17215 2283 17221
rect 2682 17212 2688 17224
rect 2740 17252 2746 17264
rect 8386 17252 8392 17264
rect 2740 17224 8392 17252
rect 2740 17212 2746 17224
rect 8386 17212 8392 17224
rect 8444 17212 8450 17264
rect 13906 17252 13912 17264
rect 13018 17224 13912 17252
rect 13906 17212 13912 17224
rect 13964 17252 13970 17264
rect 13964 17224 14490 17252
rect 13964 17212 13970 17224
rect 3145 17187 3203 17193
rect 3145 17184 3157 17187
rect 2700 17156 3157 17184
rect 1946 17076 1952 17128
rect 2004 17116 2010 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 2004 17088 2053 17116
rect 2004 17076 2010 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 2700 17057 2728 17156
rect 3145 17153 3157 17156
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17184 5411 17187
rect 5810 17184 5816 17196
rect 5399 17156 5816 17184
rect 5399 17153 5411 17156
rect 5353 17147 5411 17153
rect 5810 17144 5816 17156
rect 5868 17184 5874 17196
rect 6362 17184 6368 17196
rect 5868 17156 6368 17184
rect 5868 17144 5874 17156
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17184 13783 17187
rect 13814 17184 13820 17196
rect 13771 17156 13820 17184
rect 13771 17153 13783 17156
rect 13725 17147 13783 17153
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 15948 17193 15976 17292
rect 17218 17280 17224 17292
rect 17276 17280 17282 17332
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 17773 17323 17831 17329
rect 17773 17320 17785 17323
rect 17644 17292 17785 17320
rect 17644 17280 17650 17292
rect 17773 17289 17785 17292
rect 17819 17320 17831 17323
rect 18598 17320 18604 17332
rect 17819 17292 18604 17320
rect 17819 17289 17831 17292
rect 17773 17283 17831 17289
rect 18598 17280 18604 17292
rect 18656 17280 18662 17332
rect 18966 17280 18972 17332
rect 19024 17320 19030 17332
rect 19061 17323 19119 17329
rect 19061 17320 19073 17323
rect 19024 17292 19073 17320
rect 19024 17280 19030 17292
rect 19061 17289 19073 17292
rect 19107 17320 19119 17323
rect 19150 17320 19156 17332
rect 19107 17292 19156 17320
rect 19107 17289 19119 17292
rect 19061 17283 19119 17289
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17184 18475 17187
rect 19426 17184 19432 17196
rect 18463 17156 19432 17184
rect 18463 17153 18475 17156
rect 18417 17147 18475 17153
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 5534 17116 5540 17128
rect 5495 17088 5540 17116
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17116 13507 17119
rect 15657 17119 15715 17125
rect 13495 17088 14688 17116
rect 13495 17085 13507 17088
rect 13449 17079 13507 17085
rect 2685 17051 2743 17057
rect 2685 17017 2697 17051
rect 2731 17017 2743 17051
rect 2685 17011 2743 17017
rect 3329 17051 3387 17057
rect 3329 17017 3341 17051
rect 3375 17048 3387 17051
rect 9398 17048 9404 17060
rect 3375 17020 9404 17048
rect 3375 17017 3387 17020
rect 3329 17011 3387 17017
rect 9398 17008 9404 17020
rect 9456 17008 9462 17060
rect 14090 17008 14096 17060
rect 14148 17048 14154 17060
rect 14185 17051 14243 17057
rect 14185 17048 14197 17051
rect 14148 17020 14197 17048
rect 14148 17008 14154 17020
rect 14185 17017 14197 17020
rect 14231 17017 14243 17051
rect 14185 17011 14243 17017
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 5074 16980 5080 16992
rect 4856 16952 5080 16980
rect 4856 16940 4862 16952
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 6362 16940 6368 16992
rect 6420 16980 6426 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6420 16952 6561 16980
rect 6420 16940 6426 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 14660 16980 14688 17088
rect 15657 17085 15669 17119
rect 15703 17116 15715 17119
rect 17678 17116 17684 17128
rect 15703 17088 17684 17116
rect 15703 17085 15715 17088
rect 15657 17079 15715 17085
rect 17678 17076 17684 17088
rect 17736 17076 17742 17128
rect 17310 17008 17316 17060
rect 17368 17048 17374 17060
rect 18233 17051 18291 17057
rect 18233 17048 18245 17051
rect 17368 17020 18245 17048
rect 17368 17008 17374 17020
rect 18233 17017 18245 17020
rect 18279 17017 18291 17051
rect 18233 17011 18291 17017
rect 17034 16980 17040 16992
rect 14660 16952 17040 16980
rect 6549 16943 6607 16949
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1946 16736 1952 16788
rect 2004 16776 2010 16788
rect 2682 16776 2688 16788
rect 2004 16748 2688 16776
rect 2004 16736 2010 16748
rect 2682 16736 2688 16748
rect 2740 16776 2746 16788
rect 3053 16779 3111 16785
rect 3053 16776 3065 16779
rect 2740 16748 3065 16776
rect 2740 16736 2746 16748
rect 3053 16745 3065 16748
rect 3099 16745 3111 16779
rect 3053 16739 3111 16745
rect 13078 16736 13084 16788
rect 13136 16776 13142 16788
rect 17310 16776 17316 16788
rect 13136 16748 17316 16776
rect 13136 16736 13142 16748
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 17770 16776 17776 16788
rect 17731 16748 17776 16776
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 5074 16600 5080 16652
rect 5132 16640 5138 16652
rect 5629 16643 5687 16649
rect 5629 16640 5641 16643
rect 5132 16612 5641 16640
rect 5132 16600 5138 16612
rect 5629 16609 5641 16612
rect 5675 16609 5687 16643
rect 5902 16640 5908 16652
rect 5863 16612 5908 16640
rect 5629 16603 5687 16609
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 18506 16640 18512 16652
rect 14148 16612 18512 16640
rect 14148 16600 14154 16612
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 1854 16572 1860 16584
rect 1815 16544 1860 16572
rect 1854 16532 1860 16544
rect 1912 16532 1918 16584
rect 2314 16532 2320 16584
rect 2372 16572 2378 16584
rect 2409 16575 2467 16581
rect 2409 16572 2421 16575
rect 2372 16544 2421 16572
rect 2372 16532 2378 16544
rect 2409 16541 2421 16544
rect 2455 16541 2467 16575
rect 2409 16535 2467 16541
rect 2682 16532 2688 16584
rect 2740 16532 2746 16584
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16572 18015 16575
rect 18782 16572 18788 16584
rect 18003 16544 18788 16572
rect 18003 16541 18015 16544
rect 17957 16535 18015 16541
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 57701 16575 57759 16581
rect 57701 16541 57713 16575
rect 57747 16572 57759 16575
rect 58342 16572 58348 16584
rect 57747 16544 58348 16572
rect 57747 16541 57759 16544
rect 57701 16535 57759 16541
rect 58342 16532 58348 16544
rect 58400 16532 58406 16584
rect 2700 16504 2728 16532
rect 5534 16504 5540 16516
rect 2516 16476 2728 16504
rect 5198 16476 5540 16504
rect 2516 16448 2544 16476
rect 5534 16464 5540 16476
rect 5592 16464 5598 16516
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 2498 16396 2504 16448
rect 2556 16396 2562 16448
rect 2593 16439 2651 16445
rect 2593 16405 2605 16439
rect 2639 16436 2651 16439
rect 2682 16436 2688 16448
rect 2639 16408 2688 16436
rect 2639 16405 2651 16408
rect 2593 16399 2651 16405
rect 2682 16396 2688 16408
rect 2740 16396 2746 16448
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16436 4215 16439
rect 5258 16436 5264 16448
rect 4203 16408 5264 16436
rect 4203 16405 4215 16408
rect 4157 16399 4215 16405
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 58161 16439 58219 16445
rect 58161 16405 58173 16439
rect 58207 16436 58219 16439
rect 58802 16436 58808 16448
rect 58207 16408 58808 16436
rect 58207 16405 58219 16408
rect 58161 16399 58219 16405
rect 58802 16396 58808 16408
rect 58860 16396 58866 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 2682 16192 2688 16244
rect 2740 16232 2746 16244
rect 6546 16232 6552 16244
rect 2740 16204 6552 16232
rect 2740 16192 2746 16204
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 10410 16232 10416 16244
rect 6788 16204 10272 16232
rect 10371 16204 10416 16232
rect 6788 16192 6794 16204
rect 8941 16167 8999 16173
rect 8941 16164 8953 16167
rect 6886 16136 8953 16164
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 2038 16096 2044 16108
rect 1903 16068 2044 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 4614 15988 4620 16040
rect 4672 16028 4678 16040
rect 6886 16028 6914 16136
rect 8941 16133 8953 16136
rect 8987 16133 8999 16167
rect 10244 16164 10272 16204
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 17678 16192 17684 16244
rect 17736 16232 17742 16244
rect 18141 16235 18199 16241
rect 18141 16232 18153 16235
rect 17736 16204 18153 16232
rect 17736 16192 17742 16204
rect 18141 16201 18153 16204
rect 18187 16201 18199 16235
rect 18782 16232 18788 16244
rect 18743 16204 18788 16232
rect 18141 16195 18199 16201
rect 18782 16192 18788 16204
rect 18840 16192 18846 16244
rect 16298 16164 16304 16176
rect 10244 16136 16304 16164
rect 8941 16127 8999 16133
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 19334 16164 19340 16176
rect 18340 16136 19340 16164
rect 10042 16056 10048 16108
rect 10100 16056 10106 16108
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 18340 16105 18368 16136
rect 19334 16124 19340 16136
rect 19392 16124 19398 16176
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12860 16068 13001 16096
rect 12860 16056 12866 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16065 18383 16099
rect 18325 16059 18383 16065
rect 19153 16099 19211 16105
rect 19153 16065 19165 16099
rect 19199 16096 19211 16099
rect 20162 16096 20168 16108
rect 19199 16068 20168 16096
rect 19199 16065 19211 16068
rect 19153 16059 19211 16065
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 58342 16096 58348 16108
rect 58303 16068 58348 16096
rect 58342 16056 58348 16068
rect 58400 16056 58406 16108
rect 8662 16028 8668 16040
rect 4672 16000 6914 16028
rect 8623 16000 8668 16028
rect 4672 15988 4678 16000
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 10060 16028 10088 16056
rect 9732 16000 10088 16028
rect 9732 15988 9738 16000
rect 18598 15988 18604 16040
rect 18656 16028 18662 16040
rect 19245 16031 19303 16037
rect 19245 16028 19257 16031
rect 18656 16000 19257 16028
rect 18656 15988 18662 16000
rect 19245 15997 19257 16000
rect 19291 15997 19303 16031
rect 19426 16028 19432 16040
rect 19387 16000 19432 16028
rect 19245 15991 19303 15997
rect 19426 15988 19432 16000
rect 19484 15988 19490 16040
rect 19978 15988 19984 16040
rect 20036 15988 20042 16040
rect 11514 15920 11520 15972
rect 11572 15960 11578 15972
rect 19996 15960 20024 15988
rect 11572 15932 20024 15960
rect 11572 15920 11578 15932
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 1854 15852 1860 15904
rect 1912 15892 1918 15904
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 1912 15864 2421 15892
rect 1912 15852 1918 15864
rect 2409 15861 2421 15864
rect 2455 15892 2467 15895
rect 7650 15892 7656 15904
rect 2455 15864 7656 15892
rect 2455 15861 2467 15864
rect 2409 15855 2467 15861
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 12529 15895 12587 15901
rect 12529 15892 12541 15895
rect 12492 15864 12541 15892
rect 12492 15852 12498 15864
rect 12529 15861 12541 15864
rect 12575 15892 12587 15895
rect 12802 15892 12808 15904
rect 12575 15864 12808 15892
rect 12575 15861 12587 15864
rect 12529 15855 12587 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 14458 15892 14464 15904
rect 13872 15864 14464 15892
rect 13872 15852 13878 15864
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 19426 15852 19432 15904
rect 19484 15892 19490 15904
rect 20073 15895 20131 15901
rect 20073 15892 20085 15895
rect 19484 15864 20085 15892
rect 19484 15852 19490 15864
rect 20073 15861 20085 15864
rect 20119 15892 20131 15895
rect 20346 15892 20352 15904
rect 20119 15864 20352 15892
rect 20119 15861 20131 15864
rect 20073 15855 20131 15861
rect 20346 15852 20352 15864
rect 20404 15892 20410 15904
rect 20622 15892 20628 15904
rect 20404 15864 20628 15892
rect 20404 15852 20410 15864
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 57790 15852 57796 15904
rect 57848 15892 57854 15904
rect 58161 15895 58219 15901
rect 58161 15892 58173 15895
rect 57848 15864 58173 15892
rect 57848 15852 57854 15864
rect 58161 15861 58173 15864
rect 58207 15861 58219 15895
rect 58161 15855 58219 15861
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2498 15648 2504 15700
rect 2556 15688 2562 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 2556 15660 2789 15688
rect 2556 15648 2562 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 2777 15651 2835 15657
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 5905 15691 5963 15697
rect 5905 15688 5917 15691
rect 5684 15660 5917 15688
rect 5684 15648 5690 15660
rect 5905 15657 5917 15660
rect 5951 15657 5963 15691
rect 8018 15688 8024 15700
rect 5905 15651 5963 15657
rect 6012 15660 8024 15688
rect 2038 15620 2044 15632
rect 1951 15592 2044 15620
rect 2038 15580 2044 15592
rect 2096 15620 2102 15632
rect 6012 15620 6040 15660
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 8386 15648 8392 15700
rect 8444 15688 8450 15700
rect 10873 15691 10931 15697
rect 10873 15688 10885 15691
rect 8444 15660 10885 15688
rect 8444 15648 8450 15660
rect 10873 15657 10885 15660
rect 10919 15657 10931 15691
rect 18598 15688 18604 15700
rect 18559 15660 18604 15688
rect 10873 15651 10931 15657
rect 18598 15648 18604 15660
rect 18656 15648 18662 15700
rect 58342 15688 58348 15700
rect 58303 15660 58348 15688
rect 58342 15648 58348 15660
rect 58400 15648 58406 15700
rect 2096 15592 6040 15620
rect 2096 15580 2102 15592
rect 3050 15512 3056 15564
rect 3108 15552 3114 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 3108 15524 7389 15552
rect 3108 15512 3114 15524
rect 7377 15521 7389 15524
rect 7423 15521 7435 15555
rect 9398 15552 9404 15564
rect 9359 15524 9404 15552
rect 7377 15515 7435 15521
rect 9398 15512 9404 15524
rect 9456 15512 9462 15564
rect 57238 15552 57244 15564
rect 57199 15524 57244 15552
rect 57238 15512 57244 15524
rect 57296 15512 57302 15564
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15484 7711 15487
rect 8294 15484 8300 15496
rect 7699 15456 8300 15484
rect 7699 15453 7711 15456
rect 7653 15447 7711 15453
rect 8294 15444 8300 15456
rect 8352 15484 8358 15496
rect 8662 15484 8668 15496
rect 8352 15456 8668 15484
rect 8352 15444 8358 15456
rect 8662 15444 8668 15456
rect 8720 15484 8726 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8720 15456 9137 15484
rect 8720 15444 8726 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 19484 15456 19625 15484
rect 19484 15444 19490 15456
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 56965 15487 57023 15493
rect 56965 15484 56977 15487
rect 19613 15447 19671 15453
rect 56428 15456 56977 15484
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 5592 15388 6210 15416
rect 5592 15376 5598 15388
rect 10042 15376 10048 15428
rect 10100 15376 10106 15428
rect 56428 15360 56456 15456
rect 56965 15453 56977 15456
rect 57011 15453 57023 15487
rect 56965 15447 57023 15453
rect 4890 15308 4896 15360
rect 4948 15348 4954 15360
rect 7282 15348 7288 15360
rect 4948 15320 7288 15348
rect 4948 15308 4954 15320
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 12342 15348 12348 15360
rect 7616 15320 12348 15348
rect 7616 15308 7622 15320
rect 12342 15308 12348 15320
rect 12400 15308 12406 15360
rect 18690 15308 18696 15360
rect 18748 15348 18754 15360
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 18748 15320 19441 15348
rect 18748 15308 18754 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 20070 15348 20076 15360
rect 20031 15320 20076 15348
rect 19429 15311 19487 15317
rect 20070 15308 20076 15320
rect 20128 15308 20134 15360
rect 56410 15348 56416 15360
rect 56371 15320 56416 15348
rect 56410 15308 56416 15320
rect 56468 15308 56474 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 12342 15144 12348 15156
rect 12303 15116 12348 15144
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 18690 15144 18696 15156
rect 13872 15116 18696 15144
rect 13872 15104 13878 15116
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19613 15147 19671 15153
rect 19613 15144 19625 15147
rect 19484 15116 19625 15144
rect 19484 15104 19490 15116
rect 19613 15113 19625 15116
rect 19659 15113 19671 15147
rect 19613 15107 19671 15113
rect 2130 15076 2136 15088
rect 2043 15048 2136 15076
rect 2056 14949 2084 15048
rect 2130 15036 2136 15048
rect 2188 15076 2194 15088
rect 2498 15076 2504 15088
rect 2188 15048 2504 15076
rect 2188 15036 2194 15048
rect 2498 15036 2504 15048
rect 2556 15036 2562 15088
rect 14829 15079 14887 15085
rect 14829 15076 14841 15079
rect 13386 15048 14841 15076
rect 14829 15045 14841 15048
rect 14875 15076 14887 15079
rect 15010 15076 15016 15088
rect 14875 15048 15016 15076
rect 14875 15045 14887 15048
rect 14829 15039 14887 15045
rect 15010 15036 15016 15048
rect 15068 15076 15074 15088
rect 19886 15076 19892 15088
rect 15068 15048 17618 15076
rect 18616 15048 19892 15076
rect 15068 15036 15074 15048
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 3142 15008 3148 15020
rect 2363 14980 3148 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 9631 14980 10180 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 2280 14912 2325 14940
rect 2280 14900 2286 14912
rect 10152 14881 10180 14980
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 14424 14980 14565 15008
rect 14424 14968 14430 14980
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 14553 14971 14611 14977
rect 14660 14980 16865 15008
rect 13814 14940 13820 14952
rect 13775 14912 13820 14940
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14458 14940 14464 14952
rect 14139 14912 14464 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14458 14900 14464 14912
rect 14516 14940 14522 14952
rect 14660 14940 14688 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 14516 14912 14688 14940
rect 17129 14943 17187 14949
rect 14516 14900 14522 14912
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 18616 14940 18644 15048
rect 19886 15036 19892 15048
rect 19944 15036 19950 15088
rect 19981 15079 20039 15085
rect 19981 15045 19993 15079
rect 20027 15076 20039 15079
rect 20162 15076 20168 15088
rect 20027 15048 20168 15076
rect 20027 15045 20039 15048
rect 19981 15039 20039 15045
rect 20162 15036 20168 15048
rect 20220 15036 20226 15088
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 17175 14912 18644 14940
rect 18708 14980 18889 15008
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 10137 14875 10195 14881
rect 10137 14841 10149 14875
rect 10183 14872 10195 14875
rect 12802 14872 12808 14884
rect 10183 14844 12808 14872
rect 10183 14841 10195 14844
rect 10137 14835 10195 14841
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 2682 14804 2688 14816
rect 2643 14776 2688 14804
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 3142 14804 3148 14816
rect 3103 14776 3148 14804
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 3786 14804 3792 14816
rect 3699 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14804 3850 14816
rect 5258 14804 5264 14816
rect 3844 14776 5264 14804
rect 3844 14764 3850 14776
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 8294 14804 8300 14816
rect 8255 14776 8300 14804
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 17494 14764 17500 14816
rect 17552 14804 17558 14816
rect 18708 14804 18736 14980
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 57517 15011 57575 15017
rect 57517 14977 57529 15011
rect 57563 15008 57575 15011
rect 58342 15008 58348 15020
rect 57563 14980 58348 15008
rect 57563 14977 57575 14980
rect 57517 14971 57575 14977
rect 58342 14968 58348 14980
rect 58400 14968 58406 15020
rect 20070 14940 20076 14952
rect 20031 14912 20076 14940
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 20257 14943 20315 14949
rect 20257 14909 20269 14943
rect 20303 14940 20315 14943
rect 20622 14940 20628 14952
rect 20303 14912 20628 14940
rect 20303 14909 20315 14912
rect 20257 14903 20315 14909
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 17552 14776 18736 14804
rect 17552 14764 17558 14776
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 20622 14804 20628 14816
rect 20036 14776 20628 14804
rect 20036 14764 20042 14776
rect 20622 14764 20628 14776
rect 20680 14804 20686 14816
rect 20809 14807 20867 14813
rect 20809 14804 20821 14807
rect 20680 14776 20821 14804
rect 20680 14764 20686 14776
rect 20809 14773 20821 14776
rect 20855 14773 20867 14807
rect 20809 14767 20867 14773
rect 57330 14764 57336 14816
rect 57388 14804 57394 14816
rect 58161 14807 58219 14813
rect 58161 14804 58173 14807
rect 57388 14776 58173 14804
rect 57388 14764 57394 14776
rect 58161 14773 58173 14776
rect 58207 14773 58219 14807
rect 58161 14767 58219 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 3786 14600 3792 14612
rect 1872 14572 3792 14600
rect 1872 14405 1900 14572
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 5077 14603 5135 14609
rect 5077 14569 5089 14603
rect 5123 14600 5135 14603
rect 5166 14600 5172 14612
rect 5123 14572 5172 14600
rect 5123 14569 5135 14572
rect 5077 14563 5135 14569
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 13262 14600 13268 14612
rect 5316 14572 13268 14600
rect 5316 14560 5322 14572
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 18785 14603 18843 14609
rect 18785 14600 18797 14603
rect 18564 14572 18797 14600
rect 18564 14560 18570 14572
rect 18785 14569 18797 14572
rect 18831 14569 18843 14603
rect 18785 14563 18843 14569
rect 2590 14492 2596 14544
rect 2648 14532 2654 14544
rect 3237 14535 3295 14541
rect 2648 14504 3096 14532
rect 2648 14492 2654 14504
rect 3068 14405 3096 14504
rect 3237 14501 3249 14535
rect 3283 14532 3295 14535
rect 4614 14532 4620 14544
rect 3283 14504 4620 14532
rect 3283 14501 3295 14504
rect 3237 14495 3295 14501
rect 4614 14492 4620 14504
rect 4672 14492 4678 14544
rect 6546 14464 6552 14476
rect 6507 14436 6552 14464
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14464 6883 14467
rect 8294 14464 8300 14476
rect 6871 14436 8300 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 8294 14424 8300 14436
rect 8352 14464 8358 14476
rect 9309 14467 9367 14473
rect 9309 14464 9321 14467
rect 8352 14436 9321 14464
rect 8352 14424 8358 14436
rect 9309 14433 9321 14436
rect 9355 14433 9367 14467
rect 18800 14464 18828 14563
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19429 14603 19487 14609
rect 19429 14600 19441 14603
rect 19392 14572 19441 14600
rect 19392 14560 19398 14572
rect 19429 14569 19441 14572
rect 19475 14569 19487 14603
rect 19429 14563 19487 14569
rect 19886 14560 19892 14612
rect 19944 14600 19950 14612
rect 20809 14603 20867 14609
rect 20809 14600 20821 14603
rect 19944 14572 20821 14600
rect 19944 14560 19950 14572
rect 20809 14569 20821 14572
rect 20855 14569 20867 14603
rect 20809 14563 20867 14569
rect 19889 14467 19947 14473
rect 19889 14464 19901 14467
rect 18800 14436 19901 14464
rect 9309 14427 9367 14433
rect 19889 14433 19901 14436
rect 19935 14433 19947 14467
rect 19889 14427 19947 14433
rect 19978 14424 19984 14476
rect 20036 14464 20042 14476
rect 20530 14464 20536 14476
rect 20036 14436 20536 14464
rect 20036 14424 20042 14436
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14365 1915 14399
rect 1857 14359 1915 14365
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14365 3111 14399
rect 3053 14359 3111 14365
rect 2608 14328 2636 14359
rect 12342 14356 12348 14408
rect 12400 14396 12406 14408
rect 20070 14396 20076 14408
rect 12400 14368 20076 14396
rect 12400 14356 12406 14368
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 20993 14399 21051 14405
rect 20993 14396 21005 14399
rect 20772 14368 21005 14396
rect 20772 14356 20778 14368
rect 20993 14365 21005 14368
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 57701 14399 57759 14405
rect 57701 14365 57713 14399
rect 57747 14396 57759 14399
rect 58342 14396 58348 14408
rect 57747 14368 58348 14396
rect 57747 14365 57759 14368
rect 57701 14359 57759 14365
rect 58342 14356 58348 14368
rect 58400 14356 58406 14408
rect 2608 14300 4108 14328
rect 2406 14260 2412 14272
rect 2367 14232 2412 14260
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 4080 14269 4108 14300
rect 5166 14288 5172 14340
rect 5224 14328 5230 14340
rect 9582 14328 9588 14340
rect 5224 14300 5382 14328
rect 9543 14300 9588 14328
rect 5224 14288 5230 14300
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 11517 14331 11575 14337
rect 10810 14300 11468 14328
rect 4065 14263 4123 14269
rect 4065 14229 4077 14263
rect 4111 14260 4123 14263
rect 8938 14260 8944 14272
rect 4111 14232 8944 14260
rect 4111 14229 4123 14232
rect 4065 14223 4123 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 11054 14260 11060 14272
rect 11015 14232 11060 14260
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 11440 14260 11468 14300
rect 11517 14297 11529 14331
rect 11563 14328 11575 14331
rect 11606 14328 11612 14340
rect 11563 14300 11612 14328
rect 11563 14297 11575 14300
rect 11517 14291 11575 14297
rect 11606 14288 11612 14300
rect 11664 14288 11670 14340
rect 12618 14260 12624 14272
rect 11440 14232 12624 14260
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 12802 14260 12808 14272
rect 12763 14232 12808 14260
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 19797 14263 19855 14269
rect 19797 14229 19809 14263
rect 19843 14260 19855 14263
rect 20070 14260 20076 14272
rect 19843 14232 20076 14260
rect 19843 14229 19855 14232
rect 19797 14223 19855 14229
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 58158 14260 58164 14272
rect 58119 14232 58164 14260
rect 58158 14220 58164 14232
rect 58216 14220 58222 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 3329 14059 3387 14065
rect 3329 14025 3341 14059
rect 3375 14056 3387 14059
rect 5258 14056 5264 14068
rect 3375 14028 5264 14056
rect 3375 14025 3387 14028
rect 3329 14019 3387 14025
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 13265 14059 13323 14065
rect 13265 14025 13277 14059
rect 13311 14056 13323 14059
rect 16666 14056 16672 14068
rect 13311 14028 16672 14056
rect 13311 14025 13323 14028
rect 13265 14019 13323 14025
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 17552 14028 20177 14056
rect 17552 14016 17558 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 20714 14056 20720 14068
rect 20675 14028 20720 14056
rect 20165 14019 20223 14025
rect 2317 13991 2375 13997
rect 2317 13957 2329 13991
rect 2363 13988 2375 13991
rect 2774 13988 2780 14000
rect 2363 13960 2780 13988
rect 2363 13957 2375 13960
rect 2317 13951 2375 13957
rect 2774 13948 2780 13960
rect 2832 13988 2838 14000
rect 3878 13988 3884 14000
rect 2832 13960 3884 13988
rect 2832 13948 2838 13960
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 12618 13948 12624 14000
rect 12676 13988 12682 14000
rect 20180 13988 20208 14019
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 57238 14016 57244 14068
rect 57296 14056 57302 14068
rect 57698 14056 57704 14068
rect 57296 14028 57704 14056
rect 57296 14016 57302 14028
rect 57698 14016 57704 14028
rect 57756 14056 57762 14068
rect 58253 14059 58311 14065
rect 58253 14056 58265 14059
rect 57756 14028 58265 14056
rect 57756 14016 57762 14028
rect 58253 14025 58265 14028
rect 58299 14025 58311 14059
rect 58253 14019 58311 14025
rect 58434 14016 58440 14068
rect 58492 14056 58498 14068
rect 58986 14056 58992 14068
rect 58492 14028 58992 14056
rect 58492 14016 58498 14028
rect 58986 14016 58992 14028
rect 59044 14016 59050 14068
rect 21177 13991 21235 13997
rect 21177 13988 21189 13991
rect 12676 13960 13570 13988
rect 20180 13960 21189 13988
rect 12676 13948 12682 13960
rect 21177 13957 21189 13960
rect 21223 13957 21235 13991
rect 21177 13951 21235 13957
rect 2038 13880 2044 13932
rect 2096 13920 2102 13932
rect 2096 13892 2268 13920
rect 2096 13880 2102 13892
rect 2130 13852 2136 13864
rect 2091 13824 2136 13852
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 2240 13861 2268 13892
rect 2682 13880 2688 13932
rect 2740 13920 2746 13932
rect 3145 13923 3203 13929
rect 3145 13920 3157 13923
rect 2740 13892 3157 13920
rect 2740 13880 2746 13892
rect 3145 13889 3157 13892
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 20070 13880 20076 13932
rect 20128 13920 20134 13932
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 20128 13892 21097 13920
rect 20128 13880 20134 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 11054 13852 11060 13864
rect 2271 13824 11060 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11664 13824 11713 13852
rect 11664 13812 11670 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 15010 13852 15016 13864
rect 14971 13824 15016 13852
rect 11701 13815 11759 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 20346 13812 20352 13864
rect 20404 13852 20410 13864
rect 20404 13824 20760 13852
rect 20404 13812 20410 13824
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 2685 13719 2743 13725
rect 2685 13716 2697 13719
rect 2372 13688 2697 13716
rect 2372 13676 2378 13688
rect 2685 13685 2697 13688
rect 2731 13685 2743 13719
rect 2685 13679 2743 13685
rect 14755 13719 14813 13725
rect 14755 13685 14767 13719
rect 14801 13716 14813 13719
rect 15746 13716 15752 13728
rect 14801 13688 15752 13716
rect 14801 13685 14813 13688
rect 14755 13679 14813 13685
rect 15746 13676 15752 13688
rect 15804 13676 15810 13728
rect 20732 13716 20760 13824
rect 21100 13784 21128 13883
rect 21361 13855 21419 13861
rect 21361 13821 21373 13855
rect 21407 13852 21419 13855
rect 22094 13852 22100 13864
rect 21407 13824 22100 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 22646 13784 22652 13796
rect 21100 13756 22652 13784
rect 22646 13744 22652 13756
rect 22704 13744 22710 13796
rect 22005 13719 22063 13725
rect 22005 13716 22017 13719
rect 20732 13688 22017 13716
rect 22005 13685 22017 13688
rect 22051 13716 22063 13719
rect 22094 13716 22100 13728
rect 22051 13688 22100 13716
rect 22051 13685 22063 13688
rect 22005 13679 22063 13685
rect 22094 13676 22100 13688
rect 22152 13676 22158 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 2501 13515 2559 13521
rect 2501 13481 2513 13515
rect 2547 13512 2559 13515
rect 9582 13512 9588 13524
rect 2547 13484 9588 13512
rect 2547 13481 2559 13484
rect 2501 13475 2559 13481
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 18417 13515 18475 13521
rect 18417 13512 18429 13515
rect 15988 13484 18429 13512
rect 15988 13472 15994 13484
rect 18417 13481 18429 13484
rect 18463 13512 18475 13515
rect 19426 13512 19432 13524
rect 18463 13484 19432 13512
rect 18463 13481 18475 13484
rect 18417 13475 18475 13481
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 2130 13404 2136 13456
rect 2188 13444 2194 13456
rect 2961 13447 3019 13453
rect 2961 13444 2973 13447
rect 2188 13416 2973 13444
rect 2188 13404 2194 13416
rect 2961 13413 2973 13416
rect 3007 13413 3019 13447
rect 58618 13444 58624 13456
rect 2961 13407 3019 13413
rect 57624 13416 58624 13444
rect 57146 13376 57152 13388
rect 57107 13348 57152 13376
rect 57146 13336 57152 13348
rect 57204 13336 57210 13388
rect 57330 13385 57336 13388
rect 57308 13379 57336 13385
rect 57308 13345 57320 13379
rect 57308 13339 57336 13345
rect 57330 13336 57336 13339
rect 57388 13336 57394 13388
rect 57425 13379 57483 13385
rect 57425 13345 57437 13379
rect 57471 13376 57483 13379
rect 57624 13376 57652 13416
rect 58618 13404 58624 13416
rect 58676 13404 58682 13456
rect 57471 13348 57652 13376
rect 57471 13345 57483 13348
rect 57425 13339 57483 13345
rect 57698 13336 57704 13388
rect 57756 13376 57762 13388
rect 58161 13379 58219 13385
rect 57756 13348 57801 13376
rect 57756 13336 57762 13348
rect 58161 13345 58173 13379
rect 58207 13376 58219 13379
rect 58710 13376 58716 13388
rect 58207 13348 58716 13376
rect 58207 13345 58219 13348
rect 58161 13339 58219 13345
rect 58710 13336 58716 13348
rect 58768 13336 58774 13388
rect 1854 13308 1860 13320
rect 1815 13280 1860 13308
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 16666 13308 16672 13320
rect 16627 13280 16672 13308
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 58250 13268 58256 13320
rect 58308 13308 58314 13320
rect 58345 13311 58403 13317
rect 58345 13308 58357 13311
rect 58308 13280 58357 13308
rect 58308 13268 58314 13280
rect 58345 13277 58357 13280
rect 58391 13277 58403 13311
rect 58345 13271 58403 13277
rect 16942 13240 16948 13252
rect 16903 13212 16948 13240
rect 16942 13200 16948 13212
rect 17000 13200 17006 13252
rect 17052 13212 17434 13240
rect 1670 13172 1676 13184
rect 1631 13144 1676 13172
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 16022 13132 16028 13184
rect 16080 13172 16086 13184
rect 17052 13172 17080 13212
rect 16080 13144 17080 13172
rect 16080 13132 16086 13144
rect 55674 13132 55680 13184
rect 55732 13172 55738 13184
rect 56505 13175 56563 13181
rect 56505 13172 56517 13175
rect 55732 13144 56517 13172
rect 55732 13132 55738 13144
rect 56505 13141 56517 13144
rect 56551 13141 56563 13175
rect 56505 13135 56563 13141
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 17000 12940 18429 12968
rect 17000 12928 17006 12940
rect 18417 12937 18429 12940
rect 18463 12937 18475 12971
rect 18417 12931 18475 12937
rect 19061 12971 19119 12977
rect 19061 12937 19073 12971
rect 19107 12937 19119 12971
rect 19061 12931 19119 12937
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 1946 12832 1952 12844
rect 1903 12804 1952 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12832 18659 12835
rect 19076 12832 19104 12931
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 19521 12971 19579 12977
rect 19521 12968 19533 12971
rect 19484 12940 19533 12968
rect 19484 12928 19490 12940
rect 19521 12937 19533 12940
rect 19567 12937 19579 12971
rect 19521 12931 19579 12937
rect 57146 12928 57152 12980
rect 57204 12968 57210 12980
rect 57425 12971 57483 12977
rect 57425 12968 57437 12971
rect 57204 12940 57437 12968
rect 57204 12928 57210 12940
rect 57425 12937 57437 12940
rect 57471 12937 57483 12971
rect 57425 12931 57483 12937
rect 18647 12804 19104 12832
rect 19429 12835 19487 12841
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 19429 12801 19441 12835
rect 19475 12832 19487 12835
rect 20070 12832 20076 12844
rect 19475 12804 20076 12832
rect 19475 12801 19487 12804
rect 19429 12795 19487 12801
rect 20070 12792 20076 12804
rect 20128 12792 20134 12844
rect 57882 12792 57888 12844
rect 57940 12832 57946 12844
rect 58345 12835 58403 12841
rect 58345 12832 58357 12835
rect 57940 12804 58357 12832
rect 57940 12792 57946 12804
rect 58345 12801 58357 12804
rect 58391 12801 58403 12835
rect 58345 12795 58403 12801
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12764 19763 12767
rect 20622 12764 20628 12776
rect 19751 12736 20628 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 1854 12656 1860 12708
rect 1912 12696 1918 12708
rect 2409 12699 2467 12705
rect 2409 12696 2421 12699
rect 1912 12668 2421 12696
rect 1912 12656 1918 12668
rect 2409 12665 2421 12668
rect 2455 12696 2467 12699
rect 10870 12696 10876 12708
rect 2455 12668 10876 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 20364 12640 20392 12736
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 57330 12656 57336 12708
rect 57388 12696 57394 12708
rect 58161 12699 58219 12705
rect 58161 12696 58173 12699
rect 57388 12668 58173 12696
rect 57388 12656 57394 12668
rect 58161 12665 58173 12668
rect 58207 12665 58219 12699
rect 58161 12659 58219 12665
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 20346 12628 20352 12640
rect 20307 12600 20352 12628
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 9214 12424 9220 12436
rect 5040 12396 6914 12424
rect 9175 12396 9220 12424
rect 5040 12384 5046 12396
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 6886 12084 6914 12396
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 19426 12424 19432 12436
rect 19387 12396 19432 12424
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 57701 12427 57759 12433
rect 57701 12393 57713 12427
rect 57747 12424 57759 12427
rect 57882 12424 57888 12436
rect 57747 12396 57888 12424
rect 57747 12393 57759 12396
rect 57701 12387 57759 12393
rect 57882 12384 57888 12396
rect 57940 12384 57946 12436
rect 15838 12356 15844 12368
rect 15799 12328 15844 12356
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 9364 12260 10977 12288
rect 9364 12248 9370 12260
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 16724 12260 17601 12288
rect 16724 12248 16730 12260
rect 17589 12257 17601 12260
rect 17635 12257 17647 12291
rect 17589 12251 17647 12257
rect 58066 12248 58072 12300
rect 58124 12288 58130 12300
rect 58618 12288 58624 12300
rect 58124 12260 58624 12288
rect 58124 12248 58130 12260
rect 58618 12248 58624 12260
rect 58676 12248 58682 12300
rect 55674 12220 55680 12232
rect 55635 12192 55680 12220
rect 55674 12180 55680 12192
rect 55732 12180 55738 12232
rect 57149 12223 57207 12229
rect 57149 12189 57161 12223
rect 57195 12220 57207 12223
rect 58342 12220 58348 12232
rect 57195 12192 58348 12220
rect 57195 12189 57207 12192
rect 57149 12183 57207 12189
rect 58342 12180 58348 12192
rect 58400 12180 58406 12232
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 10689 12155 10747 12161
rect 9456 12124 9522 12152
rect 9456 12112 9462 12124
rect 10689 12121 10701 12155
rect 10735 12121 10747 12155
rect 10689 12115 10747 12121
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 6886 12056 8585 12084
rect 8573 12053 8585 12056
rect 8619 12084 8631 12087
rect 10704 12084 10732 12115
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 13170 12152 13176 12164
rect 12676 12124 13176 12152
rect 12676 12112 12682 12124
rect 13170 12112 13176 12124
rect 13228 12152 13234 12164
rect 13722 12152 13728 12164
rect 13228 12124 13728 12152
rect 13228 12112 13234 12124
rect 13722 12112 13728 12124
rect 13780 12152 13786 12164
rect 16022 12152 16028 12164
rect 13780 12124 16028 12152
rect 13780 12112 13786 12124
rect 16022 12112 16028 12124
rect 16080 12152 16086 12164
rect 17313 12155 17371 12161
rect 16080 12124 16146 12152
rect 16080 12112 16086 12124
rect 17313 12121 17325 12155
rect 17359 12152 17371 12155
rect 18690 12152 18696 12164
rect 17359 12124 18696 12152
rect 17359 12121 17371 12124
rect 17313 12115 17371 12121
rect 18690 12112 18696 12124
rect 18748 12112 18754 12164
rect 8619 12056 10732 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 42978 12044 42984 12096
rect 43036 12084 43042 12096
rect 55493 12087 55551 12093
rect 55493 12084 55505 12087
rect 43036 12056 55505 12084
rect 43036 12044 43042 12056
rect 55493 12053 55505 12056
rect 55539 12053 55551 12087
rect 55493 12047 55551 12053
rect 58066 12044 58072 12096
rect 58124 12084 58130 12096
rect 58161 12087 58219 12093
rect 58161 12084 58173 12087
rect 58124 12056 58173 12084
rect 58124 12044 58130 12056
rect 58161 12053 58173 12056
rect 58207 12053 58219 12087
rect 58161 12047 58219 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 11057 11883 11115 11889
rect 5224 11852 6914 11880
rect 5224 11840 5230 11852
rect 2498 11772 2504 11824
rect 2556 11812 2562 11824
rect 3053 11815 3111 11821
rect 3053 11812 3065 11815
rect 2556 11784 3065 11812
rect 2556 11772 2562 11784
rect 3053 11781 3065 11784
rect 3099 11812 3111 11815
rect 6270 11812 6276 11824
rect 3099 11784 6276 11812
rect 3099 11781 3111 11784
rect 3053 11775 3111 11781
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 6886 11812 6914 11852
rect 11057 11849 11069 11883
rect 11103 11880 11115 11883
rect 11330 11880 11336 11892
rect 11103 11852 11336 11880
rect 11103 11849 11115 11852
rect 11057 11843 11115 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 19061 11883 19119 11889
rect 19061 11880 19073 11883
rect 13832 11852 19073 11880
rect 13722 11812 13728 11824
rect 6886 11784 10074 11812
rect 13386 11784 13728 11812
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 13832 11821 13860 11852
rect 19061 11849 19073 11852
rect 19107 11849 19119 11883
rect 19061 11843 19119 11849
rect 13817 11815 13875 11821
rect 13817 11781 13829 11815
rect 13863 11781 13875 11815
rect 13817 11775 13875 11781
rect 15838 11772 15844 11824
rect 15896 11812 15902 11824
rect 19705 11815 19763 11821
rect 19705 11812 19717 11815
rect 15896 11784 19717 11812
rect 15896 11772 15902 11784
rect 19705 11781 19717 11784
rect 19751 11812 19763 11815
rect 19886 11812 19892 11824
rect 19751 11784 19892 11812
rect 19751 11781 19763 11784
rect 19705 11775 19763 11781
rect 19886 11772 19892 11784
rect 19944 11772 19950 11824
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 9306 11744 9312 11756
rect 1903 11716 2452 11744
rect 9267 11716 9312 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 1670 11608 1676 11620
rect 1631 11580 1676 11608
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 2424 11552 2452 11716
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 19245 11747 19303 11753
rect 19245 11713 19257 11747
rect 19291 11744 19303 11747
rect 19426 11744 19432 11756
rect 19291 11716 19432 11744
rect 19291 11713 19303 11716
rect 19245 11707 19303 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 57517 11747 57575 11753
rect 57517 11713 57529 11747
rect 57563 11744 57575 11747
rect 58342 11744 58348 11756
rect 57563 11716 58348 11744
rect 57563 11713 57575 11716
rect 57517 11707 57575 11713
rect 58342 11704 58348 11716
rect 58400 11704 58406 11756
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9180 11648 9597 11676
rect 9180 11636 9186 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11676 14151 11679
rect 14458 11676 14464 11688
rect 14139 11648 14464 11676
rect 14139 11645 14151 11648
rect 14093 11639 14151 11645
rect 14458 11636 14464 11648
rect 14516 11676 14522 11688
rect 15010 11676 15016 11688
rect 14516 11648 15016 11676
rect 14516 11636 14522 11648
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 2682 11568 2688 11620
rect 2740 11608 2746 11620
rect 3513 11611 3571 11617
rect 3513 11608 3525 11611
rect 2740 11580 3525 11608
rect 2740 11568 2746 11580
rect 3513 11577 3525 11580
rect 3559 11577 3571 11611
rect 3513 11571 3571 11577
rect 57238 11568 57244 11620
rect 57296 11608 57302 11620
rect 57422 11608 57428 11620
rect 57296 11580 57428 11608
rect 57296 11568 57302 11580
rect 57422 11568 57428 11580
rect 57480 11568 57486 11620
rect 2406 11540 2412 11552
rect 2367 11512 2412 11540
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 6822 11540 6828 11552
rect 4856 11512 6828 11540
rect 4856 11500 4862 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 12342 11540 12348 11552
rect 12303 11512 12348 11540
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 20714 11540 20720 11552
rect 20675 11512 20720 11540
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 56686 11500 56692 11552
rect 56744 11540 56750 11552
rect 58161 11543 58219 11549
rect 58161 11540 58173 11543
rect 56744 11512 58173 11540
rect 56744 11500 56750 11512
rect 58161 11509 58173 11512
rect 58207 11509 58219 11543
rect 58161 11503 58219 11509
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 12342 11336 12348 11348
rect 2464 11308 12348 11336
rect 2464 11296 2470 11308
rect 12342 11296 12348 11308
rect 12400 11336 12406 11348
rect 18506 11336 18512 11348
rect 12400 11308 18512 11336
rect 12400 11296 12406 11308
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 56505 11339 56563 11345
rect 56505 11305 56517 11339
rect 56551 11336 56563 11339
rect 57146 11336 57152 11348
rect 56551 11308 57152 11336
rect 56551 11305 56563 11308
rect 56505 11299 56563 11305
rect 57146 11296 57152 11308
rect 57204 11296 57210 11348
rect 57422 11296 57428 11348
rect 57480 11336 57486 11348
rect 58986 11336 58992 11348
rect 57480 11308 58992 11336
rect 57480 11296 57486 11308
rect 58986 11296 58992 11308
rect 59044 11296 59050 11348
rect 2685 11271 2743 11277
rect 2685 11237 2697 11271
rect 2731 11237 2743 11271
rect 2685 11231 2743 11237
rect 3329 11271 3387 11277
rect 3329 11237 3341 11271
rect 3375 11237 3387 11271
rect 6730 11268 6736 11280
rect 6691 11240 6736 11268
rect 3329 11231 3387 11237
rect 2130 11200 2136 11212
rect 2091 11172 2136 11200
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2498 11132 2504 11144
rect 2363 11104 2504 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 2700 11132 2728 11231
rect 3344 11200 3372 11231
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 19429 11271 19487 11277
rect 19429 11237 19441 11271
rect 19475 11237 19487 11271
rect 58158 11268 58164 11280
rect 19429 11231 19487 11237
rect 57624 11240 58164 11268
rect 5810 11200 5816 11212
rect 3344 11172 5816 11200
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11200 5963 11203
rect 6748 11200 6776 11228
rect 5951 11172 6776 11200
rect 5951 11169 5963 11172
rect 5905 11163 5963 11169
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 16206 11200 16212 11212
rect 6880 11172 16212 11200
rect 6880 11160 6886 11172
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 3145 11135 3203 11141
rect 3145 11132 3157 11135
rect 2700 11104 3157 11132
rect 3145 11101 3157 11104
rect 3191 11101 3203 11135
rect 3145 11095 3203 11101
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4614 11132 4620 11144
rect 4203 11104 4620 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11132 18935 11135
rect 19444 11132 19472 11231
rect 19886 11200 19892 11212
rect 19847 11172 19892 11200
rect 19886 11160 19892 11172
rect 19944 11160 19950 11212
rect 19978 11160 19984 11212
rect 20036 11200 20042 11212
rect 20073 11203 20131 11209
rect 20073 11200 20085 11203
rect 20036 11172 20085 11200
rect 20036 11160 20042 11172
rect 20073 11169 20085 11172
rect 20119 11200 20131 11203
rect 21082 11200 21088 11212
rect 20119 11172 21088 11200
rect 20119 11169 20131 11172
rect 20073 11163 20131 11169
rect 21082 11160 21088 11172
rect 21140 11160 21146 11212
rect 21545 11203 21603 11209
rect 21545 11169 21557 11203
rect 21591 11169 21603 11203
rect 21545 11163 21603 11169
rect 18923 11104 19472 11132
rect 19797 11135 19855 11141
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 20162 11132 20168 11144
rect 19843 11104 20168 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 2222 11064 2228 11076
rect 2183 11036 2228 11064
rect 2222 11024 2228 11036
rect 2280 11024 2286 11076
rect 5166 11024 5172 11076
rect 5224 11024 5230 11076
rect 5994 11024 6000 11076
rect 6052 11064 6058 11076
rect 6196 11064 6224 11095
rect 20162 11092 20168 11104
rect 20220 11132 20226 11144
rect 20622 11132 20628 11144
rect 20220 11104 20628 11132
rect 20220 11092 20226 11104
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 20772 11104 21373 11132
rect 20772 11092 20778 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 6052 11036 6224 11064
rect 6052 11024 6058 11036
rect 20806 11024 20812 11076
rect 20864 11064 20870 11076
rect 21269 11067 21327 11073
rect 21269 11064 21281 11067
rect 20864 11036 21281 11064
rect 20864 11024 20870 11036
rect 21269 11033 21281 11036
rect 21315 11033 21327 11067
rect 21560 11064 21588 11163
rect 56962 11160 56968 11212
rect 57020 11200 57026 11212
rect 57149 11203 57207 11209
rect 57149 11200 57161 11203
rect 57020 11172 57161 11200
rect 57020 11160 57026 11172
rect 57149 11169 57161 11172
rect 57195 11169 57207 11203
rect 57149 11163 57207 11169
rect 57308 11203 57366 11209
rect 57308 11169 57320 11203
rect 57354 11200 57366 11203
rect 57624 11200 57652 11240
rect 58158 11228 58164 11240
rect 58216 11228 58222 11280
rect 57354 11172 57652 11200
rect 57354 11169 57366 11172
rect 57308 11163 57366 11169
rect 57698 11160 57704 11212
rect 57756 11200 57762 11212
rect 57756 11172 57801 11200
rect 57756 11160 57762 11172
rect 57422 11132 57428 11144
rect 57383 11104 57428 11132
rect 57422 11092 57428 11104
rect 57480 11092 57486 11144
rect 57974 11092 57980 11144
rect 58032 11132 58038 11144
rect 58161 11135 58219 11141
rect 58161 11132 58173 11135
rect 58032 11104 58173 11132
rect 58032 11092 58038 11104
rect 58161 11101 58173 11104
rect 58207 11101 58219 11135
rect 58342 11132 58348 11144
rect 58303 11104 58348 11132
rect 58161 11095 58219 11101
rect 58342 11092 58348 11104
rect 58400 11092 58406 11144
rect 22094 11064 22100 11076
rect 21560 11036 22100 11064
rect 21269 11027 21327 11033
rect 22094 11024 22100 11036
rect 22152 11064 22158 11076
rect 22189 11067 22247 11073
rect 22189 11064 22201 11067
rect 22152 11036 22201 11064
rect 22152 11024 22158 11036
rect 22189 11033 22201 11036
rect 22235 11064 22247 11067
rect 22554 11064 22560 11076
rect 22235 11036 22560 11064
rect 22235 11033 22247 11036
rect 22189 11027 22247 11033
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 20714 10996 20720 11008
rect 13596 10968 20720 10996
rect 13596 10956 13602 10968
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 20898 10996 20904 11008
rect 20859 10968 20904 10996
rect 20898 10956 20904 10968
rect 20956 10956 20962 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 2685 10795 2743 10801
rect 2685 10761 2697 10795
rect 2731 10761 2743 10795
rect 2685 10755 2743 10761
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2700 10656 2728 10755
rect 14458 10752 14464 10804
rect 14516 10792 14522 10804
rect 16666 10792 16672 10804
rect 14516 10764 16672 10792
rect 14516 10752 14522 10764
rect 5166 10684 5172 10736
rect 5224 10684 5230 10736
rect 10594 10684 10600 10736
rect 10652 10724 10658 10736
rect 13081 10727 13139 10733
rect 13081 10724 13093 10727
rect 10652 10696 13093 10724
rect 10652 10684 10658 10696
rect 13081 10693 13093 10696
rect 13127 10724 13139 10727
rect 13538 10724 13544 10736
rect 13127 10696 13544 10724
rect 13127 10693 13139 10696
rect 13081 10687 13139 10693
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 13814 10684 13820 10736
rect 13872 10684 13878 10736
rect 15120 10665 15148 10764
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 19426 10752 19432 10804
rect 19484 10792 19490 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19484 10764 19625 10792
rect 19484 10752 19490 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 20165 10795 20223 10801
rect 20165 10761 20177 10795
rect 20211 10761 20223 10795
rect 56870 10792 56876 10804
rect 56831 10764 56876 10792
rect 20165 10755 20223 10761
rect 20180 10724 20208 10755
rect 56870 10752 56876 10764
rect 56928 10752 56934 10804
rect 56962 10752 56968 10804
rect 57020 10792 57026 10804
rect 57517 10795 57575 10801
rect 57517 10792 57529 10795
rect 57020 10764 57529 10792
rect 57020 10752 57026 10764
rect 57517 10761 57529 10764
rect 57563 10792 57575 10795
rect 57698 10792 57704 10804
rect 57563 10764 57704 10792
rect 57563 10761 57575 10764
rect 57517 10755 57575 10761
rect 57698 10752 57704 10764
rect 57756 10752 57762 10804
rect 17052 10696 20208 10724
rect 3145 10659 3203 10665
rect 3145 10656 3157 10659
rect 2363 10628 2636 10656
rect 2700 10628 3157 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2130 10588 2136 10600
rect 2043 10560 2136 10588
rect 2130 10548 2136 10560
rect 2188 10548 2194 10600
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2498 10588 2504 10600
rect 2271 10560 2504 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 2608 10588 2636 10628
rect 3145 10625 3157 10628
rect 3191 10625 3203 10659
rect 3145 10619 3203 10625
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 3050 10588 3056 10600
rect 2608 10560 3056 10588
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5721 10591 5779 10597
rect 5721 10588 5733 10591
rect 5316 10560 5733 10588
rect 5316 10548 5322 10560
rect 5721 10557 5733 10560
rect 5767 10557 5779 10591
rect 5994 10588 6000 10600
rect 5955 10560 6000 10588
rect 5721 10551 5779 10557
rect 5994 10548 6000 10560
rect 6052 10548 6058 10600
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 17052 10588 17080 10696
rect 18506 10616 18512 10668
rect 18564 10656 18570 10668
rect 19153 10659 19211 10665
rect 19153 10656 19165 10659
rect 18564 10628 19165 10656
rect 18564 10616 18570 10628
rect 19153 10625 19165 10628
rect 19199 10625 19211 10659
rect 19153 10619 19211 10625
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10625 19303 10659
rect 19245 10619 19303 10625
rect 20349 10659 20407 10665
rect 20349 10625 20361 10659
rect 20395 10656 20407 10659
rect 20898 10656 20904 10668
rect 20395 10628 20904 10656
rect 20395 10625 20407 10628
rect 20349 10619 20407 10625
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 14875 10560 17080 10588
rect 17972 10560 18981 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 2148 10520 2176 10548
rect 2682 10520 2688 10532
rect 2148 10492 2688 10520
rect 2682 10480 2688 10492
rect 2740 10480 2746 10532
rect 3329 10523 3387 10529
rect 3329 10489 3341 10523
rect 3375 10520 3387 10523
rect 3375 10492 4752 10520
rect 3375 10489 3387 10492
rect 3329 10483 3387 10489
rect 2314 10412 2320 10464
rect 2372 10452 2378 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 2372 10424 4261 10452
rect 2372 10412 2378 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4724 10452 4752 10492
rect 9674 10452 9680 10464
rect 4724 10424 9680 10452
rect 4249 10415 4307 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 12526 10452 12532 10464
rect 12487 10424 12532 10452
rect 12526 10412 12532 10424
rect 12584 10452 12590 10464
rect 17972 10452 18000 10560
rect 18969 10557 18981 10560
rect 19015 10588 19027 10591
rect 19058 10588 19064 10600
rect 19015 10560 19064 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 18414 10520 18420 10532
rect 18327 10492 18420 10520
rect 12584 10424 18000 10452
rect 12584 10412 12590 10424
rect 18230 10412 18236 10464
rect 18288 10452 18294 10464
rect 18340 10461 18368 10492
rect 18414 10480 18420 10492
rect 18472 10520 18478 10532
rect 19260 10520 19288 10619
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 58345 10659 58403 10665
rect 58345 10625 58357 10659
rect 58391 10656 58403 10659
rect 58434 10656 58440 10668
rect 58391 10628 58440 10656
rect 58391 10625 58403 10628
rect 58345 10619 58403 10625
rect 58434 10616 58440 10628
rect 58492 10616 58498 10668
rect 18472 10492 19288 10520
rect 18472 10480 18478 10492
rect 18325 10455 18383 10461
rect 18325 10452 18337 10455
rect 18288 10424 18337 10452
rect 18288 10412 18294 10424
rect 18325 10421 18337 10424
rect 18371 10421 18383 10455
rect 18325 10415 18383 10421
rect 57606 10412 57612 10464
rect 57664 10452 57670 10464
rect 58161 10455 58219 10461
rect 58161 10452 58173 10455
rect 57664 10424 58173 10452
rect 57664 10412 57670 10424
rect 58161 10421 58173 10424
rect 58207 10421 58219 10455
rect 58161 10415 58219 10421
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 3050 10248 3056 10260
rect 2963 10220 3056 10248
rect 3050 10208 3056 10220
rect 3108 10248 3114 10260
rect 3326 10248 3332 10260
rect 3108 10220 3332 10248
rect 3108 10208 3114 10220
rect 3326 10208 3332 10220
rect 3384 10248 3390 10260
rect 3970 10248 3976 10260
rect 3384 10220 3976 10248
rect 3384 10208 3390 10220
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15102 10248 15108 10260
rect 15059 10220 15108 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15102 10208 15108 10220
rect 15160 10248 15166 10260
rect 18506 10248 18512 10260
rect 15160 10220 18276 10248
rect 18467 10220 18512 10248
rect 15160 10208 15166 10220
rect 2038 10140 2044 10192
rect 2096 10180 2102 10192
rect 5813 10183 5871 10189
rect 5813 10180 5825 10183
rect 2096 10152 5825 10180
rect 2096 10140 2102 10152
rect 5813 10149 5825 10152
rect 5859 10149 5871 10183
rect 18248 10180 18276 10220
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19116 10220 19717 10248
rect 19116 10208 19122 10220
rect 19705 10217 19717 10220
rect 19751 10248 19763 10251
rect 20622 10248 20628 10260
rect 19751 10220 20628 10248
rect 19751 10217 19763 10220
rect 19705 10211 19763 10217
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 58250 10208 58256 10260
rect 58308 10248 58314 10260
rect 58345 10251 58403 10257
rect 58345 10248 58357 10251
rect 58308 10220 58357 10248
rect 58308 10208 58314 10220
rect 58345 10217 58357 10220
rect 58391 10217 58403 10251
rect 58345 10211 58403 10217
rect 20162 10180 20168 10192
rect 18248 10152 20168 10180
rect 5813 10143 5871 10149
rect 20162 10140 20168 10152
rect 20220 10140 20226 10192
rect 57701 10183 57759 10189
rect 57701 10149 57713 10183
rect 57747 10180 57759 10183
rect 58434 10180 58440 10192
rect 57747 10152 58440 10180
rect 57747 10149 57759 10152
rect 57701 10143 57759 10149
rect 58434 10140 58440 10152
rect 58492 10140 58498 10192
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6914 10112 6920 10124
rect 6052 10084 6920 10112
rect 6052 10072 6058 10084
rect 6914 10072 6920 10084
rect 6972 10112 6978 10124
rect 6972 10084 7604 10112
rect 6972 10072 6978 10084
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 2406 10044 2412 10056
rect 1903 10016 2412 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 7576 10053 7604 10084
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 9088 10084 12265 10112
rect 9088 10072 9094 10084
rect 12253 10081 12265 10084
rect 12299 10112 12311 10115
rect 12526 10112 12532 10124
rect 12299 10084 12532 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 16758 10112 16764 10124
rect 16719 10084 16764 10112
rect 16758 10072 16764 10084
rect 16816 10072 16822 10124
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 9306 10044 9312 10056
rect 7607 10016 9312 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10044 12127 10047
rect 12158 10044 12164 10056
rect 12115 10016 12164 10044
rect 12115 10013 12127 10016
rect 12069 10007 12127 10013
rect 12158 10004 12164 10016
rect 12216 10044 12222 10056
rect 57149 10047 57207 10053
rect 12216 10016 12434 10044
rect 12216 10004 12222 10016
rect 5166 9936 5172 9988
rect 5224 9976 5230 9988
rect 5994 9976 6000 9988
rect 5224 9948 6000 9976
rect 5224 9936 5230 9948
rect 5994 9936 6000 9948
rect 6052 9976 6058 9988
rect 7282 9976 7288 9988
rect 6052 9948 6118 9976
rect 7243 9948 7288 9976
rect 6052 9936 6058 9948
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 2501 9911 2559 9917
rect 2501 9877 2513 9911
rect 2547 9908 2559 9911
rect 2682 9908 2688 9920
rect 2547 9880 2688 9908
rect 2547 9877 2559 9880
rect 2501 9871 2559 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11701 9911 11759 9917
rect 11701 9908 11713 9911
rect 11112 9880 11713 9908
rect 11112 9868 11118 9880
rect 11701 9877 11713 9880
rect 11747 9877 11759 9911
rect 11701 9871 11759 9877
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12406 9908 12434 10016
rect 57149 10013 57161 10047
rect 57195 10044 57207 10047
rect 58158 10044 58164 10056
rect 57195 10016 58164 10044
rect 57195 10013 57207 10016
rect 57149 10007 57207 10013
rect 58158 10004 58164 10016
rect 58216 10004 58222 10056
rect 16022 9936 16028 9988
rect 16080 9936 16086 9988
rect 16485 9979 16543 9985
rect 16485 9945 16497 9979
rect 16531 9976 16543 9979
rect 17862 9976 17868 9988
rect 16531 9948 17868 9976
rect 16531 9945 16543 9948
rect 16485 9939 16543 9945
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12216 9880 12261 9908
rect 12406 9880 13001 9908
rect 12216 9868 12222 9880
rect 12989 9877 13001 9880
rect 13035 9908 13047 9911
rect 14642 9908 14648 9920
rect 13035 9880 14648 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 9030 9704 9036 9716
rect 2740 9676 9036 9704
rect 2740 9664 2746 9676
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 9306 9664 9312 9716
rect 9364 9664 9370 9716
rect 56962 9704 56968 9716
rect 56923 9676 56968 9704
rect 56962 9664 56968 9676
rect 57020 9704 57026 9716
rect 57698 9704 57704 9716
rect 57020 9676 57704 9704
rect 57020 9664 57026 9676
rect 57698 9664 57704 9676
rect 57756 9664 57762 9716
rect 5166 9596 5172 9648
rect 5224 9596 5230 9648
rect 5721 9639 5779 9645
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 5810 9636 5816 9648
rect 5767 9608 5816 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 5994 9596 6000 9648
rect 6052 9636 6058 9648
rect 9324 9636 9352 9664
rect 13814 9636 13820 9648
rect 6052 9608 8510 9636
rect 9324 9608 9996 9636
rect 13662 9608 13820 9636
rect 6052 9596 6058 9608
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 4062 9568 4068 9580
rect 1903 9540 4068 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 9968 9577 9996 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14093 9639 14151 9645
rect 14093 9605 14105 9639
rect 14139 9636 14151 9639
rect 17770 9636 17776 9648
rect 14139 9608 17776 9636
rect 14139 9605 14151 9608
rect 14093 9599 14151 9605
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 20162 9596 20168 9648
rect 20220 9636 20226 9648
rect 20806 9636 20812 9648
rect 20220 9608 20576 9636
rect 20767 9608 20812 9636
rect 20220 9596 20226 9608
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20548 9568 20576 9608
rect 20806 9596 20812 9608
rect 20864 9596 20870 9648
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 19935 9540 20484 9568
rect 20548 9540 20913 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 2406 9500 2412 9512
rect 2319 9472 2412 9500
rect 2406 9460 2412 9472
rect 2464 9500 2470 9512
rect 5997 9503 6055 9509
rect 2464 9472 5948 9500
rect 2464 9460 2470 9472
rect 1670 9432 1676 9444
rect 1631 9404 1676 9432
rect 1670 9392 1676 9404
rect 1728 9392 1734 9444
rect 2222 9392 2228 9444
rect 2280 9432 2286 9444
rect 4249 9435 4307 9441
rect 4249 9432 4261 9435
rect 2280 9404 4261 9432
rect 2280 9392 2286 9404
rect 4249 9401 4261 9404
rect 4295 9401 4307 9435
rect 5920 9432 5948 9472
rect 5997 9469 6009 9503
rect 6043 9500 6055 9503
rect 6914 9500 6920 9512
rect 6043 9472 6920 9500
rect 6043 9469 6055 9472
rect 5997 9463 6055 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 9674 9500 9680 9512
rect 9635 9472 9680 9500
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 14458 9500 14464 9512
rect 14415 9472 14464 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 5920 9404 8708 9432
rect 4249 9395 4307 9401
rect 8202 9364 8208 9376
rect 8163 9336 8208 9364
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8680 9364 8708 9404
rect 17862 9392 17868 9444
rect 17920 9432 17926 9444
rect 20456 9441 20484 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 57517 9571 57575 9577
rect 57517 9537 57529 9571
rect 57563 9568 57575 9571
rect 58158 9568 58164 9580
rect 57563 9540 58164 9568
rect 57563 9537 57575 9540
rect 57517 9531 57575 9537
rect 58158 9528 58164 9540
rect 58216 9528 58222 9580
rect 21082 9500 21088 9512
rect 21043 9472 21088 9500
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 19705 9435 19763 9441
rect 19705 9432 19717 9435
rect 17920 9404 19717 9432
rect 17920 9392 17926 9404
rect 19705 9401 19717 9404
rect 19751 9401 19763 9435
rect 19705 9395 19763 9401
rect 20441 9435 20499 9441
rect 20441 9401 20453 9435
rect 20487 9401 20499 9435
rect 58342 9432 58348 9444
rect 58303 9404 58348 9432
rect 20441 9395 20499 9401
rect 58342 9392 58348 9404
rect 58400 9392 58406 9444
rect 12621 9367 12679 9373
rect 12621 9364 12633 9367
rect 8680 9336 12633 9364
rect 12621 9333 12633 9336
rect 12667 9364 12679 9367
rect 13538 9364 13544 9376
rect 12667 9336 13544 9364
rect 12667 9333 12679 9336
rect 12621 9327 12679 9333
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2740 9132 2789 9160
rect 2740 9120 2746 9132
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 2777 9123 2835 9129
rect 5166 9120 5172 9172
rect 5224 9160 5230 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 5224 9132 5641 9160
rect 5224 9120 5230 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 6362 9160 6368 9172
rect 6323 9132 6368 9160
rect 5629 9123 5687 9129
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 12158 9160 12164 9172
rect 9232 9132 12164 9160
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 8202 9092 8208 9104
rect 2556 9064 8208 9092
rect 2556 9052 2562 9064
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 4062 8984 4068 9036
rect 4120 9024 4126 9036
rect 9232 9024 9260 9132
rect 12158 9120 12164 9132
rect 12216 9160 12222 9172
rect 12529 9163 12587 9169
rect 12529 9160 12541 9163
rect 12216 9132 12541 9160
rect 12216 9120 12222 9132
rect 12529 9129 12541 9132
rect 12575 9129 12587 9163
rect 13170 9160 13176 9172
rect 13131 9132 13176 9160
rect 12529 9123 12587 9129
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 14366 9160 14372 9172
rect 14327 9132 14372 9160
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 20162 9120 20168 9172
rect 20220 9160 20226 9172
rect 20257 9163 20315 9169
rect 20257 9160 20269 9163
rect 20220 9132 20269 9160
rect 20220 9120 20226 9132
rect 20257 9129 20269 9132
rect 20303 9129 20315 9163
rect 20257 9123 20315 9129
rect 57790 9120 57796 9172
rect 57848 9160 57854 9172
rect 57848 9132 58204 9160
rect 57848 9120 57854 9132
rect 57624 9064 58112 9092
rect 4120 8996 9260 9024
rect 4120 8984 4126 8996
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 10781 9027 10839 9033
rect 10781 9024 10793 9027
rect 9364 8996 10793 9024
rect 9364 8984 9370 8996
rect 10781 8993 10793 8996
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 20346 8984 20352 9036
rect 20404 9024 20410 9036
rect 21637 9027 21695 9033
rect 21637 9024 21649 9027
rect 20404 8996 21649 9024
rect 20404 8984 20410 8996
rect 21637 8993 21649 8996
rect 21683 9024 21695 9027
rect 22738 9024 22744 9036
rect 21683 8996 22744 9024
rect 21683 8993 21695 8996
rect 21637 8987 21695 8993
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 56045 9027 56103 9033
rect 56045 8993 56057 9027
rect 56091 9024 56103 9027
rect 56962 9024 56968 9036
rect 56091 8996 56968 9024
rect 56091 8993 56103 8996
rect 56045 8987 56103 8993
rect 56962 8984 56968 8996
rect 57020 9024 57026 9036
rect 57330 9033 57336 9036
rect 57149 9027 57207 9033
rect 57149 9024 57161 9027
rect 57020 8996 57161 9024
rect 57020 8984 57026 8996
rect 57149 8993 57161 8996
rect 57195 8993 57207 9027
rect 57149 8987 57207 8993
rect 57308 9027 57336 9033
rect 57308 8993 57320 9027
rect 57308 8987 57336 8993
rect 57330 8984 57336 8987
rect 57388 8984 57394 9036
rect 57425 9027 57483 9033
rect 57425 8993 57437 9027
rect 57471 9024 57483 9027
rect 57624 9024 57652 9064
rect 57471 8996 57652 9024
rect 57471 8993 57483 8996
rect 57425 8987 57483 8993
rect 57698 8984 57704 9036
rect 57756 9024 57762 9036
rect 57756 8996 57801 9024
rect 57756 8984 57762 8996
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8956 1915 8959
rect 2222 8956 2228 8968
rect 1903 8928 2228 8956
rect 1903 8925 1915 8928
rect 1857 8919 1915 8925
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8956 5871 8959
rect 6362 8956 6368 8968
rect 5859 8928 6368 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 6362 8916 6368 8928
rect 6420 8916 6426 8968
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10152 8888 10180 8919
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12952 8928 13001 8956
rect 12952 8916 12958 8928
rect 12989 8925 13001 8928
rect 13035 8956 13047 8959
rect 14366 8956 14372 8968
rect 13035 8928 14372 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 20806 8916 20812 8968
rect 20864 8956 20870 8968
rect 21913 8959 21971 8965
rect 21913 8956 21925 8959
rect 20864 8928 21925 8956
rect 20864 8916 20870 8928
rect 21913 8925 21925 8928
rect 21959 8956 21971 8959
rect 58084 8956 58112 9064
rect 58176 9033 58204 9132
rect 58161 9027 58219 9033
rect 58161 8993 58173 9027
rect 58207 8993 58219 9027
rect 58161 8987 58219 8993
rect 58342 8956 58348 8968
rect 21959 8928 22094 8956
rect 58084 8928 58204 8956
rect 58303 8928 58348 8956
rect 21959 8925 21971 8928
rect 21913 8919 21971 8925
rect 10962 8888 10968 8900
rect 10152 8860 10968 8888
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 11057 8891 11115 8897
rect 11057 8857 11069 8891
rect 11103 8857 11115 8891
rect 13170 8888 13176 8900
rect 12282 8860 13176 8888
rect 11057 8851 11115 8857
rect 10321 8823 10379 8829
rect 10321 8789 10333 8823
rect 10367 8820 10379 8823
rect 11072 8820 11100 8851
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 22066 8888 22094 8928
rect 22462 8888 22468 8900
rect 22066 8860 22468 8888
rect 22462 8848 22468 8860
rect 22520 8848 22526 8900
rect 58176 8888 58204 8928
rect 58342 8916 58348 8928
rect 58400 8916 58406 8968
rect 58894 8888 58900 8900
rect 58176 8860 58900 8888
rect 58894 8848 58900 8860
rect 58952 8848 58958 8900
rect 20990 8820 20996 8832
rect 10367 8792 11100 8820
rect 20951 8792 20996 8820
rect 10367 8789 10379 8792
rect 10321 8783 10379 8789
rect 20990 8780 20996 8792
rect 21048 8820 21054 8832
rect 21821 8823 21879 8829
rect 21821 8820 21833 8823
rect 21048 8792 21833 8820
rect 21048 8780 21054 8792
rect 21821 8789 21833 8792
rect 21867 8789 21879 8823
rect 21821 8783 21879 8789
rect 22186 8780 22192 8832
rect 22244 8820 22250 8832
rect 22281 8823 22339 8829
rect 22281 8820 22293 8823
rect 22244 8792 22293 8820
rect 22244 8780 22250 8792
rect 22281 8789 22293 8792
rect 22327 8789 22339 8823
rect 22738 8820 22744 8832
rect 22699 8792 22744 8820
rect 22281 8783 22339 8789
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 56502 8820 56508 8832
rect 56463 8792 56508 8820
rect 56502 8780 56508 8792
rect 56560 8780 56566 8832
rect 56870 8780 56876 8832
rect 56928 8820 56934 8832
rect 58250 8820 58256 8832
rect 56928 8792 58256 8820
rect 56928 8780 56934 8792
rect 58250 8780 58256 8792
rect 58308 8780 58314 8832
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 2685 8619 2743 8625
rect 2685 8585 2697 8619
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2700 8480 2728 8579
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3789 8619 3847 8625
rect 3789 8616 3801 8619
rect 3476 8588 3801 8616
rect 3476 8576 3482 8588
rect 3789 8585 3801 8588
rect 3835 8616 3847 8619
rect 4062 8616 4068 8628
rect 3835 8588 4068 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 6362 8576 6368 8628
rect 6420 8616 6426 8628
rect 12894 8616 12900 8628
rect 6420 8588 12900 8616
rect 6420 8576 6426 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 14458 8616 14464 8628
rect 14419 8588 14464 8616
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 57333 8619 57391 8625
rect 57333 8585 57345 8619
rect 57379 8616 57391 8619
rect 58066 8616 58072 8628
rect 57379 8588 58072 8616
rect 57379 8585 57391 8588
rect 57333 8579 57391 8585
rect 58066 8576 58072 8588
rect 58124 8576 58130 8628
rect 58342 8616 58348 8628
rect 58303 8588 58348 8616
rect 58342 8576 58348 8588
rect 58400 8576 58406 8628
rect 12529 8551 12587 8557
rect 12529 8517 12541 8551
rect 12575 8548 12587 8551
rect 12802 8548 12808 8560
rect 12575 8520 12808 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 12802 8508 12808 8520
rect 12860 8548 12866 8560
rect 12989 8551 13047 8557
rect 12989 8548 13001 8551
rect 12860 8520 13001 8548
rect 12860 8508 12866 8520
rect 12989 8517 13001 8520
rect 13035 8517 13047 8551
rect 12989 8511 13047 8517
rect 56134 8508 56140 8560
rect 56192 8548 56198 8560
rect 56229 8551 56287 8557
rect 56229 8548 56241 8551
rect 56192 8520 56241 8548
rect 56192 8508 56198 8520
rect 56229 8517 56241 8520
rect 56275 8517 56287 8551
rect 56229 8511 56287 8517
rect 56597 8551 56655 8557
rect 56597 8517 56609 8551
rect 56643 8548 56655 8551
rect 56870 8548 56876 8560
rect 56643 8520 56876 8548
rect 56643 8517 56655 8520
rect 56597 8511 56655 8517
rect 56870 8508 56876 8520
rect 56928 8508 56934 8560
rect 58526 8548 58532 8560
rect 57256 8520 58532 8548
rect 3145 8483 3203 8489
rect 3145 8480 3157 8483
rect 2700 8452 3157 8480
rect 2317 8443 2375 8449
rect 3145 8449 3157 8452
rect 3191 8449 3203 8483
rect 22186 8480 22192 8492
rect 22147 8452 22192 8480
rect 3145 8443 3203 8449
rect 2041 8415 2099 8421
rect 2041 8381 2053 8415
rect 2087 8381 2099 8415
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 2041 8375 2099 8381
rect 2056 8344 2084 8375
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2332 8412 2360 8443
rect 22186 8440 22192 8452
rect 22244 8440 22250 8492
rect 56962 8480 56968 8492
rect 56923 8452 56968 8480
rect 56962 8440 56968 8452
rect 57020 8440 57026 8492
rect 57057 8483 57115 8489
rect 57057 8449 57069 8483
rect 57103 8480 57115 8483
rect 57256 8480 57284 8520
rect 58526 8508 58532 8520
rect 58584 8508 58590 8560
rect 57103 8452 57284 8480
rect 57103 8449 57115 8452
rect 57057 8443 57115 8449
rect 58158 8440 58164 8492
rect 58216 8480 58222 8492
rect 58216 8452 58261 8480
rect 58216 8440 58222 8452
rect 3418 8412 3424 8424
rect 2332 8384 3424 8412
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 57698 8412 57704 8424
rect 57546 8384 57704 8412
rect 57698 8372 57704 8384
rect 57756 8372 57762 8424
rect 2130 8344 2136 8356
rect 2043 8316 2136 8344
rect 2130 8304 2136 8316
rect 2188 8344 2194 8356
rect 2682 8344 2688 8356
rect 2188 8316 2688 8344
rect 2188 8304 2194 8316
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 5902 8344 5908 8356
rect 3375 8316 5908 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 53834 8304 53840 8356
rect 53892 8344 53898 8356
rect 56045 8347 56103 8353
rect 56045 8344 56057 8347
rect 53892 8316 56057 8344
rect 53892 8304 53898 8316
rect 56045 8313 56057 8316
rect 56091 8313 56103 8347
rect 56045 8307 56103 8313
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 20990 8276 20996 8288
rect 15712 8248 20996 8276
rect 15712 8236 15718 8248
rect 20990 8236 20996 8248
rect 21048 8236 21054 8288
rect 22002 8276 22008 8288
rect 21963 8248 22008 8276
rect 22002 8236 22008 8248
rect 22060 8236 22066 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1670 8072 1676 8084
rect 1631 8044 1676 8072
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 2222 8032 2228 8084
rect 2280 8072 2286 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 2280 8044 4445 8072
rect 2280 8032 2286 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 4433 8035 4491 8041
rect 56962 8032 56968 8084
rect 57020 8072 57026 8084
rect 57057 8075 57115 8081
rect 57057 8072 57069 8075
rect 57020 8044 57069 8072
rect 57020 8032 57026 8044
rect 57057 8041 57069 8044
rect 57103 8041 57115 8075
rect 57698 8072 57704 8084
rect 57659 8044 57704 8072
rect 57057 8035 57115 8041
rect 57698 8032 57704 8044
rect 57756 8032 57762 8084
rect 58161 8075 58219 8081
rect 58161 8041 58173 8075
rect 58207 8072 58219 8075
rect 58250 8072 58256 8084
rect 58207 8044 58256 8072
rect 58207 8041 58219 8044
rect 58161 8035 58219 8041
rect 58250 8032 58256 8044
rect 58308 8032 58314 8084
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 3053 8007 3111 8013
rect 3053 8004 3065 8007
rect 2740 7976 3065 8004
rect 2740 7964 2746 7976
rect 3053 7973 3065 7976
rect 3099 7973 3111 8007
rect 3053 7967 3111 7973
rect 2498 7936 2504 7948
rect 1872 7908 2504 7936
rect 1872 7877 1900 7908
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 5902 7936 5908 7948
rect 5863 7908 5908 7936
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15712 7908 15853 7936
rect 15712 7896 15718 7908
rect 15841 7905 15853 7908
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 17589 7939 17647 7945
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 22002 7936 22008 7948
rect 17635 7908 22008 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 22002 7896 22008 7908
rect 22060 7896 22066 7948
rect 22554 7936 22560 7948
rect 22515 7908 22560 7936
rect 22554 7896 22560 7908
rect 22612 7896 22618 7948
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 2314 7828 2320 7880
rect 2372 7868 2378 7880
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2372 7840 2605 7868
rect 2372 7828 2378 7840
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 5350 7760 5356 7812
rect 5408 7760 5414 7812
rect 5994 7760 6000 7812
rect 6052 7800 6058 7812
rect 6196 7800 6224 7831
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 21729 7871 21787 7877
rect 17920 7840 17965 7868
rect 17920 7828 17926 7840
rect 21729 7837 21741 7871
rect 21775 7868 21787 7871
rect 22278 7868 22284 7880
rect 21775 7840 22284 7868
rect 21775 7837 21787 7840
rect 21729 7831 21787 7837
rect 22278 7828 22284 7840
rect 22336 7828 22342 7880
rect 22649 7871 22707 7877
rect 22649 7837 22661 7871
rect 22695 7837 22707 7871
rect 58342 7868 58348 7880
rect 58303 7840 58348 7868
rect 22649 7831 22707 7837
rect 6052 7772 6224 7800
rect 6052 7760 6058 7772
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 21177 7803 21235 7809
rect 13872 7772 16422 7800
rect 13872 7760 13878 7772
rect 21177 7769 21189 7803
rect 21223 7800 21235 7803
rect 22664 7800 22692 7831
rect 58342 7828 58348 7840
rect 58400 7828 58406 7880
rect 22830 7800 22836 7812
rect 21223 7772 22836 7800
rect 21223 7769 21235 7772
rect 21177 7763 21235 7769
rect 22830 7760 22836 7772
rect 22888 7760 22894 7812
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2682 7528 2688 7540
rect 2455 7500 2688 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 2777 7531 2835 7537
rect 2777 7497 2789 7531
rect 2823 7497 2835 7531
rect 2777 7491 2835 7497
rect 2792 7392 2820 7491
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 3881 7531 3939 7537
rect 3881 7528 3893 7531
rect 2924 7500 3893 7528
rect 2924 7488 2930 7500
rect 3881 7497 3893 7500
rect 3927 7528 3939 7531
rect 3970 7528 3976 7540
rect 3927 7500 3976 7528
rect 3927 7497 3939 7500
rect 3881 7491 3939 7497
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 9306 7528 9312 7540
rect 8343 7500 9312 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 10928 7500 13829 7528
rect 10928 7488 10934 7500
rect 13817 7497 13829 7500
rect 13863 7497 13875 7531
rect 19429 7531 19487 7537
rect 19429 7528 19441 7531
rect 13817 7491 13875 7497
rect 15304 7500 19441 7528
rect 3237 7395 3295 7401
rect 3237 7392 3249 7395
rect 2792 7364 3249 7392
rect 3237 7361 3249 7364
rect 3283 7361 3295 7395
rect 9582 7392 9588 7404
rect 9543 7364 9588 7392
rect 3237 7355 3295 7361
rect 9582 7352 9588 7364
rect 9640 7392 9646 7404
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9640 7364 10057 7392
rect 9640 7352 9646 7364
rect 10045 7361 10057 7364
rect 10091 7392 10103 7395
rect 12802 7392 12808 7404
rect 10091 7364 12808 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 2130 7324 2136 7336
rect 2091 7296 2136 7324
rect 2130 7284 2136 7296
rect 2188 7284 2194 7336
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 2498 7324 2504 7336
rect 2363 7296 2504 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 13832 7324 13860 7491
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 15304 7469 15332 7500
rect 19429 7497 19441 7500
rect 19475 7497 19487 7531
rect 19429 7491 19487 7497
rect 57517 7531 57575 7537
rect 57517 7497 57529 7531
rect 57563 7528 57575 7531
rect 58342 7528 58348 7540
rect 57563 7500 58348 7528
rect 57563 7497 57575 7500
rect 57517 7491 57575 7497
rect 58342 7488 58348 7500
rect 58400 7488 58406 7540
rect 15289 7463 15347 7469
rect 13964 7432 14122 7460
rect 13964 7420 13970 7432
rect 15289 7429 15301 7463
rect 15335 7429 15347 7463
rect 15289 7423 15347 7429
rect 22649 7463 22707 7469
rect 22649 7429 22661 7463
rect 22695 7460 22707 7463
rect 22738 7460 22744 7472
rect 22695 7432 22744 7460
rect 22695 7429 22707 7432
rect 22649 7423 22707 7429
rect 22738 7420 22744 7432
rect 22796 7420 22802 7472
rect 58158 7420 58164 7472
rect 58216 7460 58222 7472
rect 58253 7463 58311 7469
rect 58253 7460 58265 7463
rect 58216 7432 58265 7460
rect 58216 7420 58222 7432
rect 58253 7429 58265 7432
rect 58299 7429 58311 7463
rect 58253 7423 58311 7429
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 16850 7392 16856 7404
rect 15611 7364 16856 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 16850 7352 16856 7364
rect 16908 7392 16914 7404
rect 17862 7392 17868 7404
rect 16908 7364 17868 7392
rect 16908 7352 16914 7364
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 19978 7392 19984 7404
rect 19659 7364 19984 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 22189 7395 22247 7401
rect 22189 7392 22201 7395
rect 21499 7364 22201 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 22189 7361 22201 7364
rect 22235 7392 22247 7395
rect 22278 7392 22284 7404
rect 22235 7364 22284 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 22278 7352 22284 7364
rect 22336 7352 22342 7404
rect 22830 7392 22836 7404
rect 22791 7364 22836 7392
rect 22830 7352 22836 7364
rect 22888 7392 22894 7404
rect 23569 7395 23627 7401
rect 23569 7392 23581 7395
rect 22888 7364 23581 7392
rect 22888 7352 22894 7364
rect 23569 7361 23581 7364
rect 23615 7361 23627 7395
rect 23569 7355 23627 7361
rect 18782 7324 18788 7336
rect 13832 7296 18788 7324
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 3418 7188 3424 7200
rect 3379 7160 3424 7188
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 56962 7188 56968 7200
rect 56923 7160 56968 7188
rect 56962 7148 56968 7160
rect 57020 7148 57026 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 8309 6987 8367 6993
rect 8309 6984 8321 6987
rect 3476 6956 8321 6984
rect 3476 6944 3482 6956
rect 8309 6953 8321 6956
rect 8355 6953 8367 6987
rect 8309 6947 8367 6953
rect 21082 6944 21088 6996
rect 21140 6984 21146 6996
rect 22465 6987 22523 6993
rect 22465 6984 22477 6987
rect 21140 6956 22477 6984
rect 21140 6944 21146 6956
rect 22465 6953 22477 6956
rect 22511 6953 22523 6987
rect 22465 6947 22523 6953
rect 57054 6944 57060 6996
rect 57112 6984 57118 6996
rect 57698 6984 57704 6996
rect 57112 6956 57704 6984
rect 57112 6944 57118 6956
rect 57698 6944 57704 6956
rect 57756 6944 57762 6996
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 2225 6851 2283 6857
rect 2225 6848 2237 6851
rect 2188 6820 2237 6848
rect 2188 6808 2194 6820
rect 2225 6817 2237 6820
rect 2271 6848 2283 6851
rect 2866 6848 2872 6860
rect 2271 6820 2872 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6817 6883 6851
rect 20622 6848 20628 6860
rect 20583 6820 20628 6848
rect 6825 6811 6883 6817
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 6840 6780 6868 6811
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 22278 6848 22284 6860
rect 22020 6820 22284 6848
rect 2556 6752 6868 6780
rect 2556 6740 2562 6752
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 8628 6752 8673 6780
rect 8628 6740 8634 6752
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 22020 6789 22048 6820
rect 22278 6808 22284 6820
rect 22336 6808 22342 6860
rect 57057 6851 57115 6857
rect 57057 6848 57069 6851
rect 56888 6820 57069 6848
rect 56888 6792 56916 6820
rect 57057 6817 57069 6820
rect 57103 6848 57115 6851
rect 57698 6848 57704 6860
rect 57103 6820 57704 6848
rect 57103 6817 57115 6820
rect 57057 6811 57115 6817
rect 57698 6808 57704 6820
rect 57756 6808 57762 6860
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19484 6752 19717 6780
rect 19484 6740 19490 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 20901 6783 20959 6789
rect 20901 6749 20913 6783
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 22005 6783 22063 6789
rect 22005 6749 22017 6783
rect 22051 6749 22063 6783
rect 22005 6743 22063 6749
rect 2409 6715 2467 6721
rect 2409 6681 2421 6715
rect 2455 6712 2467 6715
rect 2455 6684 3280 6712
rect 2455 6681 2467 6684
rect 2409 6675 2467 6681
rect 3252 6656 3280 6684
rect 5350 6672 5356 6724
rect 5408 6712 5414 6724
rect 9398 6712 9404 6724
rect 5408 6684 6914 6712
rect 7866 6684 9404 6712
rect 5408 6672 5414 6684
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2774 6644 2780 6656
rect 2735 6616 2780 6644
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 3234 6604 3240 6656
rect 3292 6644 3298 6656
rect 3329 6647 3387 6653
rect 3329 6644 3341 6647
rect 3292 6616 3341 6644
rect 3292 6604 3298 6616
rect 3329 6613 3341 6616
rect 3375 6644 3387 6647
rect 3510 6644 3516 6656
rect 3375 6616 3516 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 6886 6644 6914 6684
rect 7944 6644 7972 6684
rect 9398 6672 9404 6684
rect 9456 6672 9462 6724
rect 20916 6712 20944 6743
rect 22186 6740 22192 6792
rect 22244 6780 22250 6792
rect 22922 6780 22928 6792
rect 22244 6752 22928 6780
rect 22244 6740 22250 6752
rect 22922 6740 22928 6752
rect 22980 6740 22986 6792
rect 55398 6740 55404 6792
rect 55456 6780 55462 6792
rect 55677 6783 55735 6789
rect 55677 6780 55689 6783
rect 55456 6752 55689 6780
rect 55456 6740 55462 6752
rect 55677 6749 55689 6752
rect 55723 6780 55735 6783
rect 56042 6780 56048 6792
rect 55723 6752 56048 6780
rect 55723 6749 55735 6752
rect 55677 6743 55735 6749
rect 56042 6740 56048 6752
rect 56100 6780 56106 6792
rect 56229 6783 56287 6789
rect 56229 6780 56241 6783
rect 56100 6752 56241 6780
rect 56100 6740 56106 6752
rect 56229 6749 56241 6752
rect 56275 6749 56287 6783
rect 56229 6743 56287 6749
rect 56597 6783 56655 6789
rect 56597 6749 56609 6783
rect 56643 6780 56655 6783
rect 56870 6780 56876 6792
rect 56643 6752 56876 6780
rect 56643 6749 56655 6752
rect 56597 6743 56655 6749
rect 56870 6740 56876 6752
rect 56928 6740 56934 6792
rect 56962 6740 56968 6792
rect 57020 6780 57026 6792
rect 58342 6780 58348 6792
rect 57020 6752 58348 6780
rect 57020 6740 57026 6752
rect 58342 6740 58348 6752
rect 58400 6740 58406 6792
rect 22094 6712 22100 6724
rect 20916 6684 22100 6712
rect 22094 6672 22100 6684
rect 22152 6672 22158 6724
rect 6886 6616 7972 6644
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 19521 6647 19579 6653
rect 19521 6644 19533 6647
rect 17828 6616 19533 6644
rect 17828 6604 17834 6616
rect 19521 6613 19533 6616
rect 19567 6613 19579 6647
rect 19521 6607 19579 6613
rect 21545 6647 21603 6653
rect 21545 6613 21557 6647
rect 21591 6644 21603 6647
rect 22278 6644 22284 6656
rect 21591 6616 22284 6644
rect 21591 6613 21603 6616
rect 21545 6607 21603 6613
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 58158 6644 58164 6656
rect 58119 6616 58164 6644
rect 58158 6604 58164 6616
rect 58216 6604 58222 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 4249 6443 4307 6449
rect 4249 6440 4261 6443
rect 2372 6412 4261 6440
rect 2372 6400 2378 6412
rect 4249 6409 4261 6412
rect 4295 6409 4307 6443
rect 4249 6403 4307 6409
rect 5350 6400 5356 6452
rect 5408 6400 5414 6452
rect 14734 6440 14740 6452
rect 13188 6412 14740 6440
rect 5368 6372 5396 6400
rect 9582 6372 9588 6384
rect 5290 6344 5396 6372
rect 9543 6344 9588 6372
rect 9582 6332 9588 6344
rect 9640 6372 9646 6384
rect 10045 6375 10103 6381
rect 10045 6372 10057 6375
rect 9640 6344 10057 6372
rect 9640 6332 9646 6344
rect 10045 6341 10057 6344
rect 10091 6341 10103 6375
rect 10045 6335 10103 6341
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2222 6304 2228 6316
rect 1903 6276 2228 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 2774 6304 2780 6316
rect 2639 6276 2780 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 13188 6313 13216 6412
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 19242 6440 19248 6452
rect 19203 6412 19248 6440
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 19426 6400 19432 6452
rect 19484 6440 19490 6452
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 19484 6412 19717 6440
rect 19484 6400 19490 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 58158 6440 58164 6452
rect 19705 6403 19763 6409
rect 55692 6412 58164 6440
rect 13446 6372 13452 6384
rect 13407 6344 13452 6372
rect 13446 6332 13452 6344
rect 13504 6332 13510 6384
rect 13906 6332 13912 6384
rect 13964 6332 13970 6384
rect 18693 6375 18751 6381
rect 18693 6341 18705 6375
rect 18739 6372 18751 6375
rect 20165 6375 20223 6381
rect 20165 6372 20177 6375
rect 18739 6344 20177 6372
rect 18739 6341 18751 6344
rect 18693 6335 18751 6341
rect 20165 6341 20177 6344
rect 20211 6341 20223 6375
rect 20165 6335 20223 6341
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6273 13231 6307
rect 18708 6304 18736 6335
rect 13173 6267 13231 6273
rect 14660 6276 18736 6304
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 2792 6208 5733 6236
rect 2792 6177 2820 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5994 6236 6000 6248
rect 5955 6208 6000 6236
rect 5721 6199 5779 6205
rect 5994 6196 6000 6208
rect 6052 6236 6058 6248
rect 12713 6239 12771 6245
rect 6052 6208 8340 6236
rect 6052 6196 6058 6208
rect 2777 6171 2835 6177
rect 2777 6137 2789 6171
rect 2823 6137 2835 6171
rect 2777 6131 2835 6137
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 8312 6109 8340 6208
rect 12713 6205 12725 6239
rect 12759 6236 12771 6239
rect 13446 6236 13452 6248
rect 12759 6208 13452 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 14660 6236 14688 6276
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 55692 6313 55720 6412
rect 58158 6400 58164 6412
rect 58216 6400 58222 6452
rect 20073 6307 20131 6313
rect 20073 6304 20085 6307
rect 19300 6276 20085 6304
rect 19300 6264 19306 6276
rect 20073 6273 20085 6276
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 55677 6307 55735 6313
rect 55677 6273 55689 6307
rect 55723 6273 55735 6307
rect 55677 6267 55735 6273
rect 56686 6264 56692 6316
rect 56744 6313 56750 6316
rect 56744 6307 56772 6313
rect 56760 6273 56772 6307
rect 56870 6304 56876 6316
rect 56831 6276 56876 6304
rect 56744 6267 56772 6273
rect 56744 6264 56750 6267
rect 56870 6264 56876 6276
rect 56928 6264 56934 6316
rect 58342 6304 58348 6316
rect 58303 6276 58348 6304
rect 58342 6264 58348 6276
rect 58400 6264 58406 6316
rect 14918 6236 14924 6248
rect 13596 6208 14688 6236
rect 14879 6208 14924 6236
rect 13596 6196 13602 6208
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 18690 6196 18696 6248
rect 18748 6236 18754 6248
rect 19260 6236 19288 6264
rect 18748 6208 19288 6236
rect 20349 6239 20407 6245
rect 18748 6196 18754 6208
rect 20349 6205 20361 6239
rect 20395 6236 20407 6239
rect 20622 6236 20628 6248
rect 20395 6208 20628 6236
rect 20395 6205 20407 6208
rect 20349 6199 20407 6205
rect 20622 6196 20628 6208
rect 20680 6236 20686 6248
rect 20901 6239 20959 6245
rect 20901 6236 20913 6239
rect 20680 6208 20913 6236
rect 20680 6196 20686 6208
rect 20901 6205 20913 6208
rect 20947 6205 20959 6239
rect 55858 6236 55864 6248
rect 55819 6208 55864 6236
rect 20901 6199 20959 6205
rect 55858 6196 55864 6208
rect 55916 6196 55922 6248
rect 56597 6239 56655 6245
rect 56597 6205 56609 6239
rect 56643 6236 56655 6239
rect 58802 6236 58808 6248
rect 56643 6208 58808 6236
rect 56643 6205 56655 6208
rect 56597 6199 56655 6205
rect 58802 6196 58808 6208
rect 58860 6196 58866 6248
rect 56321 6171 56379 6177
rect 56321 6137 56333 6171
rect 56367 6137 56379 6171
rect 56321 6131 56379 6137
rect 3237 6103 3295 6109
rect 3237 6100 3249 6103
rect 2924 6072 3249 6100
rect 2924 6060 2930 6072
rect 3237 6069 3249 6072
rect 3283 6069 3295 6103
rect 3237 6063 3295 6069
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 8570 6100 8576 6112
rect 8343 6072 8576 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 8570 6060 8576 6072
rect 8628 6100 8634 6112
rect 9490 6100 9496 6112
rect 8628 6072 9496 6100
rect 8628 6060 8634 6072
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 22097 6103 22155 6109
rect 22097 6069 22109 6103
rect 22143 6100 22155 6103
rect 22186 6100 22192 6112
rect 22143 6072 22192 6100
rect 22143 6069 22155 6072
rect 22097 6063 22155 6069
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 56336 6100 56364 6131
rect 57054 6100 57060 6112
rect 56336 6072 57060 6100
rect 57054 6060 57060 6072
rect 57112 6060 57118 6112
rect 57238 6060 57244 6112
rect 57296 6100 57302 6112
rect 57517 6103 57575 6109
rect 57517 6100 57529 6103
rect 57296 6072 57529 6100
rect 57296 6060 57302 6072
rect 57517 6069 57529 6072
rect 57563 6069 57575 6103
rect 58158 6100 58164 6112
rect 58119 6072 58164 6100
rect 57517 6063 57575 6069
rect 58158 6060 58164 6072
rect 58216 6060 58222 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1670 5896 1676 5908
rect 1631 5868 1676 5896
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 10796 5868 12081 5896
rect 9769 5763 9827 5769
rect 9769 5729 9781 5763
rect 9815 5760 9827 5763
rect 10796 5760 10824 5868
rect 12069 5865 12081 5868
rect 12115 5896 12127 5899
rect 13078 5896 13084 5908
rect 12115 5868 13084 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 18782 5896 18788 5908
rect 18743 5868 18788 5896
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 19705 5899 19763 5905
rect 19705 5865 19717 5899
rect 19751 5896 19763 5899
rect 19978 5896 19984 5908
rect 19751 5868 19984 5896
rect 19751 5865 19763 5868
rect 19705 5859 19763 5865
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 58158 5896 58164 5908
rect 56520 5868 58164 5896
rect 11514 5760 11520 5772
rect 9815 5732 10824 5760
rect 11475 5732 11520 5760
rect 9815 5729 9827 5732
rect 9769 5723 9827 5729
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 18800 5760 18828 5856
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 18800 5732 20177 5760
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 20349 5763 20407 5769
rect 20349 5729 20361 5763
rect 20395 5760 20407 5763
rect 22094 5760 22100 5772
rect 20395 5732 22100 5760
rect 20395 5729 20407 5732
rect 20349 5723 20407 5729
rect 22094 5720 22100 5732
rect 22152 5720 22158 5772
rect 56520 5769 56548 5868
rect 58158 5856 58164 5868
rect 58216 5856 58222 5908
rect 57054 5788 57060 5840
rect 57112 5828 57118 5840
rect 57149 5831 57207 5837
rect 57149 5828 57161 5831
rect 57112 5800 57161 5828
rect 57112 5788 57118 5800
rect 57149 5797 57161 5800
rect 57195 5797 57207 5831
rect 57149 5791 57207 5797
rect 56505 5763 56563 5769
rect 56505 5729 56517 5763
rect 56551 5729 56563 5763
rect 57422 5760 57428 5772
rect 57383 5732 57428 5760
rect 56505 5723 56563 5729
rect 57422 5720 57428 5732
rect 57480 5720 57486 5772
rect 57606 5769 57612 5772
rect 57563 5763 57612 5769
rect 57563 5729 57575 5763
rect 57609 5729 57612 5763
rect 57563 5723 57612 5729
rect 57606 5720 57612 5723
rect 57664 5720 57670 5772
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2498 5692 2504 5704
rect 1903 5664 2504 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 9490 5692 9496 5704
rect 9451 5664 9496 5692
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 20073 5695 20131 5701
rect 20073 5661 20085 5695
rect 20119 5692 20131 5695
rect 20254 5692 20260 5704
rect 20119 5664 20260 5692
rect 20119 5661 20131 5664
rect 20073 5655 20131 5661
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 56686 5692 56692 5704
rect 56647 5664 56692 5692
rect 56686 5652 56692 5664
rect 56744 5652 56750 5704
rect 57698 5692 57704 5704
rect 57659 5664 57704 5692
rect 57698 5652 57704 5664
rect 57756 5652 57762 5704
rect 9398 5584 9404 5636
rect 9456 5624 9462 5636
rect 9456 5596 10258 5624
rect 9456 5584 9462 5596
rect 56045 5559 56103 5565
rect 56045 5525 56057 5559
rect 56091 5556 56103 5559
rect 57698 5556 57704 5568
rect 56091 5528 57704 5556
rect 56091 5525 56103 5528
rect 56045 5519 56103 5525
rect 57698 5516 57704 5528
rect 57756 5516 57762 5568
rect 58250 5516 58256 5568
rect 58308 5556 58314 5568
rect 58345 5559 58403 5565
rect 58345 5556 58357 5559
rect 58308 5528 58357 5556
rect 58308 5516 58314 5528
rect 58345 5525 58357 5528
rect 58391 5525 58403 5559
rect 58345 5519 58403 5525
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 12529 5355 12587 5361
rect 12529 5321 12541 5355
rect 12575 5352 12587 5355
rect 12802 5352 12808 5364
rect 12575 5324 12808 5352
rect 12575 5321 12587 5324
rect 12529 5315 12587 5321
rect 12802 5312 12808 5324
rect 12860 5312 12866 5364
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19613 5355 19671 5361
rect 19613 5352 19625 5355
rect 19484 5324 19625 5352
rect 19484 5312 19490 5324
rect 19613 5321 19625 5324
rect 19659 5352 19671 5355
rect 20254 5352 20260 5364
rect 19659 5324 20260 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 56965 5355 57023 5361
rect 56965 5321 56977 5355
rect 57011 5352 57023 5355
rect 57054 5352 57060 5364
rect 57011 5324 57060 5352
rect 57011 5321 57023 5324
rect 56965 5315 57023 5321
rect 57054 5312 57060 5324
rect 57112 5312 57118 5364
rect 57514 5352 57520 5364
rect 57475 5324 57520 5352
rect 57514 5312 57520 5324
rect 57572 5312 57578 5364
rect 58161 5355 58219 5361
rect 58161 5321 58173 5355
rect 58207 5352 58219 5355
rect 58710 5352 58716 5364
rect 58207 5324 58716 5352
rect 58207 5321 58219 5324
rect 58161 5315 58219 5321
rect 58710 5312 58716 5324
rect 58768 5312 58774 5364
rect 9398 5244 9404 5296
rect 9456 5244 9462 5296
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5284 10103 5287
rect 12820 5284 12848 5312
rect 12989 5287 13047 5293
rect 12989 5284 13001 5287
rect 10091 5256 12388 5284
rect 12820 5256 13001 5284
rect 10091 5253 10103 5256
rect 10045 5247 10103 5253
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 2406 5216 2412 5228
rect 1903 5188 2412 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 10318 5148 10324 5160
rect 10279 5120 10324 5148
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 1670 5080 1676 5092
rect 1631 5052 1676 5080
rect 1670 5040 1676 5052
rect 1728 5040 1734 5092
rect 12360 5080 12388 5256
rect 12989 5253 13001 5256
rect 13035 5253 13047 5287
rect 12989 5247 13047 5253
rect 56413 5219 56471 5225
rect 56413 5185 56425 5219
rect 56459 5216 56471 5219
rect 58342 5216 58348 5228
rect 56459 5188 58348 5216
rect 56459 5185 56471 5188
rect 56413 5179 56471 5185
rect 58342 5176 58348 5188
rect 58400 5176 58406 5228
rect 14734 5148 14740 5160
rect 14647 5120 14740 5148
rect 14734 5108 14740 5120
rect 14792 5148 14798 5160
rect 16850 5148 16856 5160
rect 14792 5120 16856 5148
rect 14792 5108 14798 5120
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 20714 5080 20720 5092
rect 12360 5052 20720 5080
rect 20714 5040 20720 5052
rect 20772 5040 20778 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 8570 5012 8576 5024
rect 7708 4984 8576 5012
rect 7708 4972 7714 4984
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 10318 5012 10324 5024
rect 9548 4984 10324 5012
rect 9548 4972 9554 4984
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5500 4780 5917 4808
rect 5500 4768 5506 4780
rect 5905 4777 5917 4780
rect 5951 4808 5963 4811
rect 5951 4780 6914 4808
rect 5951 4777 5963 4780
rect 5905 4771 5963 4777
rect 6454 4672 6460 4684
rect 6415 4644 6460 4672
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6886 4672 6914 4780
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 21637 4811 21695 4817
rect 21637 4808 21649 4811
rect 8628 4780 21649 4808
rect 8628 4768 8634 4780
rect 21637 4777 21649 4780
rect 21683 4808 21695 4811
rect 57701 4811 57759 4817
rect 21683 4780 22692 4808
rect 21683 4777 21695 4780
rect 21637 4771 21695 4777
rect 18966 4700 18972 4752
rect 19024 4740 19030 4752
rect 19429 4743 19487 4749
rect 19429 4740 19441 4743
rect 19024 4712 19441 4740
rect 19024 4700 19030 4712
rect 19429 4709 19441 4712
rect 19475 4709 19487 4743
rect 19429 4703 19487 4709
rect 8205 4675 8263 4681
rect 8205 4672 8217 4675
rect 6886 4644 8217 4672
rect 8205 4641 8217 4644
rect 8251 4641 8263 4675
rect 8205 4635 8263 4641
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 9490 4672 9496 4684
rect 8527 4644 9496 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 16850 4672 16856 4684
rect 16811 4644 16856 4672
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 17129 4675 17187 4681
rect 17129 4641 17141 4675
rect 17175 4672 17187 4675
rect 18138 4672 18144 4684
rect 17175 4644 18144 4672
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 18874 4672 18880 4684
rect 18835 4644 18880 4672
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 22664 4681 22692 4780
rect 57701 4777 57713 4811
rect 57747 4808 57759 4811
rect 57790 4808 57796 4820
rect 57747 4780 57796 4808
rect 57747 4777 57759 4780
rect 57701 4771 57759 4777
rect 57790 4768 57796 4780
rect 57848 4768 57854 4820
rect 57974 4768 57980 4820
rect 58032 4808 58038 4820
rect 58161 4811 58219 4817
rect 58161 4808 58173 4811
rect 58032 4780 58173 4808
rect 58032 4768 58038 4780
rect 58161 4777 58173 4780
rect 58207 4777 58219 4811
rect 58161 4771 58219 4777
rect 22649 4675 22707 4681
rect 22649 4641 22661 4675
rect 22695 4641 22707 4675
rect 22649 4635 22707 4641
rect 22741 4675 22799 4681
rect 22741 4641 22753 4675
rect 22787 4641 22799 4675
rect 22741 4635 22799 4641
rect 1854 4604 1860 4616
rect 1815 4576 1860 4604
rect 1854 4564 1860 4576
rect 1912 4564 1918 4616
rect 22094 4564 22100 4616
rect 22152 4604 22158 4616
rect 22756 4604 22784 4635
rect 22152 4576 22784 4604
rect 57057 4607 57115 4613
rect 22152 4564 22158 4576
rect 57057 4573 57069 4607
rect 57103 4604 57115 4607
rect 57514 4604 57520 4616
rect 57103 4576 57520 4604
rect 57103 4573 57115 4576
rect 57057 4567 57115 4573
rect 57514 4564 57520 4576
rect 57572 4564 57578 4616
rect 58342 4604 58348 4616
rect 58303 4576 58348 4604
rect 58342 4564 58348 4576
rect 58400 4564 58406 4616
rect 8294 4536 8300 4548
rect 7774 4508 8300 4536
rect 8294 4496 8300 4508
rect 8352 4536 8358 4548
rect 9398 4536 9404 4548
rect 8352 4508 9404 4536
rect 8352 4496 8358 4508
rect 9398 4496 9404 4508
rect 9456 4496 9462 4548
rect 14734 4496 14740 4548
rect 14792 4536 14798 4548
rect 56505 4539 56563 4545
rect 14792 4508 17618 4536
rect 14792 4496 14798 4508
rect 56505 4505 56517 4539
rect 56551 4536 56563 4539
rect 58360 4536 58388 4564
rect 56551 4508 58388 4536
rect 56551 4505 56563 4508
rect 56505 4499 56563 4505
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4428 1734 4480
rect 2774 4468 2780 4480
rect 2735 4440 2780 4468
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 20070 4468 20076 4480
rect 20031 4440 20076 4468
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 22189 4471 22247 4477
rect 22189 4437 22201 4471
rect 22235 4468 22247 4471
rect 22370 4468 22376 4480
rect 22235 4440 22376 4468
rect 22235 4437 22247 4440
rect 22189 4431 22247 4437
rect 22370 4428 22376 4440
rect 22428 4428 22434 4480
rect 22557 4471 22615 4477
rect 22557 4437 22569 4471
rect 22603 4468 22615 4471
rect 22646 4468 22652 4480
rect 22603 4440 22652 4468
rect 22603 4437 22615 4440
rect 22557 4431 22615 4437
rect 22646 4428 22652 4440
rect 22704 4428 22710 4480
rect 55953 4471 56011 4477
rect 55953 4437 55965 4471
rect 55999 4468 56011 4471
rect 56318 4468 56324 4480
rect 55999 4440 56324 4468
rect 55999 4437 56011 4440
rect 55953 4431 56011 4437
rect 56318 4428 56324 4440
rect 56376 4428 56382 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 18601 4267 18659 4273
rect 18601 4264 18613 4267
rect 16040 4236 18613 4264
rect 2317 4199 2375 4205
rect 2317 4165 2329 4199
rect 2363 4196 2375 4199
rect 3234 4196 3240 4208
rect 2363 4168 3240 4196
rect 2363 4165 2375 4168
rect 2317 4159 2375 4165
rect 3234 4156 3240 4168
rect 3292 4156 3298 4208
rect 4614 4156 4620 4208
rect 4672 4196 4678 4208
rect 5445 4199 5503 4205
rect 5445 4196 5457 4199
rect 4672 4168 5457 4196
rect 4672 4156 4678 4168
rect 5445 4165 5457 4168
rect 5491 4165 5503 4199
rect 5445 4159 5503 4165
rect 13906 4156 13912 4208
rect 13964 4196 13970 4208
rect 14734 4196 14740 4208
rect 13964 4168 14740 4196
rect 13964 4156 13970 4168
rect 14734 4156 14740 4168
rect 14792 4196 14798 4208
rect 16040 4205 16068 4236
rect 18601 4233 18613 4236
rect 18647 4233 18659 4267
rect 18601 4227 18659 4233
rect 18966 4224 18972 4276
rect 19024 4264 19030 4276
rect 19613 4267 19671 4273
rect 19613 4264 19625 4267
rect 19024 4236 19625 4264
rect 19024 4224 19030 4236
rect 19613 4233 19625 4236
rect 19659 4233 19671 4267
rect 19613 4227 19671 4233
rect 16025 4199 16083 4205
rect 14792 4168 14858 4196
rect 14792 4156 14798 4168
rect 16025 4165 16037 4199
rect 16071 4165 16083 4199
rect 16850 4196 16856 4208
rect 16025 4159 16083 4165
rect 16316 4168 16856 4196
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 16316 4137 16344 4168
rect 16850 4156 16856 4168
rect 16908 4156 16914 4208
rect 57440 4168 57652 4196
rect 16301 4131 16359 4137
rect 9088 4100 14596 4128
rect 9088 4088 9094 4100
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 2406 4060 2412 4072
rect 2271 4032 2412 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 2148 3992 2176 4023
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6362 4060 6368 4072
rect 5767 4032 6368 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6362 4020 6368 4032
rect 6420 4060 6426 4072
rect 11698 4060 11704 4072
rect 6420 4032 11704 4060
rect 6420 4020 6426 4032
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 14568 4069 14596 4100
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4128 18843 4131
rect 18874 4128 18880 4140
rect 18831 4100 18880 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 20622 4088 20628 4140
rect 20680 4128 20686 4140
rect 21453 4131 21511 4137
rect 21453 4128 21465 4131
rect 20680 4100 21465 4128
rect 20680 4088 20686 4100
rect 21453 4097 21465 4100
rect 21499 4128 21511 4131
rect 22186 4128 22192 4140
rect 21499 4100 22192 4128
rect 21499 4097 21511 4100
rect 21453 4091 21511 4097
rect 22186 4088 22192 4100
rect 22244 4088 22250 4140
rect 22370 4128 22376 4140
rect 22331 4100 22376 4128
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22738 4088 22744 4140
rect 22796 4128 22802 4140
rect 23017 4131 23075 4137
rect 23017 4128 23029 4131
rect 22796 4100 23029 4128
rect 22796 4088 22802 4100
rect 23017 4097 23029 4100
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 55861 4131 55919 4137
rect 55861 4097 55873 4131
rect 55907 4128 55919 4131
rect 55950 4128 55956 4140
rect 55907 4100 55956 4128
rect 55907 4097 55919 4100
rect 55861 4091 55919 4097
rect 55950 4088 55956 4100
rect 56008 4088 56014 4140
rect 56594 4128 56600 4140
rect 56555 4100 56600 4128
rect 56594 4088 56600 4100
rect 56652 4088 56658 4140
rect 57146 4088 57152 4140
rect 57204 4128 57210 4140
rect 57440 4128 57468 4168
rect 57204 4100 57468 4128
rect 57517 4131 57575 4137
rect 57204 4088 57210 4100
rect 57517 4097 57529 4131
rect 57563 4097 57575 4131
rect 57624 4128 57652 4168
rect 58253 4131 58311 4137
rect 58253 4128 58265 4131
rect 57624 4100 58265 4128
rect 57517 4091 57575 4097
rect 58253 4097 58265 4100
rect 58299 4097 58311 4131
rect 58253 4091 58311 4097
rect 14553 4063 14611 4069
rect 14553 4029 14565 4063
rect 14599 4060 14611 4063
rect 15930 4060 15936 4072
rect 14599 4032 15936 4060
rect 14599 4029 14611 4032
rect 14553 4023 14611 4029
rect 15930 4020 15936 4032
rect 15988 4020 15994 4072
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 19705 4063 19763 4069
rect 19705 4060 19717 4063
rect 18104 4032 19717 4060
rect 18104 4020 18110 4032
rect 19705 4029 19717 4032
rect 19751 4029 19763 4063
rect 19705 4023 19763 4029
rect 19794 4020 19800 4072
rect 19852 4060 19858 4072
rect 19852 4032 19897 4060
rect 19852 4020 19858 4032
rect 56502 4020 56508 4072
rect 56560 4060 56566 4072
rect 57532 4060 57560 4091
rect 56560 4032 57560 4060
rect 56560 4020 56566 4032
rect 2774 3992 2780 4004
rect 2148 3964 2780 3992
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 9490 3952 9496 4004
rect 9548 3992 9554 4004
rect 22833 3995 22891 4001
rect 22833 3992 22845 3995
rect 9548 3964 12434 3992
rect 9548 3952 9554 3964
rect 2222 3884 2228 3936
rect 2280 3924 2286 3936
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 2280 3896 2697 3924
rect 2280 3884 2286 3896
rect 2685 3893 2697 3896
rect 2731 3893 2743 3927
rect 3234 3924 3240 3936
rect 3195 3896 3240 3924
rect 2685 3887 2743 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 12250 3924 12256 3936
rect 12211 3896 12256 3924
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 12406 3924 12434 3964
rect 16224 3964 22845 3992
rect 16224 3924 16252 3964
rect 22833 3961 22845 3964
rect 22879 3961 22891 3995
rect 22833 3955 22891 3961
rect 50154 3952 50160 4004
rect 50212 3992 50218 4004
rect 57333 3995 57391 4001
rect 57333 3992 57345 3995
rect 50212 3964 57345 3992
rect 50212 3952 50218 3964
rect 57333 3961 57345 3964
rect 57379 3961 57391 3995
rect 57333 3955 57391 3961
rect 12406 3896 16252 3924
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16853 3927 16911 3933
rect 16853 3924 16865 3927
rect 16724 3896 16865 3924
rect 16724 3884 16730 3896
rect 16853 3893 16865 3896
rect 16899 3893 16911 3927
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 16853 3887 16911 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 19245 3927 19303 3933
rect 19245 3893 19257 3927
rect 19291 3924 19303 3927
rect 19334 3924 19340 3936
rect 19291 3896 19340 3924
rect 19291 3893 19303 3896
rect 19245 3887 19303 3893
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 20404 3896 20453 3924
rect 20404 3884 20410 3896
rect 20441 3893 20453 3896
rect 20487 3893 20499 3927
rect 20441 3887 20499 3893
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 22189 3927 22247 3933
rect 22189 3924 22201 3927
rect 20772 3896 22201 3924
rect 20772 3884 20778 3896
rect 22189 3893 22201 3896
rect 22235 3893 22247 3927
rect 22189 3887 22247 3893
rect 55309 3927 55367 3933
rect 55309 3893 55321 3927
rect 55355 3924 55367 3927
rect 57422 3924 57428 3936
rect 55355 3896 57428 3924
rect 55355 3893 55367 3896
rect 55309 3887 55367 3893
rect 57422 3884 57428 3896
rect 57480 3884 57486 3936
rect 58066 3924 58072 3936
rect 58027 3896 58072 3924
rect 58066 3884 58072 3896
rect 58124 3884 58130 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 3329 3723 3387 3729
rect 3329 3689 3341 3723
rect 3375 3720 3387 3723
rect 5641 3723 5699 3729
rect 5641 3720 5653 3723
rect 3375 3692 5653 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 5641 3689 5653 3692
rect 5687 3689 5699 3723
rect 5641 3683 5699 3689
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 10744 3692 11161 3720
rect 10744 3680 10750 3692
rect 11149 3689 11161 3692
rect 11195 3689 11207 3723
rect 13354 3720 13360 3732
rect 11149 3683 11207 3689
rect 12820 3692 13360 3720
rect 1854 3612 1860 3664
rect 1912 3652 1918 3664
rect 4157 3655 4215 3661
rect 4157 3652 4169 3655
rect 1912 3624 4169 3652
rect 1912 3612 1918 3624
rect 2240 3593 2268 3624
rect 4157 3621 4169 3624
rect 4203 3621 4215 3655
rect 4157 3615 4215 3621
rect 2133 3587 2191 3593
rect 2133 3553 2145 3587
rect 2179 3553 2191 3587
rect 2133 3547 2191 3553
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3553 2283 3587
rect 2774 3584 2780 3596
rect 2225 3547 2283 3553
rect 2332 3556 2780 3584
rect 2148 3516 2176 3547
rect 2332 3516 2360 3556
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 11606 3584 11612 3596
rect 3476 3556 11612 3584
rect 3476 3544 3482 3556
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 12820 3584 12848 3692
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 18874 3720 18880 3732
rect 14752 3692 18736 3720
rect 18835 3692 18880 3720
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 14752 3661 14780 3692
rect 14737 3655 14795 3661
rect 14737 3652 14749 3655
rect 13320 3624 14749 3652
rect 13320 3612 13326 3624
rect 14737 3621 14749 3624
rect 14783 3621 14795 3655
rect 18708 3652 18736 3692
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 22738 3720 22744 3732
rect 22699 3692 22744 3720
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 20346 3652 20352 3664
rect 18708 3624 20352 3652
rect 14737 3615 14795 3621
rect 20346 3612 20352 3624
rect 20404 3652 20410 3664
rect 20714 3652 20720 3664
rect 20404 3624 20720 3652
rect 20404 3612 20410 3624
rect 20714 3612 20720 3624
rect 20772 3612 20778 3664
rect 21358 3612 21364 3664
rect 21416 3652 21422 3664
rect 40129 3655 40187 3661
rect 21416 3624 22324 3652
rect 21416 3612 21422 3624
rect 12667 3556 12848 3584
rect 12897 3587 12955 3593
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 12897 3553 12909 3587
rect 12943 3584 12955 3587
rect 15654 3584 15660 3596
rect 12943 3556 15660 3584
rect 12943 3553 12955 3556
rect 12897 3547 12955 3553
rect 15654 3544 15660 3556
rect 15712 3584 15718 3596
rect 16485 3587 16543 3593
rect 16485 3584 16497 3587
rect 15712 3556 16497 3584
rect 15712 3544 15718 3556
rect 16485 3553 16497 3556
rect 16531 3584 16543 3587
rect 16850 3584 16856 3596
rect 16531 3556 16856 3584
rect 16531 3553 16543 3556
rect 16485 3547 16543 3553
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 18325 3587 18383 3593
rect 18325 3553 18337 3587
rect 18371 3584 18383 3587
rect 19794 3584 19800 3596
rect 18371 3556 19800 3584
rect 18371 3553 18383 3556
rect 18325 3547 18383 3553
rect 19794 3544 19800 3556
rect 19852 3584 19858 3596
rect 20901 3587 20959 3593
rect 20901 3584 20913 3587
rect 19852 3556 20913 3584
rect 19852 3544 19858 3556
rect 20901 3553 20913 3556
rect 20947 3553 20959 3587
rect 22094 3584 22100 3596
rect 22007 3556 22100 3584
rect 20901 3547 20959 3553
rect 2148 3488 2360 3516
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 2317 3451 2375 3457
rect 2317 3417 2329 3451
rect 2363 3448 2375 3451
rect 2958 3448 2964 3460
rect 2363 3420 2964 3448
rect 2363 3417 2375 3420
rect 2317 3411 2375 3417
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 2685 3383 2743 3389
rect 2685 3349 2697 3383
rect 2731 3380 2743 3383
rect 3160 3380 3188 3479
rect 5902 3476 5908 3528
rect 5960 3516 5966 3528
rect 6825 3519 6883 3525
rect 6825 3516 6837 3519
rect 5960 3488 6005 3516
rect 6104 3488 6837 3516
rect 5960 3476 5966 3488
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 6104 3448 6132 3488
rect 6825 3485 6837 3488
rect 6871 3516 6883 3519
rect 8294 3516 8300 3528
rect 6871 3488 8300 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 17681 3519 17739 3525
rect 14792 3488 15134 3516
rect 14792 3476 14798 3488
rect 17681 3485 17693 3519
rect 17727 3516 17739 3519
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 17727 3488 18521 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 18509 3485 18521 3488
rect 18555 3516 18567 3519
rect 19889 3519 19947 3525
rect 18555 3488 19840 3516
rect 18555 3485 18567 3488
rect 18509 3479 18567 3485
rect 5224 3420 6132 3448
rect 5224 3408 5230 3420
rect 6362 3408 6368 3460
rect 6420 3448 6426 3460
rect 6457 3451 6515 3457
rect 6457 3448 6469 3451
rect 6420 3420 6469 3448
rect 6420 3408 6426 3420
rect 6457 3417 6469 3420
rect 6503 3417 6515 3451
rect 6457 3411 6515 3417
rect 8018 3408 8024 3460
rect 8076 3448 8082 3460
rect 8076 3420 9260 3448
rect 8076 3408 8082 3420
rect 7282 3380 7288 3392
rect 2731 3352 3188 3380
rect 7243 3352 7288 3380
rect 2731 3349 2743 3352
rect 2685 3343 2743 3349
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 9125 3383 9183 3389
rect 9125 3380 9137 3383
rect 8996 3352 9137 3380
rect 8996 3340 9002 3352
rect 9125 3349 9137 3352
rect 9171 3349 9183 3383
rect 9232 3380 9260 3420
rect 12158 3408 12164 3460
rect 12216 3408 12222 3460
rect 16209 3451 16267 3457
rect 12406 3420 14964 3448
rect 12406 3380 12434 3420
rect 9232 3352 12434 3380
rect 14936 3380 14964 3420
rect 16209 3417 16221 3451
rect 16255 3448 16267 3451
rect 19812 3448 19840 3488
rect 19889 3485 19901 3519
rect 19935 3516 19947 3519
rect 20717 3519 20775 3525
rect 19935 3488 20392 3516
rect 19935 3485 19947 3488
rect 19889 3479 19947 3485
rect 20254 3448 20260 3460
rect 16255 3420 19748 3448
rect 19812 3420 20260 3448
rect 16255 3417 16267 3420
rect 16209 3411 16267 3417
rect 15838 3380 15844 3392
rect 14936 3352 15844 3380
rect 9125 3343 9183 3349
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 19720 3389 19748 3420
rect 20254 3408 20260 3420
rect 20312 3408 20318 3460
rect 20364 3389 20392 3488
rect 20717 3485 20729 3519
rect 20763 3516 20775 3519
rect 20806 3516 20812 3528
rect 20763 3488 20812 3516
rect 20763 3485 20775 3488
rect 20717 3479 20775 3485
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 20916 3516 20944 3547
rect 22066 3544 22100 3556
rect 22152 3544 22158 3596
rect 22296 3593 22324 3624
rect 40129 3621 40141 3655
rect 40175 3652 40187 3655
rect 53834 3652 53840 3664
rect 40175 3624 53840 3652
rect 40175 3621 40187 3624
rect 40129 3615 40187 3621
rect 22281 3587 22339 3593
rect 22281 3553 22293 3587
rect 22327 3553 22339 3587
rect 22281 3547 22339 3553
rect 22066 3516 22094 3544
rect 20916 3488 22094 3516
rect 22373 3519 22431 3525
rect 22373 3485 22385 3519
rect 22419 3516 22431 3519
rect 22462 3516 22468 3528
rect 22419 3488 22468 3516
rect 22419 3485 22431 3488
rect 22373 3479 22431 3485
rect 22462 3476 22468 3488
rect 22520 3476 22526 3528
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 22612 3488 23213 3516
rect 22612 3476 22618 3488
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 39117 3519 39175 3525
rect 39117 3485 39129 3519
rect 39163 3516 39175 3519
rect 40144 3516 40172 3615
rect 53834 3612 53840 3624
rect 53892 3612 53898 3664
rect 44818 3544 44824 3596
rect 44876 3584 44882 3596
rect 58618 3584 58624 3596
rect 44876 3556 58624 3584
rect 44876 3544 44882 3556
rect 58618 3544 58624 3556
rect 58676 3544 58682 3596
rect 39163 3488 40172 3516
rect 46477 3519 46535 3525
rect 39163 3485 39175 3488
rect 39117 3479 39175 3485
rect 46477 3485 46489 3519
rect 46523 3485 46535 3519
rect 48498 3516 48504 3528
rect 48459 3488 48504 3516
rect 46477 3479 46535 3485
rect 20824 3448 20852 3476
rect 21082 3448 21088 3460
rect 20824 3420 21088 3448
rect 21082 3408 21088 3420
rect 21140 3408 21146 3460
rect 46492 3448 46520 3479
rect 48498 3476 48504 3488
rect 48556 3516 48562 3528
rect 48961 3519 49019 3525
rect 48961 3516 48973 3519
rect 48556 3488 48973 3516
rect 48556 3476 48562 3488
rect 48961 3485 48973 3488
rect 49007 3485 49019 3519
rect 53098 3516 53104 3528
rect 53059 3488 53104 3516
rect 48961 3479 49019 3485
rect 53098 3476 53104 3488
rect 53156 3516 53162 3528
rect 53561 3519 53619 3525
rect 53561 3516 53573 3519
rect 53156 3488 53573 3516
rect 53156 3476 53162 3488
rect 53561 3485 53573 3488
rect 53607 3485 53619 3519
rect 53561 3479 53619 3485
rect 54573 3519 54631 3525
rect 54573 3485 54585 3519
rect 54619 3516 54631 3519
rect 54662 3516 54668 3528
rect 54619 3488 54668 3516
rect 54619 3485 54631 3488
rect 54573 3479 54631 3485
rect 54662 3476 54668 3488
rect 54720 3476 54726 3528
rect 55677 3519 55735 3525
rect 55677 3485 55689 3519
rect 55723 3516 55735 3519
rect 55950 3516 55956 3528
rect 55723 3488 55956 3516
rect 55723 3485 55735 3488
rect 55677 3479 55735 3485
rect 55950 3476 55956 3488
rect 56008 3476 56014 3528
rect 56505 3519 56563 3525
rect 56505 3485 56517 3519
rect 56551 3516 56563 3519
rect 56594 3516 56600 3528
rect 56551 3488 56600 3516
rect 56551 3485 56563 3488
rect 56505 3479 56563 3485
rect 56594 3476 56600 3488
rect 56652 3476 56658 3528
rect 57149 3519 57207 3525
rect 57149 3485 57161 3519
rect 57195 3516 57207 3519
rect 57238 3516 57244 3528
rect 57195 3488 57244 3516
rect 57195 3485 57207 3488
rect 57149 3479 57207 3485
rect 57238 3476 57244 3488
rect 57296 3476 57302 3528
rect 57606 3516 57612 3528
rect 57567 3488 57612 3516
rect 57606 3476 57612 3488
rect 57664 3476 57670 3528
rect 47029 3451 47087 3457
rect 47029 3448 47041 3451
rect 46492 3420 47041 3448
rect 47029 3417 47041 3420
rect 47075 3448 47087 3451
rect 55582 3448 55588 3460
rect 47075 3420 55588 3448
rect 47075 3417 47087 3420
rect 47029 3411 47087 3417
rect 55582 3408 55588 3420
rect 55640 3408 55646 3460
rect 17037 3383 17095 3389
rect 17037 3380 17049 3383
rect 15988 3352 17049 3380
rect 15988 3340 15994 3352
rect 17037 3349 17049 3352
rect 17083 3380 17095 3383
rect 18417 3383 18475 3389
rect 18417 3380 18429 3383
rect 17083 3352 18429 3380
rect 17083 3349 17095 3352
rect 17037 3343 17095 3349
rect 18417 3349 18429 3352
rect 18463 3349 18475 3383
rect 18417 3343 18475 3349
rect 19705 3383 19763 3389
rect 19705 3349 19717 3383
rect 19751 3349 19763 3383
rect 19705 3343 19763 3349
rect 20349 3383 20407 3389
rect 20349 3349 20361 3383
rect 20395 3349 20407 3383
rect 20349 3343 20407 3349
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 20809 3383 20867 3389
rect 20809 3380 20821 3383
rect 20772 3352 20821 3380
rect 20772 3340 20778 3352
rect 20809 3349 20821 3352
rect 20855 3349 20867 3383
rect 20809 3343 20867 3349
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 23385 3383 23443 3389
rect 23385 3380 23397 3383
rect 22152 3352 23397 3380
rect 22152 3340 22158 3352
rect 23385 3349 23397 3352
rect 23431 3349 23443 3383
rect 38930 3380 38936 3392
rect 38891 3352 38936 3380
rect 23385 3343 23443 3349
rect 38930 3340 38936 3352
rect 38988 3340 38994 3392
rect 45738 3340 45744 3392
rect 45796 3380 45802 3392
rect 46293 3383 46351 3389
rect 46293 3380 46305 3383
rect 45796 3352 46305 3380
rect 45796 3340 45802 3352
rect 46293 3349 46305 3352
rect 46339 3349 46351 3383
rect 48314 3380 48320 3392
rect 48275 3352 48320 3380
rect 46293 3343 46351 3349
rect 48314 3340 48320 3352
rect 48372 3340 48378 3392
rect 52914 3380 52920 3392
rect 52875 3352 52920 3380
rect 52914 3340 52920 3352
rect 52972 3340 52978 3392
rect 54386 3380 54392 3392
rect 54347 3352 54392 3380
rect 54386 3340 54392 3352
rect 54444 3340 54450 3392
rect 55490 3380 55496 3392
rect 55451 3352 55496 3380
rect 55490 3340 55496 3352
rect 55548 3340 55554 3392
rect 55766 3340 55772 3392
rect 55824 3380 55830 3392
rect 56321 3383 56379 3389
rect 56321 3380 56333 3383
rect 55824 3352 56333 3380
rect 55824 3340 55830 3352
rect 56321 3349 56333 3352
rect 56367 3349 56379 3383
rect 56962 3380 56968 3392
rect 56923 3352 56968 3380
rect 56321 3343 56379 3349
rect 56962 3340 56968 3352
rect 57020 3340 57026 3392
rect 57790 3380 57796 3392
rect 57751 3352 57796 3380
rect 57790 3340 57796 3352
rect 57848 3340 57854 3392
rect 58342 3380 58348 3392
rect 58303 3352 58348 3380
rect 58342 3340 58348 3352
rect 58400 3340 58406 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 2464 3148 4077 3176
rect 2464 3136 2470 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 4890 3176 4896 3188
rect 4065 3139 4123 3145
rect 4264 3148 4896 3176
rect 2774 3068 2780 3120
rect 2832 3108 2838 3120
rect 3513 3111 3571 3117
rect 3513 3108 3525 3111
rect 2832 3080 3525 3108
rect 2832 3068 2838 3080
rect 3513 3077 3525 3080
rect 3559 3077 3571 3111
rect 3513 3071 3571 3077
rect 2222 3040 2228 3052
rect 2183 3012 2228 3040
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 2958 3040 2964 3052
rect 2919 3012 2964 3040
rect 2958 3000 2964 3012
rect 3016 3040 3022 3052
rect 4264 3040 4292 3148
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 5166 3136 5172 3188
rect 5224 3136 5230 3188
rect 6362 3136 6368 3188
rect 6420 3176 6426 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6420 3148 6561 3176
rect 6420 3136 6426 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 8018 3176 8024 3188
rect 7979 3148 8024 3176
rect 6549 3139 6607 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 11698 3176 11704 3188
rect 11659 3148 11704 3176
rect 11698 3136 11704 3148
rect 11756 3176 11762 3188
rect 19153 3179 19211 3185
rect 19153 3176 19165 3179
rect 11756 3148 12434 3176
rect 11756 3136 11762 3148
rect 5184 3108 5212 3136
rect 9490 3108 9496 3120
rect 5106 3080 5212 3108
rect 9451 3080 9496 3108
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 12158 3068 12164 3120
rect 12216 3108 12222 3120
rect 12253 3111 12311 3117
rect 12253 3108 12265 3111
rect 12216 3080 12265 3108
rect 12216 3068 12222 3080
rect 12253 3077 12265 3080
rect 12299 3077 12311 3111
rect 12406 3108 12434 3148
rect 15396 3148 19165 3176
rect 12621 3111 12679 3117
rect 12621 3108 12633 3111
rect 12406 3080 12633 3108
rect 12253 3071 12311 3077
rect 12621 3077 12633 3080
rect 12667 3077 12679 3111
rect 12621 3071 12679 3077
rect 3016 3012 4292 3040
rect 5813 3043 5871 3049
rect 3016 3000 3022 3012
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5902 3040 5908 3052
rect 5859 3012 5908 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 8386 3000 8392 3052
rect 8444 3000 8450 3052
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 10318 3040 10324 3052
rect 9815 3012 10324 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 12268 3040 12296 3071
rect 14734 3068 14740 3120
rect 14792 3068 14798 3120
rect 15396 3117 15424 3148
rect 19153 3145 19165 3148
rect 19199 3145 19211 3179
rect 22554 3176 22560 3188
rect 22515 3148 22560 3176
rect 19153 3139 19211 3145
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 23934 3136 23940 3188
rect 23992 3176 23998 3188
rect 27249 3179 27307 3185
rect 27249 3176 27261 3179
rect 23992 3148 27261 3176
rect 23992 3136 23998 3148
rect 27249 3145 27261 3148
rect 27295 3145 27307 3179
rect 28718 3176 28724 3188
rect 28679 3148 28724 3176
rect 27249 3139 27307 3145
rect 15381 3111 15439 3117
rect 15381 3077 15393 3111
rect 15427 3077 15439 3111
rect 15381 3071 15439 3077
rect 15838 3068 15844 3120
rect 15896 3108 15902 3120
rect 21358 3108 21364 3120
rect 15896 3080 21364 3108
rect 15896 3068 15902 3080
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 13906 3040 13912 3052
rect 12268 3012 13912 3040
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 18046 3040 18052 3052
rect 15712 3012 15757 3040
rect 16224 3012 18052 3040
rect 15712 3000 15718 3012
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 2424 2944 5549 2972
rect 2424 2913 2452 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 16224 2972 16252 3012
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3040 18199 3043
rect 18966 3040 18972 3052
rect 18187 3012 18972 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 19334 3040 19340 3052
rect 19295 3012 19340 3040
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 20070 3040 20076 3052
rect 20031 3012 20076 3040
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 20349 3043 20407 3049
rect 20349 3009 20361 3043
rect 20395 3040 20407 3043
rect 20438 3040 20444 3052
rect 20395 3012 20444 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 22189 3043 22247 3049
rect 22189 3040 22201 3043
rect 20680 3012 22201 3040
rect 20680 3000 20686 3012
rect 22189 3009 22201 3012
rect 22235 3009 22247 3043
rect 22370 3040 22376 3052
rect 22331 3012 22376 3040
rect 22189 3003 22247 3009
rect 22370 3000 22376 3012
rect 22428 3040 22434 3052
rect 23017 3043 23075 3049
rect 23017 3040 23029 3043
rect 22428 3012 23029 3040
rect 22428 3000 22434 3012
rect 23017 3009 23029 3012
rect 23063 3009 23075 3043
rect 27264 3040 27292 3139
rect 28718 3136 28724 3148
rect 28776 3136 28782 3188
rect 29822 3176 29828 3188
rect 29783 3148 29828 3176
rect 29822 3136 29828 3148
rect 29880 3136 29886 3188
rect 30926 3176 30932 3188
rect 30887 3148 30932 3176
rect 30926 3136 30932 3148
rect 30984 3136 30990 3188
rect 33134 3176 33140 3188
rect 33095 3148 33140 3176
rect 33134 3136 33140 3148
rect 33192 3136 33198 3188
rect 42978 3176 42984 3188
rect 42939 3148 42984 3176
rect 42978 3136 42984 3148
rect 43036 3136 43042 3188
rect 43714 3176 43720 3188
rect 43675 3148 43720 3176
rect 43714 3136 43720 3148
rect 43772 3136 43778 3188
rect 44818 3176 44824 3188
rect 44779 3148 44824 3176
rect 44818 3136 44824 3148
rect 44876 3136 44882 3188
rect 51442 3176 51448 3188
rect 51403 3148 51448 3176
rect 51442 3136 51448 3148
rect 51500 3136 51506 3188
rect 54662 3176 54668 3188
rect 54623 3148 54668 3176
rect 54662 3136 54668 3148
rect 54720 3136 54726 3188
rect 55858 3176 55864 3188
rect 55819 3148 55864 3176
rect 55858 3136 55864 3148
rect 55916 3136 55922 3188
rect 56505 3179 56563 3185
rect 56505 3145 56517 3179
rect 56551 3176 56563 3179
rect 56686 3176 56692 3188
rect 56551 3148 56692 3176
rect 56551 3145 56563 3148
rect 56505 3139 56563 3145
rect 56686 3136 56692 3148
rect 56744 3136 56750 3188
rect 30282 3068 30288 3120
rect 30340 3108 30346 3120
rect 32306 3108 32312 3120
rect 30340 3080 32312 3108
rect 30340 3068 30346 3080
rect 32306 3068 32312 3080
rect 32364 3068 32370 3120
rect 37734 3068 37740 3120
rect 37792 3108 37798 3120
rect 37921 3111 37979 3117
rect 37921 3108 37933 3111
rect 37792 3080 37933 3108
rect 37792 3068 37798 3080
rect 37921 3077 37933 3080
rect 37967 3108 37979 3111
rect 58342 3108 58348 3120
rect 37967 3080 54616 3108
rect 37967 3077 37979 3080
rect 37921 3071 37979 3077
rect 27801 3043 27859 3049
rect 27801 3040 27813 3043
rect 27264 3012 27813 3040
rect 23017 3003 23075 3009
rect 27801 3009 27813 3012
rect 27847 3009 27859 3043
rect 27801 3003 27859 3009
rect 5537 2935 5595 2941
rect 6886 2944 16252 2972
rect 16301 2975 16359 2981
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2873 2467 2907
rect 2409 2867 2467 2873
rect 2516 2876 3188 2904
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 2516 2836 2544 2876
rect 2004 2808 2544 2836
rect 3160 2836 3188 2876
rect 6886 2836 6914 2944
rect 13924 2913 13952 2944
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 17770 2972 17776 2984
rect 16347 2944 17776 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 17770 2932 17776 2944
rect 17828 2972 17834 2984
rect 17865 2975 17923 2981
rect 17865 2972 17877 2975
rect 17828 2944 17877 2972
rect 17828 2932 17834 2944
rect 17865 2941 17877 2944
rect 17911 2941 17923 2975
rect 17865 2935 17923 2941
rect 40310 2932 40316 2984
rect 40368 2972 40374 2984
rect 40497 2975 40555 2981
rect 40497 2972 40509 2975
rect 40368 2944 40509 2972
rect 40368 2932 40374 2944
rect 40497 2941 40509 2944
rect 40543 2972 40555 2975
rect 50154 2972 50160 2984
rect 40543 2944 50160 2972
rect 40543 2941 40555 2944
rect 40497 2935 40555 2941
rect 50154 2932 50160 2944
rect 50212 2932 50218 2984
rect 50614 2932 50620 2984
rect 50672 2972 50678 2984
rect 50801 2975 50859 2981
rect 50801 2972 50813 2975
rect 50672 2944 50813 2972
rect 50672 2932 50678 2944
rect 50801 2941 50813 2944
rect 50847 2972 50859 2975
rect 54478 2972 54484 2984
rect 50847 2944 54484 2972
rect 50847 2941 50859 2944
rect 50801 2935 50859 2941
rect 54478 2932 54484 2944
rect 54536 2932 54542 2984
rect 54588 2972 54616 3080
rect 56704 3080 58348 3108
rect 55401 3043 55459 3049
rect 55401 3009 55413 3043
rect 55447 3040 55459 3043
rect 56042 3040 56048 3052
rect 55447 3012 56048 3040
rect 55447 3009 55459 3012
rect 55401 3003 55459 3009
rect 56042 3000 56048 3012
rect 56100 3000 56106 3052
rect 56704 3049 56732 3080
rect 58342 3068 58348 3080
rect 58400 3068 58406 3120
rect 56689 3043 56747 3049
rect 56689 3009 56701 3043
rect 56735 3009 56747 3043
rect 57330 3040 57336 3052
rect 57291 3012 57336 3040
rect 56689 3003 56747 3009
rect 57330 3000 57336 3012
rect 57388 3000 57394 3052
rect 58250 3040 58256 3052
rect 58211 3012 58256 3040
rect 58250 3000 58256 3012
rect 58308 3000 58314 3052
rect 54588 2944 58112 2972
rect 13909 2907 13967 2913
rect 13909 2873 13921 2907
rect 13955 2873 13967 2907
rect 38654 2904 38660 2916
rect 38567 2876 38660 2904
rect 13909 2867 13967 2873
rect 38654 2864 38660 2876
rect 38712 2904 38718 2916
rect 56962 2904 56968 2916
rect 38712 2876 56968 2904
rect 38712 2864 38718 2876
rect 56962 2864 56968 2876
rect 57020 2864 57026 2916
rect 58084 2913 58112 2944
rect 58069 2907 58127 2913
rect 58069 2873 58081 2907
rect 58115 2873 58127 2907
rect 58069 2867 58127 2873
rect 3160 2808 6914 2836
rect 7469 2839 7527 2845
rect 2004 2796 2010 2808
rect 7469 2805 7481 2839
rect 7515 2836 7527 2839
rect 7834 2836 7840 2848
rect 7515 2808 7840 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 10100 2808 10241 2836
rect 10100 2796 10106 2808
rect 10229 2805 10241 2808
rect 10275 2805 10287 2839
rect 11146 2836 11152 2848
rect 11107 2808 11152 2836
rect 10229 2799 10287 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 13449 2839 13507 2845
rect 13449 2805 13461 2839
rect 13495 2836 13507 2839
rect 13814 2836 13820 2848
rect 13495 2808 13820 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 17405 2839 17463 2845
rect 17405 2805 17417 2839
rect 17451 2836 17463 2839
rect 18874 2836 18880 2848
rect 17451 2808 18880 2836
rect 17451 2805 17463 2808
rect 17405 2799 17463 2805
rect 18874 2796 18880 2808
rect 18932 2796 18938 2848
rect 23290 2796 23296 2848
rect 23348 2836 23354 2848
rect 23845 2839 23903 2845
rect 23845 2836 23857 2839
rect 23348 2808 23857 2836
rect 23348 2796 23354 2808
rect 23845 2805 23857 2808
rect 23891 2805 23903 2839
rect 24394 2836 24400 2848
rect 24355 2808 24400 2836
rect 23845 2799 23903 2805
rect 24394 2796 24400 2808
rect 24452 2796 24458 2848
rect 25498 2836 25504 2848
rect 25459 2808 25504 2836
rect 25498 2796 25504 2808
rect 25556 2796 25562 2848
rect 27706 2796 27712 2848
rect 27764 2836 27770 2848
rect 27985 2839 28043 2845
rect 27985 2836 27997 2839
rect 27764 2808 27997 2836
rect 27764 2796 27770 2808
rect 27985 2805 27997 2808
rect 28031 2805 28043 2839
rect 35986 2836 35992 2848
rect 35947 2808 35992 2836
rect 27985 2799 28043 2805
rect 35986 2796 35992 2808
rect 36044 2796 36050 2848
rect 54205 2839 54263 2845
rect 54205 2805 54217 2839
rect 54251 2836 54263 2839
rect 55950 2836 55956 2848
rect 54251 2808 55956 2836
rect 54251 2805 54263 2808
rect 54205 2799 54263 2805
rect 55950 2796 55956 2808
rect 56008 2796 56014 2848
rect 57146 2836 57152 2848
rect 57107 2808 57152 2836
rect 57146 2796 57152 2808
rect 57204 2796 57210 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 2593 2635 2651 2641
rect 2593 2601 2605 2635
rect 2639 2632 2651 2635
rect 4614 2632 4620 2644
rect 2639 2604 4620 2632
rect 2639 2601 2651 2604
rect 2593 2595 2651 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 4798 2632 4804 2644
rect 4759 2604 4804 2632
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 14642 2632 14648 2644
rect 14603 2604 14648 2632
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 15841 2635 15899 2641
rect 15841 2601 15853 2635
rect 15887 2632 15899 2635
rect 18690 2632 18696 2644
rect 15887 2604 18696 2632
rect 15887 2601 15899 2604
rect 15841 2595 15899 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 22462 2632 22468 2644
rect 22423 2604 22468 2632
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 24949 2635 25007 2641
rect 24949 2601 24961 2635
rect 24995 2632 25007 2635
rect 28902 2632 28908 2644
rect 24995 2604 28908 2632
rect 24995 2601 25007 2604
rect 24949 2595 25007 2601
rect 28902 2592 28908 2604
rect 28960 2592 28966 2644
rect 55398 2632 55404 2644
rect 39776 2604 55404 2632
rect 4890 2524 4896 2576
rect 4948 2564 4954 2576
rect 6825 2567 6883 2573
rect 6825 2564 6837 2567
rect 4948 2536 6837 2564
rect 4948 2524 4954 2536
rect 6825 2533 6837 2536
rect 6871 2533 6883 2567
rect 6825 2527 6883 2533
rect 17129 2567 17187 2573
rect 17129 2533 17141 2567
rect 17175 2564 17187 2567
rect 18230 2564 18236 2576
rect 17175 2536 18236 2564
rect 17175 2533 17187 2536
rect 17129 2527 17187 2533
rect 18230 2524 18236 2536
rect 18288 2524 18294 2576
rect 25777 2567 25835 2573
rect 25777 2533 25789 2567
rect 25823 2564 25835 2567
rect 39666 2564 39672 2576
rect 25823 2536 39672 2564
rect 25823 2533 25835 2536
rect 25777 2527 25835 2533
rect 39666 2524 39672 2536
rect 39724 2524 39730 2576
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 4028 2468 4752 2496
rect 4028 2456 4034 2468
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2314 2428 2320 2440
rect 1995 2400 2320 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2314 2388 2320 2400
rect 2372 2428 2378 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2372 2400 2421 2428
rect 2372 2388 2378 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4522 2428 4528 2440
rect 3467 2400 4528 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4522 2388 4528 2400
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4724 2428 4752 2468
rect 4908 2468 9413 2496
rect 4908 2428 4936 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 18874 2496 18880 2508
rect 18835 2468 18880 2496
rect 9401 2459 9459 2465
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19613 2499 19671 2505
rect 19613 2465 19625 2499
rect 19659 2496 19671 2499
rect 20625 2499 20683 2505
rect 20625 2496 20637 2499
rect 19659 2468 20637 2496
rect 19659 2465 19671 2468
rect 19613 2459 19671 2465
rect 20625 2465 20637 2468
rect 20671 2496 20683 2499
rect 21082 2496 21088 2508
rect 20671 2468 21088 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 21082 2456 21088 2468
rect 21140 2456 21146 2508
rect 22646 2456 22652 2508
rect 22704 2496 22710 2508
rect 23477 2499 23535 2505
rect 23477 2496 23489 2499
rect 22704 2468 23489 2496
rect 22704 2456 22710 2468
rect 23477 2465 23489 2468
rect 23523 2465 23535 2499
rect 23477 2459 23535 2465
rect 27985 2499 28043 2505
rect 27985 2465 27997 2499
rect 28031 2496 28043 2499
rect 29730 2496 29736 2508
rect 28031 2468 29736 2496
rect 28031 2465 28043 2468
rect 27985 2459 28043 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 36357 2499 36415 2505
rect 36357 2465 36369 2499
rect 36403 2496 36415 2499
rect 39776 2496 39804 2604
rect 55398 2592 55404 2604
rect 55456 2592 55462 2644
rect 56689 2635 56747 2641
rect 56689 2601 56701 2635
rect 56735 2632 56747 2635
rect 57606 2632 57612 2644
rect 56735 2604 57612 2632
rect 56735 2601 56747 2604
rect 56689 2595 56747 2601
rect 57606 2592 57612 2604
rect 57664 2592 57670 2644
rect 56134 2524 56140 2576
rect 56192 2564 56198 2576
rect 57333 2567 57391 2573
rect 57333 2564 57345 2567
rect 56192 2536 57345 2564
rect 56192 2524 56198 2536
rect 57333 2533 57345 2536
rect 57379 2533 57391 2567
rect 57333 2527 57391 2533
rect 57146 2496 57152 2508
rect 36403 2468 39804 2496
rect 41156 2468 42012 2496
rect 36403 2465 36415 2468
rect 36357 2459 36415 2465
rect 4724 2400 4936 2428
rect 4617 2391 4675 2397
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 5721 2431 5779 2437
rect 5721 2428 5733 2431
rect 5684 2400 5733 2428
rect 5684 2388 5690 2400
rect 5721 2397 5733 2400
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6972 2400 7021 2428
rect 6972 2388 6978 2400
rect 7009 2397 7021 2400
rect 7055 2428 7067 2431
rect 7282 2428 7288 2440
rect 7055 2400 7288 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 7392 2400 10149 2428
rect 4157 2363 4215 2369
rect 4157 2329 4169 2363
rect 4203 2360 4215 2363
rect 5644 2360 5672 2388
rect 7392 2360 7420 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12216 2400 12357 2428
rect 12216 2388 12222 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12492 2400 12541 2428
rect 12492 2388 12498 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 13354 2388 13360 2440
rect 13412 2428 13418 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 13412 2400 13461 2428
rect 13412 2388 13418 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14458 2428 14464 2440
rect 13872 2400 14464 2428
rect 13872 2388 13878 2400
rect 14458 2388 14464 2400
rect 14516 2428 14522 2440
rect 14737 2431 14795 2437
rect 14737 2428 14749 2431
rect 14516 2400 14749 2428
rect 14516 2388 14522 2400
rect 14737 2397 14749 2400
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15620 2400 15761 2428
rect 15620 2388 15626 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 18601 2431 18659 2437
rect 18601 2397 18613 2431
rect 18647 2428 18659 2431
rect 19426 2428 19432 2440
rect 18647 2400 19432 2428
rect 18647 2397 18659 2400
rect 18601 2391 18659 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2428 20959 2431
rect 20990 2428 20996 2440
rect 20947 2400 20996 2428
rect 20947 2397 20959 2400
rect 20901 2391 20959 2397
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 22281 2431 22339 2437
rect 22281 2397 22293 2431
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2428 23259 2431
rect 23290 2428 23296 2440
rect 23247 2400 23296 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 4203 2332 5672 2360
rect 5736 2332 7420 2360
rect 4203 2329 4215 2332
rect 4157 2323 4215 2329
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 5736 2292 5764 2332
rect 7834 2320 7840 2372
rect 7892 2360 7898 2372
rect 8021 2363 8079 2369
rect 8021 2360 8033 2363
rect 7892 2332 8033 2360
rect 7892 2320 7898 2332
rect 8021 2329 8033 2332
rect 8067 2329 8079 2363
rect 8021 2323 8079 2329
rect 8938 2320 8944 2372
rect 8996 2360 9002 2372
rect 9217 2363 9275 2369
rect 9217 2360 9229 2363
rect 8996 2332 9229 2360
rect 8996 2320 9002 2332
rect 9217 2329 9229 2332
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 10042 2320 10048 2372
rect 10100 2360 10106 2372
rect 10321 2363 10379 2369
rect 10321 2360 10333 2363
rect 10100 2332 10333 2360
rect 10100 2320 10106 2332
rect 10321 2329 10333 2332
rect 10367 2329 10379 2363
rect 10321 2323 10379 2329
rect 11057 2363 11115 2369
rect 11057 2329 11069 2363
rect 11103 2360 11115 2363
rect 11146 2360 11152 2372
rect 11103 2332 11152 2360
rect 11103 2329 11115 2332
rect 11057 2323 11115 2329
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 13372 2360 13400 2388
rect 12406 2332 13400 2360
rect 5902 2292 5908 2304
rect 4120 2264 5764 2292
rect 5863 2264 5908 2292
rect 4120 2252 4126 2264
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 8110 2292 8116 2304
rect 8071 2264 8116 2292
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 10962 2292 10968 2304
rect 10923 2264 10968 2292
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2292 11943 2295
rect 12406 2292 12434 2332
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 16945 2363 17003 2369
rect 16945 2360 16957 2363
rect 16724 2332 16957 2360
rect 16724 2320 16730 2332
rect 16945 2329 16957 2332
rect 16991 2329 17003 2363
rect 16945 2323 17003 2329
rect 20165 2363 20223 2369
rect 20165 2329 20177 2363
rect 20211 2360 20223 2363
rect 22186 2360 22192 2372
rect 20211 2332 22192 2360
rect 20211 2329 20223 2332
rect 20165 2323 20223 2329
rect 22186 2320 22192 2332
rect 22244 2360 22250 2372
rect 22296 2360 22324 2391
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 25498 2388 25504 2440
rect 25556 2428 25562 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 25556 2400 25605 2428
rect 25556 2388 25562 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 28718 2388 28724 2440
rect 28776 2428 28782 2440
rect 28905 2431 28963 2437
rect 28905 2428 28917 2431
rect 28776 2400 28917 2428
rect 28776 2388 28782 2400
rect 28905 2397 28917 2400
rect 28951 2397 28963 2431
rect 28905 2391 28963 2397
rect 29822 2388 29828 2440
rect 29880 2428 29886 2440
rect 30009 2431 30067 2437
rect 30009 2428 30021 2431
rect 29880 2400 30021 2428
rect 29880 2388 29886 2400
rect 30009 2397 30021 2400
rect 30055 2397 30067 2431
rect 30009 2391 30067 2397
rect 30926 2388 30932 2440
rect 30984 2428 30990 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 30984 2400 31125 2428
rect 30984 2388 30990 2400
rect 31113 2397 31125 2400
rect 31159 2397 31171 2431
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 31113 2391 31171 2397
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33321 2431 33379 2437
rect 33321 2428 33333 2431
rect 33192 2400 33333 2428
rect 33192 2388 33198 2400
rect 33321 2397 33333 2400
rect 33367 2397 33379 2431
rect 34977 2431 35035 2437
rect 34977 2428 34989 2431
rect 33321 2391 33379 2397
rect 34348 2400 34989 2428
rect 22244 2332 22324 2360
rect 22244 2320 22250 2332
rect 24394 2320 24400 2372
rect 24452 2360 24458 2372
rect 24673 2363 24731 2369
rect 24673 2360 24685 2363
rect 24452 2332 24685 2360
rect 24452 2320 24458 2332
rect 24673 2329 24685 2332
rect 24719 2329 24731 2363
rect 24673 2323 24731 2329
rect 27157 2363 27215 2369
rect 27157 2329 27169 2363
rect 27203 2329 27215 2363
rect 27157 2323 27215 2329
rect 13630 2292 13636 2304
rect 11931 2264 12434 2292
rect 13591 2264 13636 2292
rect 11931 2261 11943 2264
rect 11885 2255 11943 2261
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 26602 2292 26608 2304
rect 26563 2264 26608 2292
rect 26602 2252 26608 2264
rect 26660 2292 26666 2304
rect 27172 2292 27200 2323
rect 34348 2304 34376 2400
rect 34977 2397 34989 2400
rect 35023 2397 35035 2431
rect 34977 2391 35035 2397
rect 35986 2388 35992 2440
rect 36044 2428 36050 2440
rect 36081 2431 36139 2437
rect 36081 2428 36093 2431
rect 36044 2400 36093 2428
rect 36044 2388 36050 2400
rect 36081 2397 36093 2400
rect 36127 2397 36139 2431
rect 37734 2428 37740 2440
rect 37695 2400 37740 2428
rect 36081 2391 36139 2397
rect 37734 2388 37740 2400
rect 37792 2388 37798 2440
rect 38473 2431 38531 2437
rect 38473 2397 38485 2431
rect 38519 2428 38531 2431
rect 38654 2428 38660 2440
rect 38519 2400 38660 2428
rect 38519 2397 38531 2400
rect 38473 2391 38531 2397
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 38930 2428 38936 2440
rect 38891 2400 38936 2428
rect 38930 2388 38936 2400
rect 38988 2388 38994 2440
rect 40310 2428 40316 2440
rect 40271 2400 40316 2428
rect 40310 2388 40316 2400
rect 40368 2388 40374 2440
rect 35529 2363 35587 2369
rect 35529 2329 35541 2363
rect 35575 2360 35587 2363
rect 41156 2360 41184 2468
rect 41325 2431 41383 2437
rect 41325 2397 41337 2431
rect 41371 2428 41383 2431
rect 41371 2400 41920 2428
rect 41371 2397 41383 2400
rect 41325 2391 41383 2397
rect 35575 2332 41184 2360
rect 35575 2329 35587 2332
rect 35529 2323 35587 2329
rect 41892 2304 41920 2400
rect 41984 2360 42012 2468
rect 46860 2468 57152 2496
rect 42889 2431 42947 2437
rect 42889 2397 42901 2431
rect 42935 2428 42947 2431
rect 42978 2428 42984 2440
rect 42935 2400 42984 2428
rect 42935 2397 42947 2400
rect 42889 2391 42947 2397
rect 42978 2388 42984 2400
rect 43036 2388 43042 2440
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43714 2428 43720 2440
rect 43671 2400 43720 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43714 2388 43720 2400
rect 43772 2388 43778 2440
rect 44637 2431 44695 2437
rect 44637 2397 44649 2431
rect 44683 2428 44695 2431
rect 44818 2428 44824 2440
rect 44683 2400 44824 2428
rect 44683 2397 44695 2400
rect 44637 2391 44695 2397
rect 44818 2388 44824 2400
rect 44876 2388 44882 2440
rect 45738 2428 45744 2440
rect 45699 2400 45744 2428
rect 45738 2388 45744 2400
rect 45796 2388 45802 2440
rect 46860 2437 46888 2468
rect 57146 2456 57152 2468
rect 57204 2456 57210 2508
rect 46845 2431 46903 2437
rect 46845 2397 46857 2431
rect 46891 2397 46903 2431
rect 46845 2391 46903 2397
rect 48041 2431 48099 2437
rect 48041 2397 48053 2431
rect 48087 2428 48099 2431
rect 48314 2428 48320 2440
rect 48087 2400 48320 2428
rect 48087 2397 48099 2400
rect 48041 2391 48099 2397
rect 48314 2388 48320 2400
rect 48372 2388 48378 2440
rect 49050 2428 49056 2440
rect 49011 2400 49056 2428
rect 49050 2388 49056 2400
rect 49108 2428 49114 2440
rect 49513 2431 49571 2437
rect 49513 2428 49525 2431
rect 49108 2400 49525 2428
rect 49108 2388 49114 2400
rect 49513 2397 49525 2400
rect 49559 2397 49571 2431
rect 50614 2428 50620 2440
rect 50575 2400 50620 2428
rect 49513 2391 49571 2397
rect 50614 2388 50620 2400
rect 50672 2388 50678 2440
rect 51353 2431 51411 2437
rect 51353 2397 51365 2431
rect 51399 2428 51411 2431
rect 51442 2428 51448 2440
rect 51399 2400 51448 2428
rect 51399 2397 51411 2400
rect 51353 2391 51411 2397
rect 51442 2388 51448 2400
rect 51500 2388 51506 2440
rect 52365 2431 52423 2437
rect 52365 2397 52377 2431
rect 52411 2428 52423 2431
rect 52914 2428 52920 2440
rect 52411 2400 52920 2428
rect 52411 2397 52423 2400
rect 52365 2391 52423 2397
rect 52914 2388 52920 2400
rect 52972 2388 52978 2440
rect 53469 2431 53527 2437
rect 53469 2397 53481 2431
rect 53515 2428 53527 2431
rect 54386 2428 54392 2440
rect 53515 2400 54392 2428
rect 53515 2397 53527 2400
rect 53469 2391 53527 2397
rect 54386 2388 54392 2400
rect 54444 2388 54450 2440
rect 54573 2431 54631 2437
rect 54573 2397 54585 2431
rect 54619 2428 54631 2431
rect 55490 2428 55496 2440
rect 54619 2400 55496 2428
rect 54619 2397 54631 2400
rect 54573 2391 54631 2397
rect 55490 2388 55496 2400
rect 55548 2388 55554 2440
rect 55766 2428 55772 2440
rect 55727 2400 55772 2428
rect 55766 2388 55772 2400
rect 55824 2388 55830 2440
rect 55950 2388 55956 2440
rect 56008 2428 56014 2440
rect 56410 2428 56416 2440
rect 56008 2400 56416 2428
rect 56008 2388 56014 2400
rect 56410 2388 56416 2400
rect 56468 2428 56474 2440
rect 56505 2431 56563 2437
rect 56505 2428 56517 2431
rect 56468 2400 56517 2428
rect 56468 2388 56474 2400
rect 56505 2397 56517 2400
rect 56551 2397 56563 2431
rect 56505 2391 56563 2397
rect 57517 2431 57575 2437
rect 57517 2397 57529 2431
rect 57563 2397 57575 2431
rect 57517 2391 57575 2397
rect 56226 2360 56232 2372
rect 41984 2332 56232 2360
rect 56226 2320 56232 2332
rect 56284 2320 56290 2372
rect 56318 2320 56324 2372
rect 56376 2360 56382 2372
rect 57532 2360 57560 2391
rect 57790 2388 57796 2440
rect 57848 2428 57854 2440
rect 58069 2431 58127 2437
rect 58069 2428 58081 2431
rect 57848 2400 58081 2428
rect 57848 2388 57854 2400
rect 58069 2397 58081 2400
rect 58115 2397 58127 2431
rect 58069 2391 58127 2397
rect 56376 2332 57560 2360
rect 56376 2320 56382 2332
rect 26660 2264 27200 2292
rect 26660 2252 26666 2264
rect 28810 2252 28816 2304
rect 28868 2292 28874 2304
rect 29089 2295 29147 2301
rect 29089 2292 29101 2295
rect 28868 2264 29101 2292
rect 28868 2252 28874 2264
rect 29089 2261 29101 2264
rect 29135 2261 29147 2295
rect 29089 2255 29147 2261
rect 29914 2252 29920 2304
rect 29972 2292 29978 2304
rect 30193 2295 30251 2301
rect 30193 2292 30205 2295
rect 29972 2264 30205 2292
rect 29972 2252 29978 2264
rect 30193 2261 30205 2264
rect 30239 2261 30251 2295
rect 30193 2255 30251 2261
rect 31018 2252 31024 2304
rect 31076 2292 31082 2304
rect 31297 2295 31355 2301
rect 31297 2292 31309 2295
rect 31076 2264 31309 2292
rect 31076 2252 31082 2264
rect 31297 2261 31309 2264
rect 31343 2261 31355 2295
rect 31297 2255 31355 2261
rect 32122 2252 32128 2304
rect 32180 2292 32186 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 32180 2264 32505 2292
rect 32180 2252 32186 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 33226 2252 33232 2304
rect 33284 2292 33290 2304
rect 33505 2295 33563 2301
rect 33505 2292 33517 2295
rect 33284 2264 33517 2292
rect 33284 2252 33290 2264
rect 33505 2261 33517 2264
rect 33551 2261 33563 2295
rect 34330 2292 34336 2304
rect 34291 2264 34336 2292
rect 33505 2255 33563 2261
rect 34330 2252 34336 2264
rect 34388 2252 34394 2304
rect 36538 2252 36544 2304
rect 36596 2292 36602 2304
rect 37553 2295 37611 2301
rect 37553 2292 37565 2295
rect 36596 2264 37565 2292
rect 36596 2252 36602 2264
rect 37553 2261 37565 2264
rect 37599 2261 37611 2295
rect 37553 2255 37611 2261
rect 37642 2252 37648 2304
rect 37700 2292 37706 2304
rect 38289 2295 38347 2301
rect 38289 2292 38301 2295
rect 37700 2264 38301 2292
rect 37700 2252 37706 2264
rect 38289 2261 38301 2264
rect 38335 2261 38347 2295
rect 38289 2255 38347 2261
rect 38746 2252 38752 2304
rect 38804 2292 38810 2304
rect 39117 2295 39175 2301
rect 39117 2292 39129 2295
rect 38804 2264 39129 2292
rect 38804 2252 38810 2264
rect 39117 2261 39129 2264
rect 39163 2261 39175 2295
rect 39117 2255 39175 2261
rect 39850 2252 39856 2304
rect 39908 2292 39914 2304
rect 40129 2295 40187 2301
rect 40129 2292 40141 2295
rect 39908 2264 40141 2292
rect 39908 2252 39914 2264
rect 40129 2261 40141 2264
rect 40175 2261 40187 2295
rect 40129 2255 40187 2261
rect 40954 2252 40960 2304
rect 41012 2292 41018 2304
rect 41141 2295 41199 2301
rect 41141 2292 41153 2295
rect 41012 2264 41153 2292
rect 41012 2252 41018 2264
rect 41141 2261 41153 2264
rect 41187 2261 41199 2295
rect 41874 2292 41880 2304
rect 41835 2264 41880 2292
rect 41141 2255 41199 2261
rect 41874 2252 41880 2264
rect 41932 2252 41938 2304
rect 42058 2252 42064 2304
rect 42116 2292 42122 2304
rect 42705 2295 42763 2301
rect 42705 2292 42717 2295
rect 42116 2264 42717 2292
rect 42116 2252 42122 2264
rect 42705 2261 42717 2264
rect 42751 2261 42763 2295
rect 42705 2255 42763 2261
rect 43162 2252 43168 2304
rect 43220 2292 43226 2304
rect 43441 2295 43499 2301
rect 43441 2292 43453 2295
rect 43220 2264 43453 2292
rect 43220 2252 43226 2264
rect 43441 2261 43453 2264
rect 43487 2261 43499 2295
rect 43441 2255 43499 2261
rect 44266 2252 44272 2304
rect 44324 2292 44330 2304
rect 44453 2295 44511 2301
rect 44453 2292 44465 2295
rect 44324 2264 44465 2292
rect 44324 2252 44330 2264
rect 44453 2261 44465 2264
rect 44499 2261 44511 2295
rect 44453 2255 44511 2261
rect 45370 2252 45376 2304
rect 45428 2292 45434 2304
rect 45557 2295 45615 2301
rect 45557 2292 45569 2295
rect 45428 2264 45569 2292
rect 45428 2252 45434 2264
rect 45557 2261 45569 2264
rect 45603 2261 45615 2295
rect 45557 2255 45615 2261
rect 46474 2252 46480 2304
rect 46532 2292 46538 2304
rect 46661 2295 46719 2301
rect 46661 2292 46673 2295
rect 46532 2264 46673 2292
rect 46532 2252 46538 2264
rect 46661 2261 46673 2264
rect 46707 2261 46719 2295
rect 46661 2255 46719 2261
rect 47578 2252 47584 2304
rect 47636 2292 47642 2304
rect 47857 2295 47915 2301
rect 47857 2292 47869 2295
rect 47636 2264 47869 2292
rect 47636 2252 47642 2264
rect 47857 2261 47869 2264
rect 47903 2261 47915 2295
rect 47857 2255 47915 2261
rect 48682 2252 48688 2304
rect 48740 2292 48746 2304
rect 48869 2295 48927 2301
rect 48869 2292 48881 2295
rect 48740 2264 48881 2292
rect 48740 2252 48746 2264
rect 48869 2261 48881 2264
rect 48915 2261 48927 2295
rect 48869 2255 48927 2261
rect 49786 2252 49792 2304
rect 49844 2292 49850 2304
rect 50433 2295 50491 2301
rect 50433 2292 50445 2295
rect 49844 2264 50445 2292
rect 49844 2252 49850 2264
rect 50433 2261 50445 2264
rect 50479 2261 50491 2295
rect 50433 2255 50491 2261
rect 50890 2252 50896 2304
rect 50948 2292 50954 2304
rect 51169 2295 51227 2301
rect 51169 2292 51181 2295
rect 50948 2264 51181 2292
rect 50948 2252 50954 2264
rect 51169 2261 51181 2264
rect 51215 2261 51227 2295
rect 51169 2255 51227 2261
rect 51994 2252 52000 2304
rect 52052 2292 52058 2304
rect 52181 2295 52239 2301
rect 52181 2292 52193 2295
rect 52052 2264 52193 2292
rect 52052 2252 52058 2264
rect 52181 2261 52193 2264
rect 52227 2261 52239 2295
rect 52181 2255 52239 2261
rect 53098 2252 53104 2304
rect 53156 2292 53162 2304
rect 53285 2295 53343 2301
rect 53285 2292 53297 2295
rect 53156 2264 53297 2292
rect 53156 2252 53162 2264
rect 53285 2261 53297 2264
rect 53331 2261 53343 2295
rect 53285 2255 53343 2261
rect 54202 2252 54208 2304
rect 54260 2292 54266 2304
rect 54389 2295 54447 2301
rect 54389 2292 54401 2295
rect 54260 2264 54401 2292
rect 54260 2252 54266 2264
rect 54389 2261 54401 2264
rect 54435 2261 54447 2295
rect 54389 2255 54447 2261
rect 55306 2252 55312 2304
rect 55364 2292 55370 2304
rect 55585 2295 55643 2301
rect 55585 2292 55597 2295
rect 55364 2264 55597 2292
rect 55364 2252 55370 2264
rect 55585 2261 55597 2264
rect 55631 2261 55643 2295
rect 55585 2255 55643 2261
rect 57514 2252 57520 2304
rect 57572 2292 57578 2304
rect 58253 2295 58311 2301
rect 58253 2292 58265 2295
rect 57572 2264 58265 2292
rect 57572 2252 57578 2264
rect 58253 2261 58265 2264
rect 58299 2261 58311 2295
rect 58253 2255 58311 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 4798 2048 4804 2100
rect 4856 2088 4862 2100
rect 22370 2088 22376 2100
rect 4856 2060 22376 2088
rect 4856 2048 4862 2060
rect 22370 2048 22376 2060
rect 22428 2048 22434 2100
rect 41874 2048 41880 2100
rect 41932 2088 41938 2100
rect 58066 2088 58072 2100
rect 41932 2060 58072 2088
rect 41932 2048 41938 2060
rect 58066 2048 58072 2060
rect 58124 2048 58130 2100
rect 3234 1980 3240 2032
rect 3292 2020 3298 2032
rect 8110 2020 8116 2032
rect 3292 1992 8116 2020
rect 3292 1980 3298 1992
rect 8110 1980 8116 1992
rect 8168 1980 8174 2032
rect 5902 1912 5908 1964
rect 5960 1952 5966 1964
rect 20622 1952 20628 1964
rect 5960 1924 20628 1952
rect 5960 1912 5966 1924
rect 20622 1912 20628 1924
rect 20680 1912 20686 1964
rect 3326 1844 3332 1896
rect 3384 1884 3390 1896
rect 12158 1884 12164 1896
rect 3384 1856 12164 1884
rect 3384 1844 3390 1856
rect 12158 1844 12164 1856
rect 12216 1844 12222 1896
rect 6178 1776 6184 1828
rect 6236 1816 6242 1828
rect 13630 1816 13636 1828
rect 6236 1788 13636 1816
rect 6236 1776 6242 1788
rect 13630 1776 13636 1788
rect 13688 1776 13694 1828
rect 3510 1708 3516 1760
rect 3568 1748 3574 1760
rect 10962 1748 10968 1760
rect 3568 1720 10968 1748
rect 3568 1708 3574 1720
rect 10962 1708 10968 1720
rect 11020 1708 11026 1760
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 11428 57536 11480 57588
rect 13820 57536 13872 57588
rect 16212 57579 16264 57588
rect 16212 57545 16221 57579
rect 16221 57545 16255 57579
rect 16255 57545 16264 57579
rect 16212 57536 16264 57545
rect 20720 57536 20772 57588
rect 20904 57468 20956 57520
rect 25780 57536 25832 57588
rect 26976 57536 27028 57588
rect 29368 57536 29420 57588
rect 34152 57536 34204 57588
rect 1860 57400 1912 57452
rect 3056 57400 3108 57452
rect 4252 57400 4304 57452
rect 4620 57400 4672 57452
rect 5540 57400 5592 57452
rect 7840 57400 7892 57452
rect 8484 57400 8536 57452
rect 9036 57400 9088 57452
rect 10232 57400 10284 57452
rect 11428 57400 11480 57452
rect 12624 57400 12676 57452
rect 13820 57400 13872 57452
rect 15016 57400 15068 57452
rect 16212 57400 16264 57452
rect 17408 57400 17460 57452
rect 18604 57400 18656 57452
rect 19984 57400 20036 57452
rect 20996 57400 21048 57452
rect 22192 57400 22244 57452
rect 23388 57400 23440 57452
rect 24584 57400 24636 57452
rect 3148 57375 3200 57384
rect 3148 57341 3157 57375
rect 3157 57341 3191 57375
rect 3191 57341 3200 57375
rect 3148 57332 3200 57341
rect 5724 57375 5776 57384
rect 5724 57341 5733 57375
rect 5733 57341 5767 57375
rect 5767 57341 5776 57375
rect 5724 57332 5776 57341
rect 8300 57375 8352 57384
rect 8300 57341 8309 57375
rect 8309 57341 8343 57375
rect 8343 57341 8352 57375
rect 8300 57332 8352 57341
rect 20536 57332 20588 57384
rect 24952 57332 25004 57384
rect 28172 57400 28224 57452
rect 30564 57400 30616 57452
rect 31760 57400 31812 57452
rect 32128 57400 32180 57452
rect 32956 57400 33008 57452
rect 38752 57536 38804 57588
rect 38844 57468 38896 57520
rect 42708 57536 42760 57588
rect 35348 57400 35400 57452
rect 36544 57400 36596 57452
rect 37740 57400 37792 57452
rect 38936 57400 38988 57452
rect 40132 57400 40184 57452
rect 41328 57400 41380 57452
rect 42800 57443 42852 57452
rect 42800 57409 42809 57443
rect 42809 57409 42843 57443
rect 42843 57409 42852 57443
rect 42800 57400 42852 57409
rect 43720 57400 43772 57452
rect 44916 57400 44968 57452
rect 46112 57400 46164 57452
rect 47308 57400 47360 57452
rect 48504 57400 48556 57452
rect 49700 57400 49752 57452
rect 50344 57400 50396 57452
rect 51080 57400 51132 57452
rect 52092 57400 52144 57452
rect 53288 57400 53340 57452
rect 54484 57400 54536 57452
rect 55680 57400 55732 57452
rect 56876 57400 56928 57452
rect 58072 57400 58124 57452
rect 30380 57332 30432 57384
rect 38384 57332 38436 57384
rect 25044 57264 25096 57316
rect 5448 57196 5500 57248
rect 9312 57239 9364 57248
rect 9312 57205 9321 57239
rect 9321 57205 9355 57239
rect 9355 57205 9364 57239
rect 9312 57196 9364 57205
rect 10508 57239 10560 57248
rect 10508 57205 10517 57239
rect 10517 57205 10551 57239
rect 10551 57205 10560 57239
rect 10508 57196 10560 57205
rect 11888 57239 11940 57248
rect 11888 57205 11897 57239
rect 11897 57205 11931 57239
rect 11931 57205 11940 57239
rect 11888 57196 11940 57205
rect 12900 57239 12952 57248
rect 12900 57205 12909 57239
rect 12909 57205 12943 57239
rect 12943 57205 12952 57239
rect 12900 57196 12952 57205
rect 14464 57239 14516 57248
rect 14464 57205 14473 57239
rect 14473 57205 14507 57239
rect 14507 57205 14516 57239
rect 14464 57196 14516 57205
rect 18880 57239 18932 57248
rect 18880 57205 18889 57239
rect 18889 57205 18923 57239
rect 18923 57205 18932 57239
rect 18880 57196 18932 57205
rect 20076 57239 20128 57248
rect 20076 57205 20085 57239
rect 20085 57205 20119 57239
rect 20119 57205 20128 57239
rect 20076 57196 20128 57205
rect 21272 57239 21324 57248
rect 21272 57205 21281 57239
rect 21281 57205 21315 57239
rect 21315 57205 21324 57239
rect 21272 57196 21324 57205
rect 24860 57239 24912 57248
rect 24860 57205 24869 57239
rect 24869 57205 24903 57239
rect 24903 57205 24912 57239
rect 24860 57196 24912 57205
rect 25872 57239 25924 57248
rect 25872 57205 25881 57239
rect 25881 57205 25915 57239
rect 25915 57205 25924 57239
rect 25872 57196 25924 57205
rect 26148 57196 26200 57248
rect 28356 57196 28408 57248
rect 29736 57239 29788 57248
rect 29736 57205 29745 57239
rect 29745 57205 29779 57239
rect 29779 57205 29788 57239
rect 29736 57196 29788 57205
rect 36452 57264 36504 57316
rect 32312 57196 32364 57248
rect 32956 57196 33008 57248
rect 33232 57239 33284 57248
rect 33232 57205 33241 57239
rect 33241 57205 33275 57239
rect 33275 57205 33284 57239
rect 33232 57196 33284 57205
rect 34704 57196 34756 57248
rect 35808 57196 35860 57248
rect 35900 57196 35952 57248
rect 37648 57196 37700 57248
rect 38660 57196 38712 57248
rect 44548 57332 44600 57384
rect 42800 57264 42852 57316
rect 44640 57264 44692 57316
rect 48596 57239 48648 57248
rect 48596 57205 48605 57239
rect 48605 57205 48639 57239
rect 48639 57205 48648 57239
rect 48596 57196 48648 57205
rect 48688 57196 48740 57248
rect 52184 57239 52236 57248
rect 52184 57205 52193 57239
rect 52193 57205 52227 57239
rect 52227 57205 52236 57239
rect 52184 57196 52236 57205
rect 53380 57239 53432 57248
rect 53380 57205 53389 57239
rect 53389 57205 53423 57239
rect 53423 57205 53432 57239
rect 53380 57196 53432 57205
rect 54576 57239 54628 57248
rect 54576 57205 54585 57239
rect 54585 57205 54619 57239
rect 54619 57205 54628 57239
rect 54576 57196 54628 57205
rect 55772 57239 55824 57248
rect 55772 57205 55781 57239
rect 55781 57205 55815 57239
rect 55815 57205 55824 57239
rect 55772 57196 55824 57205
rect 56968 57239 57020 57248
rect 56968 57205 56977 57239
rect 56977 57205 57011 57239
rect 57011 57205 57020 57239
rect 56968 57196 57020 57205
rect 58164 57239 58216 57248
rect 58164 57205 58173 57239
rect 58173 57205 58207 57239
rect 58207 57205 58216 57239
rect 58164 57196 58216 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 1860 57035 1912 57044
rect 1860 57001 1869 57035
rect 1869 57001 1903 57035
rect 1903 57001 1912 57035
rect 1860 56992 1912 57001
rect 3056 56992 3108 57044
rect 4620 56992 4672 57044
rect 8484 57035 8536 57044
rect 8484 57001 8493 57035
rect 8493 57001 8527 57035
rect 8527 57001 8536 57035
rect 8484 56992 8536 57001
rect 9036 56992 9088 57044
rect 12624 57035 12676 57044
rect 12624 57001 12633 57035
rect 12633 57001 12667 57035
rect 12667 57001 12676 57035
rect 12624 56992 12676 57001
rect 15016 57035 15068 57044
rect 15016 57001 15025 57035
rect 15025 57001 15059 57035
rect 15059 57001 15068 57035
rect 15016 56992 15068 57001
rect 17408 57035 17460 57044
rect 17408 57001 17417 57035
rect 17417 57001 17451 57035
rect 17451 57001 17460 57035
rect 17408 56992 17460 57001
rect 19984 56992 20036 57044
rect 22192 57035 22244 57044
rect 22192 57001 22201 57035
rect 22201 57001 22235 57035
rect 22235 57001 22244 57035
rect 22192 56992 22244 57001
rect 24584 57035 24636 57044
rect 24584 57001 24593 57035
rect 24593 57001 24627 57035
rect 24627 57001 24636 57035
rect 24584 56992 24636 57001
rect 28172 57035 28224 57044
rect 28172 57001 28181 57035
rect 28181 57001 28215 57035
rect 28215 57001 28224 57035
rect 28172 56992 28224 57001
rect 32128 57035 32180 57044
rect 32128 57001 32137 57035
rect 32137 57001 32171 57035
rect 32171 57001 32180 57035
rect 32128 56992 32180 57001
rect 35348 57035 35400 57044
rect 35348 57001 35357 57035
rect 35357 57001 35391 57035
rect 35391 57001 35400 57035
rect 35348 56992 35400 57001
rect 36544 57035 36596 57044
rect 36544 57001 36553 57035
rect 36553 57001 36587 57035
rect 36587 57001 36596 57035
rect 36544 56992 36596 57001
rect 38936 56992 38988 57044
rect 41328 57035 41380 57044
rect 41328 57001 41337 57035
rect 41337 57001 41371 57035
rect 41371 57001 41380 57035
rect 41328 56992 41380 57001
rect 44916 56992 44968 57044
rect 47308 56992 47360 57044
rect 50344 57035 50396 57044
rect 50344 57001 50353 57035
rect 50353 57001 50387 57035
rect 50387 57001 50396 57035
rect 50344 56992 50396 57001
rect 52092 57035 52144 57044
rect 52092 57001 52101 57035
rect 52101 57001 52135 57035
rect 52135 57001 52144 57035
rect 52092 56992 52144 57001
rect 54484 57035 54536 57044
rect 54484 57001 54493 57035
rect 54493 57001 54527 57035
rect 54527 57001 54536 57035
rect 54484 56992 54536 57001
rect 56876 56992 56928 57044
rect 9312 56924 9364 56976
rect 17224 56924 17276 56976
rect 29184 56924 29236 56976
rect 37832 56924 37884 56976
rect 44732 56924 44784 56976
rect 48596 56924 48648 56976
rect 6644 56856 6696 56908
rect 10508 56856 10560 56908
rect 17960 56856 18012 56908
rect 20076 56856 20128 56908
rect 26240 56856 26292 56908
rect 29736 56899 29788 56908
rect 29736 56865 29745 56899
rect 29745 56865 29779 56899
rect 29779 56865 29788 56899
rect 29736 56856 29788 56865
rect 7012 56831 7064 56840
rect 7012 56797 7021 56831
rect 7021 56797 7055 56831
rect 7055 56797 7064 56831
rect 7012 56788 7064 56797
rect 11888 56788 11940 56840
rect 19340 56788 19392 56840
rect 21272 56788 21324 56840
rect 29368 56788 29420 56840
rect 29828 56831 29880 56840
rect 29828 56797 29837 56831
rect 29837 56797 29871 56831
rect 29871 56797 29880 56831
rect 29828 56788 29880 56797
rect 38752 56831 38804 56840
rect 12900 56720 12952 56772
rect 20812 56720 20864 56772
rect 21180 56763 21232 56772
rect 21180 56729 21189 56763
rect 21189 56729 21223 56763
rect 21223 56729 21232 56763
rect 21180 56720 21232 56729
rect 14464 56652 14516 56704
rect 29460 56720 29512 56772
rect 38752 56797 38764 56831
rect 38764 56797 38798 56831
rect 38798 56797 38804 56831
rect 38752 56788 38804 56797
rect 39028 56797 39030 56818
rect 39030 56797 39080 56818
rect 39028 56766 39080 56797
rect 39120 56831 39172 56840
rect 39120 56797 39129 56831
rect 39129 56797 39163 56831
rect 39163 56797 39172 56831
rect 39120 56788 39172 56797
rect 43352 56788 43404 56840
rect 48688 56856 48740 56908
rect 43628 56763 43680 56772
rect 43628 56729 43637 56763
rect 43637 56729 43671 56763
rect 43671 56729 43680 56763
rect 43628 56720 43680 56729
rect 43904 56831 43956 56840
rect 43904 56797 43913 56831
rect 43913 56797 43947 56831
rect 43947 56797 43956 56831
rect 57060 56831 57112 56840
rect 43904 56788 43956 56797
rect 57060 56797 57069 56831
rect 57069 56797 57103 56831
rect 57103 56797 57112 56831
rect 57060 56788 57112 56797
rect 57520 56831 57572 56840
rect 57520 56797 57529 56831
rect 57529 56797 57563 56831
rect 57563 56797 57572 56831
rect 57520 56788 57572 56797
rect 58348 56831 58400 56840
rect 58348 56797 58357 56831
rect 58357 56797 58391 56831
rect 58391 56797 58400 56831
rect 58348 56788 58400 56797
rect 56968 56720 57020 56772
rect 30196 56695 30248 56704
rect 30196 56661 30205 56695
rect 30205 56661 30239 56695
rect 30239 56661 30248 56695
rect 30196 56652 30248 56661
rect 35992 56652 36044 56704
rect 38752 56652 38804 56704
rect 56876 56695 56928 56704
rect 56876 56661 56885 56695
rect 56885 56661 56919 56695
rect 56919 56661 56928 56695
rect 56876 56652 56928 56661
rect 57704 56695 57756 56704
rect 57704 56661 57713 56695
rect 57713 56661 57747 56695
rect 57747 56661 57756 56695
rect 57704 56652 57756 56661
rect 59176 56652 59228 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 17224 56448 17276 56500
rect 17960 56380 18012 56432
rect 24952 56448 25004 56500
rect 21180 56312 21232 56364
rect 21916 56312 21968 56364
rect 23756 56355 23808 56364
rect 23756 56321 23760 56355
rect 23760 56321 23794 56355
rect 23794 56321 23808 56355
rect 23756 56312 23808 56321
rect 25320 56380 25372 56432
rect 27436 56448 27488 56500
rect 20720 56244 20772 56296
rect 24216 56355 24268 56364
rect 24216 56321 24225 56355
rect 24225 56321 24259 56355
rect 24259 56321 24268 56355
rect 24216 56312 24268 56321
rect 24860 56312 24912 56364
rect 25228 56355 25280 56364
rect 25228 56321 25237 56355
rect 25237 56321 25271 56355
rect 25271 56321 25280 56355
rect 25228 56312 25280 56321
rect 25780 56312 25832 56364
rect 29368 56380 29420 56432
rect 24584 56244 24636 56296
rect 26424 56312 26476 56364
rect 26884 56244 26936 56296
rect 27344 56244 27396 56296
rect 27528 56355 27580 56364
rect 27528 56321 27542 56355
rect 27542 56321 27576 56355
rect 27576 56321 27580 56355
rect 27528 56312 27580 56321
rect 28540 56244 28592 56296
rect 28816 56355 28868 56364
rect 28816 56321 28826 56355
rect 28826 56321 28860 56355
rect 28860 56321 28868 56355
rect 28816 56312 28868 56321
rect 28954 56355 29006 56370
rect 28954 56321 28963 56355
rect 28963 56321 28997 56355
rect 28997 56321 29006 56355
rect 28954 56318 29006 56321
rect 30472 56448 30524 56500
rect 31024 56380 31076 56432
rect 31392 56448 31444 56500
rect 34980 56448 35032 56500
rect 35992 56448 36044 56500
rect 38016 56448 38068 56500
rect 32312 56380 32364 56432
rect 30196 56355 30248 56364
rect 30196 56321 30203 56355
rect 30203 56321 30248 56355
rect 30196 56312 30248 56321
rect 30380 56355 30432 56364
rect 30380 56321 30389 56355
rect 30389 56321 30423 56355
rect 30423 56321 30432 56355
rect 30380 56312 30432 56321
rect 30472 56355 30524 56364
rect 30472 56321 30486 56355
rect 30486 56321 30520 56355
rect 30520 56321 30524 56355
rect 30472 56312 30524 56321
rect 30656 56312 30708 56364
rect 31208 56312 31260 56364
rect 31668 56312 31720 56364
rect 32772 56355 32824 56364
rect 32772 56321 32776 56355
rect 32776 56321 32810 56355
rect 32810 56321 32824 56355
rect 32772 56312 32824 56321
rect 33048 56312 33100 56364
rect 34520 56380 34572 56432
rect 34704 56423 34756 56432
rect 34704 56389 34713 56423
rect 34713 56389 34747 56423
rect 34747 56389 34756 56423
rect 34704 56380 34756 56389
rect 35808 56423 35860 56432
rect 33324 56312 33376 56364
rect 34612 56355 34664 56364
rect 34612 56321 34616 56355
rect 34616 56321 34650 56355
rect 34650 56321 34664 56355
rect 34612 56312 34664 56321
rect 34980 56355 35032 56364
rect 34980 56321 34988 56355
rect 34988 56321 35022 56355
rect 35022 56321 35032 56355
rect 34980 56312 35032 56321
rect 35072 56355 35124 56364
rect 35072 56321 35081 56355
rect 35081 56321 35115 56355
rect 35115 56321 35124 56355
rect 35072 56312 35124 56321
rect 35532 56312 35584 56364
rect 30840 56244 30892 56296
rect 35808 56389 35817 56423
rect 35817 56389 35851 56423
rect 35851 56389 35860 56423
rect 35808 56380 35860 56389
rect 37832 56380 37884 56432
rect 35716 56355 35768 56364
rect 35716 56321 35720 56355
rect 35720 56321 35754 56355
rect 35754 56321 35768 56355
rect 36084 56355 36136 56364
rect 35716 56312 35768 56321
rect 36084 56321 36092 56355
rect 36092 56321 36126 56355
rect 36126 56321 36136 56355
rect 36084 56312 36136 56321
rect 36176 56355 36228 56364
rect 36176 56321 36185 56355
rect 36185 56321 36219 56355
rect 36219 56321 36228 56355
rect 37648 56355 37700 56364
rect 36176 56312 36228 56321
rect 37648 56321 37657 56355
rect 37657 56321 37691 56355
rect 37691 56321 37700 56355
rect 37648 56312 37700 56321
rect 37740 56355 37792 56364
rect 37740 56321 37749 56355
rect 37749 56321 37783 56355
rect 37783 56321 37792 56355
rect 37740 56312 37792 56321
rect 38016 56355 38068 56364
rect 38016 56321 38025 56355
rect 38025 56321 38059 56355
rect 38059 56321 38068 56355
rect 38660 56355 38712 56364
rect 38016 56312 38068 56321
rect 38660 56321 38669 56355
rect 38669 56321 38703 56355
rect 38703 56321 38712 56355
rect 38660 56312 38712 56321
rect 38752 56355 38804 56364
rect 38752 56321 38761 56355
rect 38761 56321 38795 56355
rect 38795 56321 38804 56355
rect 38936 56355 38988 56364
rect 38752 56312 38804 56321
rect 38936 56321 38945 56355
rect 38945 56321 38979 56355
rect 38979 56321 38988 56355
rect 38936 56312 38988 56321
rect 39028 56355 39080 56364
rect 39028 56321 39037 56355
rect 39037 56321 39071 56355
rect 39071 56321 39080 56355
rect 40776 56355 40828 56364
rect 39028 56312 39080 56321
rect 40776 56321 40780 56355
rect 40780 56321 40814 56355
rect 40814 56321 40828 56355
rect 40776 56312 40828 56321
rect 40500 56244 40552 56296
rect 23388 56108 23440 56160
rect 23572 56151 23624 56160
rect 23572 56117 23581 56151
rect 23581 56117 23615 56151
rect 23615 56117 23624 56151
rect 23572 56108 23624 56117
rect 25136 56108 25188 56160
rect 25320 56108 25372 56160
rect 28632 56176 28684 56228
rect 28724 56108 28776 56160
rect 33140 56176 33192 56228
rect 33324 56176 33376 56228
rect 35072 56176 35124 56228
rect 35164 56176 35216 56228
rect 35624 56176 35676 56228
rect 40960 56355 41012 56364
rect 40960 56321 40969 56355
rect 40969 56321 41003 56355
rect 41003 56321 41012 56355
rect 42708 56380 42760 56432
rect 42984 56380 43036 56432
rect 43628 56380 43680 56432
rect 40960 56312 41012 56321
rect 41236 56355 41288 56364
rect 41236 56321 41245 56355
rect 41245 56321 41279 56355
rect 41279 56321 41288 56355
rect 41236 56312 41288 56321
rect 42616 56312 42668 56364
rect 43352 56312 43404 56364
rect 44640 56448 44692 56500
rect 57060 56448 57112 56500
rect 57520 56380 57572 56432
rect 43904 56312 43956 56364
rect 58072 56312 58124 56364
rect 58440 56312 58492 56364
rect 58164 56244 58216 56296
rect 53380 56176 53432 56228
rect 29920 56108 29972 56160
rect 32588 56151 32640 56160
rect 32588 56117 32597 56151
rect 32597 56117 32631 56151
rect 32631 56117 32640 56151
rect 32588 56108 32640 56117
rect 33048 56108 33100 56160
rect 37556 56108 37608 56160
rect 38660 56108 38712 56160
rect 41144 56108 41196 56160
rect 43168 56151 43220 56160
rect 43168 56117 43177 56151
rect 43177 56117 43211 56151
rect 43211 56117 43220 56151
rect 43168 56108 43220 56117
rect 58164 56151 58216 56160
rect 58164 56117 58173 56151
rect 58173 56117 58207 56151
rect 58207 56117 58216 56151
rect 58164 56108 58216 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 20904 55904 20956 55956
rect 23664 55904 23716 55956
rect 24584 55947 24636 55956
rect 24584 55913 24593 55947
rect 24593 55913 24627 55947
rect 24627 55913 24636 55947
rect 24584 55904 24636 55913
rect 28816 55947 28868 55956
rect 23940 55879 23992 55888
rect 23940 55845 23949 55879
rect 23949 55845 23983 55879
rect 23983 55845 23992 55879
rect 23940 55836 23992 55845
rect 8300 55768 8352 55820
rect 20536 55700 20588 55752
rect 23388 55743 23440 55752
rect 23388 55709 23397 55743
rect 23397 55709 23431 55743
rect 23431 55709 23440 55743
rect 23388 55700 23440 55709
rect 23572 55743 23624 55752
rect 23572 55709 23581 55743
rect 23581 55709 23615 55743
rect 23615 55709 23624 55743
rect 23572 55700 23624 55709
rect 23664 55743 23716 55752
rect 23664 55709 23673 55743
rect 23673 55709 23707 55743
rect 23707 55709 23716 55743
rect 23664 55700 23716 55709
rect 24676 55700 24728 55752
rect 25228 55836 25280 55888
rect 25412 55836 25464 55888
rect 25780 55836 25832 55888
rect 26608 55836 26660 55888
rect 25044 55811 25096 55820
rect 25044 55777 25053 55811
rect 25053 55777 25087 55811
rect 25087 55777 25096 55811
rect 25044 55768 25096 55777
rect 28356 55811 28408 55820
rect 28356 55777 28365 55811
rect 28365 55777 28399 55811
rect 28399 55777 28408 55811
rect 28356 55768 28408 55777
rect 28816 55913 28825 55947
rect 28825 55913 28859 55947
rect 28859 55913 28868 55947
rect 28816 55904 28868 55913
rect 28908 55904 28960 55956
rect 36084 55904 36136 55956
rect 38614 55904 38666 55956
rect 40960 55904 41012 55956
rect 41512 55904 41564 55956
rect 58440 55904 58492 55956
rect 30288 55879 30340 55888
rect 30288 55845 30297 55879
rect 30297 55845 30331 55879
rect 30331 55845 30340 55879
rect 30288 55836 30340 55845
rect 31024 55836 31076 55888
rect 31208 55768 31260 55820
rect 37556 55836 37608 55888
rect 38292 55836 38344 55888
rect 41144 55879 41196 55888
rect 41144 55845 41153 55879
rect 41153 55845 41187 55879
rect 41187 55845 41196 55879
rect 41144 55836 41196 55845
rect 25136 55700 25188 55752
rect 25780 55700 25832 55752
rect 26976 55743 27028 55752
rect 26976 55709 26985 55743
rect 26985 55709 27019 55743
rect 27019 55709 27028 55743
rect 26976 55700 27028 55709
rect 27344 55700 27396 55752
rect 28448 55743 28500 55752
rect 28448 55709 28457 55743
rect 28457 55709 28491 55743
rect 28491 55709 28500 55743
rect 28448 55700 28500 55709
rect 1676 55607 1728 55616
rect 1676 55573 1685 55607
rect 1685 55573 1719 55607
rect 1719 55573 1728 55607
rect 1676 55564 1728 55573
rect 2320 55607 2372 55616
rect 2320 55573 2329 55607
rect 2329 55573 2363 55607
rect 2363 55573 2372 55607
rect 2320 55564 2372 55573
rect 28356 55632 28408 55684
rect 29184 55700 29236 55752
rect 29920 55743 29972 55752
rect 29920 55709 29929 55743
rect 29929 55709 29963 55743
rect 29963 55709 29972 55743
rect 29920 55700 29972 55709
rect 32864 55743 32916 55752
rect 21916 55564 21968 55616
rect 25228 55564 25280 55616
rect 25964 55564 26016 55616
rect 29460 55632 29512 55684
rect 30012 55675 30064 55684
rect 30012 55641 30021 55675
rect 30021 55641 30055 55675
rect 30055 55641 30064 55675
rect 30012 55632 30064 55641
rect 28816 55564 28868 55616
rect 32864 55709 32868 55743
rect 32868 55709 32902 55743
rect 32902 55709 32916 55743
rect 32864 55700 32916 55709
rect 32956 55743 33008 55752
rect 32956 55709 32965 55743
rect 32965 55709 32999 55743
rect 32999 55709 33008 55743
rect 32956 55700 33008 55709
rect 33324 55743 33376 55752
rect 33324 55709 33333 55743
rect 33333 55709 33367 55743
rect 33367 55709 33376 55743
rect 33324 55700 33376 55709
rect 34612 55700 34664 55752
rect 35716 55700 35768 55752
rect 35900 55743 35952 55752
rect 35900 55709 35909 55743
rect 35909 55709 35943 55743
rect 35943 55709 35952 55743
rect 35900 55700 35952 55709
rect 31760 55632 31812 55684
rect 35624 55632 35676 55684
rect 36268 55743 36320 55752
rect 36268 55709 36277 55743
rect 36277 55709 36311 55743
rect 36311 55709 36320 55743
rect 36268 55700 36320 55709
rect 37740 55700 37792 55752
rect 38476 55700 38528 55752
rect 38844 55768 38896 55820
rect 37464 55632 37516 55684
rect 38752 55709 38761 55730
rect 38761 55709 38795 55730
rect 38795 55709 38804 55730
rect 38752 55678 38804 55709
rect 38844 55632 38896 55684
rect 40500 55700 40552 55752
rect 41052 55700 41104 55752
rect 52184 55768 52236 55820
rect 39028 55632 39080 55684
rect 41512 55675 41564 55684
rect 41512 55641 41521 55675
rect 41521 55641 41555 55675
rect 41555 55641 41564 55675
rect 41512 55632 41564 55641
rect 41788 55743 41840 55752
rect 41788 55709 41797 55743
rect 41797 55709 41831 55743
rect 41831 55709 41840 55743
rect 41788 55700 41840 55709
rect 42616 55700 42668 55752
rect 43628 55743 43680 55752
rect 43628 55709 43637 55743
rect 43637 55709 43671 55743
rect 43671 55709 43680 55743
rect 43628 55700 43680 55709
rect 42800 55632 42852 55684
rect 43904 55743 43956 55752
rect 43904 55709 43913 55743
rect 43913 55709 43947 55743
rect 43947 55709 43956 55743
rect 43904 55700 43956 55709
rect 58348 55743 58400 55752
rect 58348 55709 58357 55743
rect 58357 55709 58391 55743
rect 58391 55709 58400 55743
rect 58348 55700 58400 55709
rect 43168 55564 43220 55616
rect 44732 55632 44784 55684
rect 55772 55632 55824 55684
rect 59544 55564 59596 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 25780 55360 25832 55412
rect 28448 55360 28500 55412
rect 29000 55360 29052 55412
rect 29828 55360 29880 55412
rect 34520 55360 34572 55412
rect 38292 55360 38344 55412
rect 7012 55292 7064 55344
rect 30012 55292 30064 55344
rect 2412 55267 2464 55276
rect 2412 55233 2421 55267
rect 2421 55233 2455 55267
rect 2455 55233 2464 55267
rect 2412 55224 2464 55233
rect 20812 55224 20864 55276
rect 21916 55224 21968 55276
rect 26056 55224 26108 55276
rect 26608 55224 26660 55276
rect 28540 55224 28592 55276
rect 38752 55224 38804 55276
rect 35624 55156 35676 55208
rect 40316 55292 40368 55344
rect 41236 55292 41288 55344
rect 41788 55292 41840 55344
rect 43352 55360 43404 55412
rect 43904 55360 43956 55412
rect 56692 55360 56744 55412
rect 54576 55292 54628 55344
rect 39580 55267 39632 55276
rect 39580 55233 39589 55267
rect 39589 55233 39623 55267
rect 39623 55233 39632 55267
rect 39580 55224 39632 55233
rect 40868 55224 40920 55276
rect 42616 55224 42668 55276
rect 42984 55267 43036 55276
rect 42984 55233 42993 55267
rect 42993 55233 43027 55267
rect 43027 55233 43036 55267
rect 42984 55224 43036 55233
rect 41512 55156 41564 55208
rect 43352 55224 43404 55276
rect 44548 55224 44600 55276
rect 57980 55224 58032 55276
rect 1676 55063 1728 55072
rect 1676 55029 1685 55063
rect 1685 55029 1719 55063
rect 1719 55029 1728 55063
rect 1676 55020 1728 55029
rect 32404 55063 32456 55072
rect 32404 55029 32413 55063
rect 32413 55029 32447 55063
rect 32447 55029 32456 55063
rect 32404 55020 32456 55029
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 25780 54816 25832 54868
rect 19340 54612 19392 54664
rect 21916 54544 21968 54596
rect 32496 54748 32548 54800
rect 25964 54612 26016 54664
rect 26148 54655 26200 54664
rect 26148 54621 26157 54655
rect 26157 54621 26191 54655
rect 26191 54621 26200 54655
rect 26608 54655 26660 54664
rect 26148 54612 26200 54621
rect 26608 54621 26617 54655
rect 26617 54621 26651 54655
rect 26651 54621 26660 54655
rect 26608 54612 26660 54621
rect 31392 54680 31444 54732
rect 32864 54816 32916 54868
rect 34612 54816 34664 54868
rect 37464 54859 37516 54868
rect 37464 54825 37473 54859
rect 37473 54825 37507 54859
rect 37507 54825 37516 54859
rect 37464 54816 37516 54825
rect 26240 54544 26292 54596
rect 22928 54476 22980 54528
rect 23756 54476 23808 54528
rect 24400 54476 24452 54528
rect 27436 54544 27488 54596
rect 34704 54680 34756 54732
rect 37556 54680 37608 54732
rect 32404 54655 32456 54664
rect 32404 54621 32413 54655
rect 32413 54621 32447 54655
rect 32447 54621 32456 54655
rect 32404 54612 32456 54621
rect 34612 54612 34664 54664
rect 35440 54655 35492 54664
rect 35440 54621 35448 54655
rect 35448 54621 35482 54655
rect 35482 54621 35492 54655
rect 35440 54612 35492 54621
rect 35532 54655 35584 54664
rect 35532 54621 35541 54655
rect 35541 54621 35575 54655
rect 35575 54621 35584 54655
rect 38384 54680 38436 54732
rect 35532 54612 35584 54621
rect 37924 54655 37976 54664
rect 33232 54544 33284 54596
rect 35624 54544 35676 54596
rect 37556 54544 37608 54596
rect 37924 54621 37933 54655
rect 37933 54621 37967 54655
rect 37967 54621 37976 54655
rect 37924 54612 37976 54621
rect 38016 54655 38068 54664
rect 38016 54621 38025 54655
rect 38025 54621 38059 54655
rect 38059 54621 38068 54655
rect 38660 54655 38712 54664
rect 38016 54612 38068 54621
rect 38660 54621 38669 54655
rect 38669 54621 38703 54655
rect 38703 54621 38712 54655
rect 38660 54612 38712 54621
rect 39580 54544 39632 54596
rect 27344 54476 27396 54528
rect 31852 54519 31904 54528
rect 31852 54485 31861 54519
rect 31861 54485 31895 54519
rect 31895 54485 31904 54519
rect 31852 54476 31904 54485
rect 32772 54519 32824 54528
rect 32772 54485 32781 54519
rect 32781 54485 32815 54519
rect 32815 54485 32824 54519
rect 32772 54476 32824 54485
rect 34888 54519 34940 54528
rect 34888 54485 34897 54519
rect 34897 54485 34931 54519
rect 34931 54485 34940 54519
rect 34888 54476 34940 54485
rect 37924 54476 37976 54528
rect 38936 54476 38988 54528
rect 39672 54476 39724 54528
rect 58348 54519 58400 54528
rect 58348 54485 58357 54519
rect 58357 54485 58391 54519
rect 58391 54485 58400 54519
rect 58348 54476 58400 54485
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 1676 54043 1728 54052
rect 1676 54009 1685 54043
rect 1685 54009 1719 54043
rect 1719 54009 1728 54043
rect 1676 54000 1728 54009
rect 2872 53932 2924 53984
rect 5724 53932 5776 53984
rect 18880 54204 18932 54256
rect 24400 54179 24452 54188
rect 24400 54145 24404 54179
rect 24404 54145 24438 54179
rect 24438 54145 24452 54179
rect 24400 54136 24452 54145
rect 25412 54136 25464 54188
rect 25964 54204 26016 54256
rect 27344 54247 27396 54256
rect 27344 54213 27353 54247
rect 27353 54213 27387 54247
rect 27387 54213 27396 54247
rect 27344 54204 27396 54213
rect 30932 54272 30984 54324
rect 31852 54272 31904 54324
rect 32496 54315 32548 54324
rect 32496 54281 32505 54315
rect 32505 54281 32539 54315
rect 32539 54281 32548 54315
rect 32496 54272 32548 54281
rect 35348 54272 35400 54324
rect 35440 54272 35492 54324
rect 38016 54272 38068 54324
rect 39028 54272 39080 54324
rect 40316 54315 40368 54324
rect 40316 54281 40325 54315
rect 40325 54281 40359 54315
rect 40359 54281 40368 54315
rect 40316 54272 40368 54281
rect 40868 54272 40920 54324
rect 32312 54204 32364 54256
rect 32588 54204 32640 54256
rect 25688 54179 25740 54188
rect 25688 54145 25697 54179
rect 25697 54145 25731 54179
rect 25731 54145 25740 54179
rect 25688 54136 25740 54145
rect 25872 54136 25924 54188
rect 26056 54136 26108 54188
rect 27528 54179 27580 54188
rect 27528 54145 27542 54179
rect 27542 54145 27576 54179
rect 27576 54145 27580 54179
rect 27528 54136 27580 54145
rect 30564 54136 30616 54188
rect 32680 54179 32732 54188
rect 24676 54068 24728 54120
rect 32680 54145 32689 54179
rect 32689 54145 32723 54179
rect 32723 54145 32732 54179
rect 32680 54136 32732 54145
rect 29736 54068 29788 54120
rect 31852 54068 31904 54120
rect 32312 54111 32364 54120
rect 32312 54077 32321 54111
rect 32321 54077 32355 54111
rect 32355 54077 32364 54111
rect 32312 54068 32364 54077
rect 32404 54068 32456 54120
rect 34704 54136 34756 54188
rect 35348 54136 35400 54188
rect 36544 54179 36596 54188
rect 36544 54145 36545 54179
rect 36545 54145 36579 54179
rect 36579 54145 36596 54179
rect 37924 54204 37976 54256
rect 36544 54136 36596 54145
rect 36820 54179 36872 54188
rect 36820 54145 36829 54179
rect 36829 54145 36863 54179
rect 36863 54145 36872 54179
rect 38660 54204 38712 54256
rect 36820 54136 36872 54145
rect 39672 54136 39724 54188
rect 39580 54068 39632 54120
rect 58348 54179 58400 54188
rect 58348 54145 58357 54179
rect 58357 54145 58391 54179
rect 58391 54145 58400 54179
rect 58348 54136 58400 54145
rect 34888 54000 34940 54052
rect 36452 54000 36504 54052
rect 39672 54000 39724 54052
rect 24768 53932 24820 53984
rect 29460 53932 29512 53984
rect 29920 53932 29972 53984
rect 32312 53932 32364 53984
rect 36820 53932 36872 53984
rect 39580 53932 39632 53984
rect 58900 53932 58952 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 30840 53728 30892 53780
rect 29828 53660 29880 53712
rect 30472 53703 30524 53712
rect 30472 53669 30481 53703
rect 30481 53669 30515 53703
rect 30515 53669 30524 53703
rect 30472 53660 30524 53669
rect 24676 53592 24728 53644
rect 31760 53728 31812 53780
rect 37556 53771 37608 53780
rect 37556 53737 37565 53771
rect 37565 53737 37599 53771
rect 37599 53737 37608 53771
rect 37556 53728 37608 53737
rect 38476 53771 38528 53780
rect 38476 53737 38485 53771
rect 38485 53737 38519 53771
rect 38519 53737 38528 53771
rect 38476 53728 38528 53737
rect 39672 53728 39724 53780
rect 32588 53660 32640 53712
rect 1676 53431 1728 53440
rect 1676 53397 1685 53431
rect 1685 53397 1719 53431
rect 1719 53397 1728 53431
rect 1676 53388 1728 53397
rect 22928 53524 22980 53576
rect 24768 53567 24820 53576
rect 24768 53533 24777 53567
rect 24777 53533 24811 53567
rect 24811 53533 24820 53567
rect 24768 53524 24820 53533
rect 29736 53567 29788 53576
rect 29736 53533 29745 53567
rect 29745 53533 29779 53567
rect 29779 53533 29788 53567
rect 29736 53524 29788 53533
rect 29920 53524 29972 53576
rect 32772 53592 32824 53644
rect 36544 53660 36596 53712
rect 39580 53660 39632 53712
rect 41512 53728 41564 53780
rect 30564 53567 30616 53576
rect 30564 53533 30573 53567
rect 30573 53533 30607 53567
rect 30607 53533 30616 53567
rect 30564 53524 30616 53533
rect 2504 53388 2556 53440
rect 5448 53388 5500 53440
rect 32312 53524 32364 53576
rect 32588 53567 32640 53576
rect 32588 53533 32597 53567
rect 32597 53533 32631 53567
rect 32631 53533 32640 53567
rect 32588 53524 32640 53533
rect 32680 53524 32732 53576
rect 38660 53524 38712 53576
rect 58348 53567 58400 53576
rect 35348 53456 35400 53508
rect 37556 53456 37608 53508
rect 58348 53533 58357 53567
rect 58357 53533 58391 53567
rect 58391 53533 58400 53567
rect 58348 53524 58400 53533
rect 32588 53388 32640 53440
rect 58532 53388 58584 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 29000 53184 29052 53236
rect 32772 53184 32824 53236
rect 39580 53184 39632 53236
rect 2412 53048 2464 53100
rect 10600 53048 10652 53100
rect 32404 53116 32456 53168
rect 29920 53091 29972 53100
rect 29920 53057 29929 53091
rect 29929 53057 29963 53091
rect 29963 53057 29972 53091
rect 29920 53048 29972 53057
rect 32312 53048 32364 53100
rect 29736 52980 29788 53032
rect 28816 52887 28868 52896
rect 28816 52853 28825 52887
rect 28825 52853 28859 52887
rect 28859 52853 28868 52887
rect 28816 52844 28868 52853
rect 39672 52887 39724 52896
rect 39672 52853 39681 52887
rect 39681 52853 39715 52887
rect 39715 52853 39724 52887
rect 39672 52844 39724 52853
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 29736 52640 29788 52692
rect 1676 52615 1728 52624
rect 1676 52581 1685 52615
rect 1685 52581 1719 52615
rect 1719 52581 1728 52615
rect 1676 52572 1728 52581
rect 58716 52572 58768 52624
rect 2780 52436 2832 52488
rect 55496 52436 55548 52488
rect 56876 52436 56928 52488
rect 58348 52479 58400 52488
rect 58348 52445 58357 52479
rect 58357 52445 58391 52479
rect 58391 52445 58400 52479
rect 58348 52436 58400 52445
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 1676 51799 1728 51808
rect 1676 51765 1685 51799
rect 1685 51765 1719 51799
rect 1719 51765 1728 51799
rect 1676 51756 1728 51765
rect 58348 52003 58400 52012
rect 58348 51969 58357 52003
rect 58357 51969 58391 52003
rect 58391 51969 58400 52003
rect 58348 51960 58400 51969
rect 4804 51756 4856 51808
rect 59084 51756 59136 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 58348 51255 58400 51264
rect 58348 51221 58357 51255
rect 58357 51221 58391 51255
rect 58391 51221 58400 51255
rect 58348 51212 58400 51221
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 2504 51008 2556 51060
rect 3608 51008 3660 51060
rect 58348 50915 58400 50924
rect 1676 50779 1728 50788
rect 1676 50745 1685 50779
rect 1685 50745 1719 50779
rect 1719 50745 1728 50779
rect 1676 50736 1728 50745
rect 58348 50881 58357 50915
rect 58357 50881 58391 50915
rect 58391 50881 58400 50915
rect 58348 50872 58400 50881
rect 2596 50668 2648 50720
rect 58808 50668 58860 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 2780 50328 2832 50380
rect 19064 50328 19116 50380
rect 1952 50260 2004 50312
rect 58348 50303 58400 50312
rect 58348 50269 58357 50303
rect 58357 50269 58391 50303
rect 58391 50269 58400 50303
rect 58348 50260 58400 50269
rect 1676 50167 1728 50176
rect 1676 50133 1685 50167
rect 1685 50133 1719 50167
rect 1719 50133 1728 50167
rect 1676 50124 1728 50133
rect 58440 50124 58492 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 10784 49172 10836 49224
rect 58348 49215 58400 49224
rect 58348 49181 58357 49215
rect 58357 49181 58391 49215
rect 58391 49181 58400 49215
rect 58348 49172 58400 49181
rect 1676 49079 1728 49088
rect 1676 49045 1685 49079
rect 1685 49045 1719 49079
rect 1719 49045 1728 49079
rect 1676 49036 1728 49045
rect 57980 49036 58032 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 2044 48696 2096 48748
rect 58348 48739 58400 48748
rect 58348 48705 58357 48739
rect 58357 48705 58391 48739
rect 58391 48705 58400 48739
rect 58348 48696 58400 48705
rect 1676 48535 1728 48544
rect 1676 48501 1685 48535
rect 1685 48501 1719 48535
rect 1719 48501 1728 48535
rect 1676 48492 1728 48501
rect 2044 48492 2096 48544
rect 57336 48492 57388 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 58348 47991 58400 48000
rect 58348 47957 58357 47991
rect 58357 47957 58391 47991
rect 58391 47957 58400 47991
rect 58348 47948 58400 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 58348 47651 58400 47660
rect 1676 47515 1728 47524
rect 1676 47481 1685 47515
rect 1685 47481 1719 47515
rect 1719 47481 1728 47515
rect 1676 47472 1728 47481
rect 58348 47617 58357 47651
rect 58357 47617 58391 47651
rect 58391 47617 58400 47651
rect 58348 47608 58400 47617
rect 2872 47540 2924 47592
rect 15200 47540 15252 47592
rect 4712 47404 4764 47456
rect 58256 47404 58308 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 58624 47132 58676 47184
rect 58348 47039 58400 47048
rect 58348 47005 58357 47039
rect 58357 47005 58391 47039
rect 58391 47005 58400 47039
rect 58348 46996 58400 47005
rect 2136 46928 2188 46980
rect 1676 46903 1728 46912
rect 1676 46869 1685 46903
rect 1685 46869 1719 46903
rect 1719 46869 1728 46903
rect 1676 46860 1728 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 1676 45815 1728 45824
rect 1676 45781 1685 45815
rect 1685 45781 1719 45815
rect 1719 45781 1728 45815
rect 1676 45772 1728 45781
rect 58348 45951 58400 45960
rect 58348 45917 58357 45951
rect 58357 45917 58391 45951
rect 58391 45917 58400 45951
rect 58348 45908 58400 45917
rect 3056 45772 3108 45824
rect 59636 45772 59688 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 1676 45271 1728 45280
rect 1676 45237 1685 45271
rect 1685 45237 1719 45271
rect 1719 45237 1728 45271
rect 1676 45228 1728 45237
rect 58348 45475 58400 45484
rect 58348 45441 58357 45475
rect 58357 45441 58391 45475
rect 58391 45441 58400 45475
rect 58348 45432 58400 45441
rect 9588 45228 9640 45280
rect 59268 45228 59320 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 2412 44820 2464 44872
rect 17408 44820 17460 44872
rect 58348 44727 58400 44736
rect 58348 44693 58357 44727
rect 58357 44693 58391 44727
rect 58391 44693 58400 44727
rect 58348 44684 58400 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 58348 44387 58400 44396
rect 1676 44251 1728 44260
rect 1676 44217 1685 44251
rect 1685 44217 1719 44251
rect 1719 44217 1728 44251
rect 1676 44208 1728 44217
rect 58348 44353 58357 44387
rect 58357 44353 58391 44387
rect 58391 44353 58400 44387
rect 58348 44344 58400 44353
rect 6184 44140 6236 44192
rect 59360 44140 59412 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 1676 43639 1728 43648
rect 1676 43605 1685 43639
rect 1685 43605 1719 43639
rect 1719 43605 1728 43639
rect 1676 43596 1728 43605
rect 58348 43775 58400 43784
rect 58348 43741 58357 43775
rect 58357 43741 58391 43775
rect 58391 43741 58400 43775
rect 58348 43732 58400 43741
rect 3976 43596 4028 43648
rect 56784 43596 56836 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 15936 42644 15988 42696
rect 58348 42687 58400 42696
rect 58348 42653 58357 42687
rect 58357 42653 58391 42687
rect 58391 42653 58400 42687
rect 58348 42644 58400 42653
rect 1676 42551 1728 42560
rect 1676 42517 1685 42551
rect 1685 42517 1719 42551
rect 1719 42517 1728 42551
rect 1676 42508 1728 42517
rect 57796 42508 57848 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 14464 42168 14516 42220
rect 58348 42211 58400 42220
rect 58348 42177 58357 42211
rect 58357 42177 58391 42211
rect 58391 42177 58400 42211
rect 58348 42168 58400 42177
rect 1676 42007 1728 42016
rect 1676 41973 1685 42007
rect 1685 41973 1719 42007
rect 1719 41973 1728 42007
rect 1676 41964 1728 41973
rect 58992 41964 59044 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 58348 41463 58400 41472
rect 58348 41429 58357 41463
rect 58357 41429 58391 41463
rect 58391 41429 58400 41463
rect 58348 41420 58400 41429
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 58348 41123 58400 41132
rect 1676 40987 1728 40996
rect 1676 40953 1685 40987
rect 1685 40953 1719 40987
rect 1719 40953 1728 40987
rect 1676 40944 1728 40953
rect 58348 41089 58357 41123
rect 58357 41089 58391 41123
rect 58391 41089 58400 41123
rect 58348 41080 58400 41089
rect 7564 40876 7616 40928
rect 57612 40876 57664 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 1676 40375 1728 40384
rect 1676 40341 1685 40375
rect 1685 40341 1719 40375
rect 1719 40341 1728 40375
rect 1676 40332 1728 40341
rect 58348 40511 58400 40520
rect 58348 40477 58357 40511
rect 58357 40477 58391 40511
rect 58391 40477 58400 40511
rect 58348 40468 58400 40477
rect 6276 40332 6328 40384
rect 57060 40332 57112 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 57244 40128 57296 40180
rect 57888 40060 57940 40112
rect 56416 39831 56468 39840
rect 56416 39797 56425 39831
rect 56425 39797 56459 39831
rect 56459 39797 56468 39831
rect 56416 39788 56468 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 56048 39448 56100 39500
rect 56416 39448 56468 39500
rect 57244 39423 57296 39432
rect 1676 39287 1728 39296
rect 1676 39253 1685 39287
rect 1685 39253 1719 39287
rect 1719 39253 1728 39287
rect 1676 39244 1728 39253
rect 57244 39389 57253 39423
rect 57253 39389 57287 39423
rect 57287 39389 57296 39423
rect 57244 39380 57296 39389
rect 57704 39423 57756 39432
rect 57704 39389 57713 39423
rect 57713 39389 57747 39423
rect 57747 39389 57756 39423
rect 57704 39380 57756 39389
rect 57980 39355 58032 39364
rect 57980 39321 57989 39355
rect 57989 39321 58023 39355
rect 58023 39321 58032 39355
rect 57980 39312 58032 39321
rect 7656 39244 7708 39296
rect 56140 39287 56192 39296
rect 56140 39253 56149 39287
rect 56149 39253 56183 39287
rect 56183 39253 56192 39287
rect 56140 39244 56192 39253
rect 56600 39244 56652 39296
rect 56876 39287 56928 39296
rect 56876 39253 56885 39287
rect 56885 39253 56919 39287
rect 56919 39253 56928 39287
rect 56876 39244 56928 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 57152 39040 57204 39092
rect 57336 39040 57388 39092
rect 1676 38743 1728 38752
rect 1676 38709 1685 38743
rect 1685 38709 1719 38743
rect 1719 38709 1728 38743
rect 1676 38700 1728 38709
rect 55404 38904 55456 38956
rect 56140 38904 56192 38956
rect 58164 38904 58216 38956
rect 58348 38947 58400 38956
rect 58348 38913 58357 38947
rect 58357 38913 58391 38947
rect 58391 38913 58400 38947
rect 58348 38904 58400 38913
rect 56048 38836 56100 38888
rect 2780 38700 2832 38752
rect 55404 38743 55456 38752
rect 55404 38709 55413 38743
rect 55413 38709 55447 38743
rect 55447 38709 55456 38743
rect 55404 38700 55456 38709
rect 55956 38743 56008 38752
rect 55956 38709 55965 38743
rect 55965 38709 55999 38743
rect 55999 38709 56008 38743
rect 55956 38700 56008 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 57060 38539 57112 38548
rect 57060 38505 57069 38539
rect 57069 38505 57103 38539
rect 57103 38505 57112 38539
rect 57060 38496 57112 38505
rect 58164 38496 58216 38548
rect 56048 38156 56100 38208
rect 58348 38199 58400 38208
rect 58348 38165 58357 38199
rect 58357 38165 58391 38199
rect 58391 38165 58400 38199
rect 58348 38156 58400 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 54852 37884 54904 37936
rect 55496 37927 55548 37936
rect 55496 37893 55505 37927
rect 55505 37893 55539 37927
rect 55539 37893 55548 37927
rect 55496 37884 55548 37893
rect 1676 37723 1728 37732
rect 1676 37689 1685 37723
rect 1685 37689 1719 37723
rect 1719 37689 1728 37723
rect 1676 37680 1728 37689
rect 55404 37859 55456 37868
rect 55404 37825 55413 37859
rect 55413 37825 55447 37859
rect 55447 37825 55456 37859
rect 55404 37816 55456 37825
rect 55864 37884 55916 37936
rect 58256 37884 58308 37936
rect 58348 37859 58400 37868
rect 58348 37825 58357 37859
rect 58357 37825 58391 37859
rect 58391 37825 58400 37859
rect 58348 37816 58400 37825
rect 2780 37748 2832 37800
rect 4620 37748 4672 37800
rect 56048 37748 56100 37800
rect 56508 37748 56560 37800
rect 2412 37655 2464 37664
rect 2412 37621 2421 37655
rect 2421 37621 2455 37655
rect 2455 37621 2464 37655
rect 2412 37612 2464 37621
rect 54576 37612 54628 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2412 37408 2464 37460
rect 13636 37408 13688 37460
rect 56048 37408 56100 37460
rect 57888 37272 57940 37324
rect 58348 37247 58400 37256
rect 58348 37213 58357 37247
rect 58357 37213 58391 37247
rect 58391 37213 58400 37247
rect 58348 37204 58400 37213
rect 1676 37111 1728 37120
rect 1676 37077 1685 37111
rect 1685 37077 1719 37111
rect 1719 37077 1728 37111
rect 1676 37068 1728 37077
rect 2412 37111 2464 37120
rect 2412 37077 2421 37111
rect 2421 37077 2455 37111
rect 2455 37077 2464 37111
rect 2412 37068 2464 37077
rect 57428 37068 57480 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 2412 36864 2464 36916
rect 16580 36864 16632 36916
rect 57980 36864 58032 36916
rect 59176 36864 59228 36916
rect 57888 36728 57940 36780
rect 56508 36524 56560 36576
rect 58072 36524 58124 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 53104 36252 53156 36304
rect 56508 36184 56560 36236
rect 8484 36116 8536 36168
rect 57428 36159 57480 36168
rect 57428 36125 57437 36159
rect 57437 36125 57471 36159
rect 57471 36125 57480 36159
rect 57428 36116 57480 36125
rect 57980 36116 58032 36168
rect 55404 36048 55456 36100
rect 56324 36091 56376 36100
rect 56324 36057 56333 36091
rect 56333 36057 56367 36091
rect 56367 36057 56376 36091
rect 56324 36048 56376 36057
rect 1676 36023 1728 36032
rect 1676 35989 1685 36023
rect 1685 35989 1719 36023
rect 1719 35989 1728 36023
rect 1676 35980 1728 35989
rect 59452 36048 59504 36100
rect 58624 35980 58676 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 57980 35776 58032 35828
rect 59544 35776 59596 35828
rect 11704 35640 11756 35692
rect 58348 35683 58400 35692
rect 58348 35649 58357 35683
rect 58357 35649 58391 35683
rect 58391 35649 58400 35683
rect 58348 35640 58400 35649
rect 1676 35479 1728 35488
rect 1676 35445 1685 35479
rect 1685 35445 1719 35479
rect 1719 35445 1728 35479
rect 1676 35436 1728 35445
rect 56416 35436 56468 35488
rect 57520 35436 57572 35488
rect 58164 35479 58216 35488
rect 58164 35445 58173 35479
rect 58173 35445 58207 35479
rect 58207 35445 58216 35479
rect 58164 35436 58216 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 57152 35232 57204 35284
rect 59636 35232 59688 35284
rect 6276 35164 6328 35216
rect 16028 35164 16080 35216
rect 55772 35096 55824 35148
rect 56324 35096 56376 35148
rect 57152 35139 57204 35148
rect 57152 35105 57170 35139
rect 57170 35105 57204 35139
rect 57152 35096 57204 35105
rect 57980 35164 58032 35216
rect 57520 35139 57572 35148
rect 57520 35105 57529 35139
rect 57529 35105 57563 35139
rect 57563 35105 57572 35139
rect 57520 35096 57572 35105
rect 58072 35096 58124 35148
rect 52368 34960 52420 35012
rect 58072 34960 58124 35012
rect 55036 34892 55088 34944
rect 55772 34935 55824 34944
rect 55772 34901 55781 34935
rect 55781 34901 55815 34935
rect 55815 34901 55824 34935
rect 55772 34892 55824 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 55312 34688 55364 34740
rect 56692 34731 56744 34740
rect 56692 34697 56701 34731
rect 56701 34697 56735 34731
rect 56735 34697 56744 34731
rect 56692 34688 56744 34697
rect 52368 34595 52420 34604
rect 52368 34561 52377 34595
rect 52377 34561 52411 34595
rect 52411 34561 52420 34595
rect 52368 34552 52420 34561
rect 55312 34595 55364 34604
rect 55312 34561 55321 34595
rect 55321 34561 55355 34595
rect 55355 34561 55364 34595
rect 55312 34552 55364 34561
rect 58164 34620 58216 34672
rect 58348 34595 58400 34604
rect 58348 34561 58357 34595
rect 58357 34561 58391 34595
rect 58391 34561 58400 34595
rect 58348 34552 58400 34561
rect 6920 34484 6972 34536
rect 51448 34484 51500 34536
rect 55036 34527 55088 34536
rect 55036 34493 55045 34527
rect 55045 34493 55079 34527
rect 55079 34493 55088 34527
rect 55036 34484 55088 34493
rect 1676 34459 1728 34468
rect 1676 34425 1685 34459
rect 1685 34425 1719 34459
rect 1719 34425 1728 34459
rect 1676 34416 1728 34425
rect 55588 34459 55640 34468
rect 55588 34425 55597 34459
rect 55597 34425 55631 34459
rect 55631 34425 55640 34459
rect 55864 34484 55916 34536
rect 59268 34484 59320 34536
rect 55588 34416 55640 34425
rect 54392 34391 54444 34400
rect 54392 34357 54401 34391
rect 54401 34357 54435 34391
rect 54435 34357 54444 34391
rect 54392 34348 54444 34357
rect 56416 34348 56468 34400
rect 58164 34391 58216 34400
rect 58164 34357 58173 34391
rect 58173 34357 58207 34391
rect 58207 34357 58216 34391
rect 58164 34348 58216 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 55588 34144 55640 34196
rect 56968 34076 57020 34128
rect 2504 33940 2556 33992
rect 58348 33983 58400 33992
rect 58348 33949 58357 33983
rect 58357 33949 58391 33983
rect 58391 33949 58400 33983
rect 58348 33940 58400 33949
rect 1676 33847 1728 33856
rect 1676 33813 1685 33847
rect 1685 33813 1719 33847
rect 1719 33813 1728 33847
rect 1676 33804 1728 33813
rect 57796 33804 57848 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 57980 33600 58032 33652
rect 58532 33600 58584 33652
rect 54392 33464 54444 33516
rect 57796 33464 57848 33516
rect 54760 33439 54812 33448
rect 54760 33405 54769 33439
rect 54769 33405 54803 33439
rect 54803 33405 54812 33439
rect 54760 33396 54812 33405
rect 56876 33260 56928 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 48504 32988 48556 33040
rect 1676 32759 1728 32768
rect 1676 32725 1685 32759
rect 1685 32725 1719 32759
rect 1719 32725 1728 32759
rect 1676 32716 1728 32725
rect 56416 32852 56468 32904
rect 56968 32895 57020 32904
rect 56968 32861 56977 32895
rect 56977 32861 57011 32895
rect 57011 32861 57020 32895
rect 56968 32852 57020 32861
rect 57980 32852 58032 32904
rect 56784 32784 56836 32836
rect 2688 32716 2740 32768
rect 55772 32759 55824 32768
rect 55772 32725 55781 32759
rect 55781 32725 55815 32759
rect 55815 32725 55824 32759
rect 55772 32716 55824 32725
rect 57060 32716 57112 32768
rect 57520 32784 57572 32836
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 55772 32512 55824 32564
rect 57520 32512 57572 32564
rect 12440 32376 12492 32428
rect 58348 32419 58400 32428
rect 58348 32385 58357 32419
rect 58357 32385 58391 32419
rect 58391 32385 58400 32419
rect 58348 32376 58400 32385
rect 1676 32215 1728 32224
rect 1676 32181 1685 32215
rect 1685 32181 1719 32215
rect 1719 32181 1728 32215
rect 1676 32172 1728 32181
rect 56416 32172 56468 32224
rect 57428 32172 57480 32224
rect 58256 32172 58308 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 56968 31968 57020 32020
rect 59360 31968 59412 32020
rect 55772 31943 55824 31952
rect 55772 31909 55781 31943
rect 55781 31909 55815 31943
rect 55815 31909 55824 31943
rect 55772 31900 55824 31909
rect 56232 31900 56284 31952
rect 56968 31832 57020 31884
rect 57520 31900 57572 31952
rect 58900 31900 58952 31952
rect 57428 31875 57480 31884
rect 57428 31841 57437 31875
rect 57437 31841 57471 31875
rect 57471 31841 57480 31875
rect 57428 31832 57480 31841
rect 58164 31832 58216 31884
rect 54484 31764 54536 31816
rect 57980 31764 58032 31816
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 57520 31467 57572 31476
rect 57520 31433 57529 31467
rect 57529 31433 57563 31467
rect 57563 31433 57572 31467
rect 57520 31424 57572 31433
rect 56968 31356 57020 31408
rect 59084 31356 59136 31408
rect 2228 31288 2280 31340
rect 54484 31288 54536 31340
rect 58164 31331 58216 31340
rect 58164 31297 58173 31331
rect 58173 31297 58207 31331
rect 58207 31297 58216 31331
rect 58164 31288 58216 31297
rect 49056 31220 49108 31272
rect 1676 31195 1728 31204
rect 1676 31161 1685 31195
rect 1685 31161 1719 31195
rect 1719 31161 1728 31195
rect 1676 31152 1728 31161
rect 2228 31084 2280 31136
rect 56416 31084 56468 31136
rect 58532 31084 58584 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 58164 30880 58216 30932
rect 57520 30812 57572 30864
rect 58440 30812 58492 30864
rect 58440 30676 58492 30728
rect 1676 30583 1728 30592
rect 1676 30549 1685 30583
rect 1685 30549 1719 30583
rect 1719 30549 1728 30583
rect 1676 30540 1728 30549
rect 2412 30583 2464 30592
rect 2412 30549 2421 30583
rect 2421 30549 2455 30583
rect 2455 30549 2464 30583
rect 2412 30540 2464 30549
rect 58348 30583 58400 30592
rect 58348 30549 58357 30583
rect 58357 30549 58391 30583
rect 58391 30549 58400 30583
rect 58348 30540 58400 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 58440 30336 58492 30388
rect 12440 30268 12492 30320
rect 12624 30268 12676 30320
rect 14464 30268 14516 30320
rect 15660 30268 15712 30320
rect 56968 30311 57020 30320
rect 56968 30277 56977 30311
rect 56977 30277 57011 30311
rect 57011 30277 57020 30311
rect 56968 30268 57020 30277
rect 11060 30200 11112 30252
rect 12348 30175 12400 30184
rect 12348 30141 12357 30175
rect 12357 30141 12391 30175
rect 12391 30141 12400 30175
rect 12348 30132 12400 30141
rect 57152 30132 57204 30184
rect 57612 30132 57664 30184
rect 11060 30039 11112 30048
rect 11060 30005 11069 30039
rect 11069 30005 11103 30039
rect 11103 30005 11112 30039
rect 11060 29996 11112 30005
rect 11428 29996 11480 30048
rect 57152 29996 57204 30048
rect 57428 30039 57480 30048
rect 57428 30005 57437 30039
rect 57437 30005 57471 30039
rect 57471 30005 57480 30039
rect 57428 29996 57480 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 57704 29724 57756 29776
rect 11152 29656 11204 29708
rect 11428 29631 11480 29640
rect 11428 29597 11437 29631
rect 11437 29597 11471 29631
rect 11471 29597 11480 29631
rect 11428 29588 11480 29597
rect 58256 29588 58308 29640
rect 9220 29520 9272 29572
rect 9772 29563 9824 29572
rect 9772 29529 9781 29563
rect 9781 29529 9815 29563
rect 9815 29529 9824 29563
rect 9772 29520 9824 29529
rect 56140 29520 56192 29572
rect 57152 29520 57204 29572
rect 1676 29495 1728 29504
rect 1676 29461 1685 29495
rect 1685 29461 1719 29495
rect 1719 29461 1728 29495
rect 1676 29452 1728 29461
rect 11244 29495 11296 29504
rect 11244 29461 11253 29495
rect 11253 29461 11287 29495
rect 11287 29461 11296 29495
rect 11244 29452 11296 29461
rect 12348 29452 12400 29504
rect 55588 29452 55640 29504
rect 56968 29452 57020 29504
rect 58992 29520 59044 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 8484 29291 8536 29300
rect 8484 29257 8493 29291
rect 8493 29257 8527 29291
rect 8527 29257 8536 29291
rect 8484 29248 8536 29257
rect 10784 29248 10836 29300
rect 11980 29248 12032 29300
rect 57336 29291 57388 29300
rect 57336 29257 57345 29291
rect 57345 29257 57379 29291
rect 57379 29257 57388 29291
rect 57336 29248 57388 29257
rect 57612 29248 57664 29300
rect 15016 29180 15068 29232
rect 11152 29112 11204 29164
rect 1676 29019 1728 29028
rect 1676 28985 1685 29019
rect 1685 28985 1719 29019
rect 1719 28985 1728 29019
rect 1676 28976 1728 28985
rect 5908 28976 5960 29028
rect 9772 29044 9824 29096
rect 9956 28976 10008 29028
rect 58440 29112 58492 29164
rect 10968 28976 11020 29028
rect 57152 28976 57204 29028
rect 6828 28951 6880 28960
rect 6828 28917 6837 28951
rect 6837 28917 6871 28951
rect 6871 28917 6880 28951
rect 6828 28908 6880 28917
rect 7656 28908 7708 28960
rect 56968 28908 57020 28960
rect 57336 28908 57388 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 3792 28704 3844 28756
rect 5908 28611 5960 28620
rect 5908 28577 5917 28611
rect 5917 28577 5951 28611
rect 5951 28577 5960 28611
rect 5908 28568 5960 28577
rect 7932 28704 7984 28756
rect 8760 28636 8812 28688
rect 9588 28611 9640 28620
rect 6000 28500 6052 28552
rect 6828 28500 6880 28552
rect 7656 28543 7708 28552
rect 7656 28509 7665 28543
rect 7665 28509 7699 28543
rect 7699 28509 7708 28543
rect 7656 28500 7708 28509
rect 9588 28577 9597 28611
rect 9597 28577 9631 28611
rect 9631 28577 9640 28611
rect 9588 28568 9640 28577
rect 16580 28747 16632 28756
rect 16580 28713 16589 28747
rect 16589 28713 16623 28747
rect 16623 28713 16632 28747
rect 16580 28704 16632 28713
rect 9772 28636 9824 28688
rect 10968 28568 11020 28620
rect 12348 28611 12400 28620
rect 12348 28577 12357 28611
rect 12357 28577 12391 28611
rect 12391 28577 12400 28611
rect 12348 28568 12400 28577
rect 57704 28568 57756 28620
rect 9496 28543 9548 28552
rect 9496 28509 9505 28543
rect 9505 28509 9539 28543
rect 9539 28509 9548 28543
rect 9496 28500 9548 28509
rect 10508 28500 10560 28552
rect 11704 28500 11756 28552
rect 6920 28432 6972 28484
rect 7104 28432 7156 28484
rect 57336 28500 57388 28552
rect 57428 28500 57480 28552
rect 58716 28500 58768 28552
rect 57888 28475 57940 28484
rect 1952 28407 2004 28416
rect 1952 28373 1961 28407
rect 1961 28373 1995 28407
rect 1995 28373 2004 28407
rect 1952 28364 2004 28373
rect 4068 28364 4120 28416
rect 6828 28364 6880 28416
rect 9128 28407 9180 28416
rect 9128 28373 9137 28407
rect 9137 28373 9171 28407
rect 9171 28373 9180 28407
rect 9128 28364 9180 28373
rect 11152 28364 11204 28416
rect 12164 28407 12216 28416
rect 12164 28373 12173 28407
rect 12173 28373 12207 28407
rect 12207 28373 12216 28407
rect 12164 28364 12216 28373
rect 56784 28407 56836 28416
rect 56784 28373 56793 28407
rect 56793 28373 56827 28407
rect 56827 28373 56836 28407
rect 56784 28364 56836 28373
rect 57888 28441 57897 28475
rect 57897 28441 57931 28475
rect 57931 28441 57940 28475
rect 57888 28432 57940 28441
rect 57336 28364 57388 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 4712 28203 4764 28212
rect 4712 28169 4721 28203
rect 4721 28169 4755 28203
rect 4755 28169 4764 28203
rect 4712 28160 4764 28169
rect 6184 28160 6236 28212
rect 6460 28092 6512 28144
rect 1676 27931 1728 27940
rect 1676 27897 1685 27931
rect 1685 27897 1719 27931
rect 1719 27897 1728 27931
rect 1676 27888 1728 27897
rect 6000 28024 6052 28076
rect 6828 28067 6880 28076
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 3424 27956 3476 28008
rect 4068 27956 4120 28008
rect 7840 27999 7892 28008
rect 7840 27965 7849 27999
rect 7849 27965 7883 27999
rect 7883 27965 7892 27999
rect 7840 27956 7892 27965
rect 8116 28067 8168 28076
rect 8116 28033 8125 28067
rect 8125 28033 8159 28067
rect 8159 28033 8168 28067
rect 8116 28024 8168 28033
rect 12072 28160 12124 28212
rect 12348 28160 12400 28212
rect 9496 28092 9548 28144
rect 11060 28092 11112 28144
rect 11428 28092 11480 28144
rect 11704 28135 11756 28144
rect 11704 28101 11713 28135
rect 11713 28101 11747 28135
rect 11747 28101 11756 28135
rect 11704 28092 11756 28101
rect 16580 28092 16632 28144
rect 17224 28067 17276 28076
rect 5264 27888 5316 27940
rect 17224 28033 17233 28067
rect 17233 28033 17267 28067
rect 17267 28033 17276 28067
rect 17224 28024 17276 28033
rect 57152 28160 57204 28212
rect 57428 28160 57480 28212
rect 57704 28160 57756 28212
rect 56784 28092 56836 28144
rect 58716 28092 58768 28144
rect 58440 28024 58492 28076
rect 2780 27820 2832 27872
rect 3424 27863 3476 27872
rect 3424 27829 3433 27863
rect 3433 27829 3467 27863
rect 3467 27829 3476 27863
rect 3424 27820 3476 27829
rect 5172 27863 5224 27872
rect 5172 27829 5181 27863
rect 5181 27829 5215 27863
rect 5215 27829 5224 27863
rect 5172 27820 5224 27829
rect 8576 27820 8628 27872
rect 9680 27863 9732 27872
rect 9680 27829 9689 27863
rect 9689 27829 9723 27863
rect 9723 27829 9732 27863
rect 9680 27820 9732 27829
rect 10968 27820 11020 27872
rect 13544 27863 13596 27872
rect 13544 27829 13553 27863
rect 13553 27829 13587 27863
rect 13587 27829 13596 27863
rect 13544 27820 13596 27829
rect 15752 27863 15804 27872
rect 15752 27829 15761 27863
rect 15761 27829 15795 27863
rect 15795 27829 15804 27863
rect 15752 27820 15804 27829
rect 54852 27888 54904 27940
rect 19432 27820 19484 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 6000 27616 6052 27668
rect 2780 27523 2832 27532
rect 2780 27489 2789 27523
rect 2789 27489 2823 27523
rect 2823 27489 2832 27523
rect 2780 27480 2832 27489
rect 3056 27480 3108 27532
rect 4068 27480 4120 27532
rect 8116 27548 8168 27600
rect 10416 27548 10468 27600
rect 1952 27412 2004 27464
rect 2044 27412 2096 27464
rect 3240 27344 3292 27396
rect 3884 27412 3936 27464
rect 5172 27455 5224 27464
rect 5172 27421 5181 27455
rect 5181 27421 5215 27455
rect 5215 27421 5224 27455
rect 5172 27412 5224 27421
rect 5356 27412 5408 27464
rect 9128 27412 9180 27464
rect 9864 27344 9916 27396
rect 11336 27523 11388 27532
rect 11336 27489 11345 27523
rect 11345 27489 11379 27523
rect 11379 27489 11388 27523
rect 11336 27480 11388 27489
rect 13544 27548 13596 27600
rect 57704 27591 57756 27600
rect 57704 27557 57713 27591
rect 57713 27557 57747 27591
rect 57747 27557 57756 27591
rect 57704 27548 57756 27557
rect 15108 27480 15160 27532
rect 57152 27523 57204 27532
rect 57152 27489 57161 27523
rect 57161 27489 57195 27523
rect 57195 27489 57204 27523
rect 57152 27480 57204 27489
rect 57244 27480 57296 27532
rect 57612 27480 57664 27532
rect 58348 27523 58400 27532
rect 58348 27489 58357 27523
rect 58357 27489 58391 27523
rect 58391 27489 58400 27523
rect 58348 27480 58400 27489
rect 11060 27412 11112 27464
rect 58164 27455 58216 27464
rect 10784 27344 10836 27396
rect 58164 27421 58173 27455
rect 58173 27421 58207 27455
rect 58207 27421 58216 27455
rect 58164 27412 58216 27421
rect 17224 27344 17276 27396
rect 19248 27344 19300 27396
rect 1676 27319 1728 27328
rect 1676 27285 1685 27319
rect 1685 27285 1719 27319
rect 1719 27285 1728 27319
rect 1676 27276 1728 27285
rect 3332 27319 3384 27328
rect 3332 27285 3341 27319
rect 3341 27285 3375 27319
rect 3375 27285 3384 27319
rect 3332 27276 3384 27285
rect 5448 27276 5500 27328
rect 9036 27276 9088 27328
rect 10876 27276 10928 27328
rect 11060 27319 11112 27328
rect 11060 27285 11069 27319
rect 11069 27285 11103 27319
rect 11103 27285 11112 27319
rect 11060 27276 11112 27285
rect 12256 27276 12308 27328
rect 12992 27276 13044 27328
rect 14280 27319 14332 27328
rect 14280 27285 14289 27319
rect 14289 27285 14323 27319
rect 14323 27285 14332 27319
rect 14280 27276 14332 27285
rect 14924 27276 14976 27328
rect 18052 27276 18104 27328
rect 56508 27319 56560 27328
rect 56508 27285 56517 27319
rect 56517 27285 56551 27319
rect 56551 27285 56560 27319
rect 56508 27276 56560 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 2320 27072 2372 27124
rect 6644 27072 6696 27124
rect 11060 27072 11112 27124
rect 15108 27115 15160 27124
rect 15108 27081 15117 27115
rect 15117 27081 15151 27115
rect 15151 27081 15160 27115
rect 15108 27072 15160 27081
rect 18236 27072 18288 27124
rect 57152 27072 57204 27124
rect 57704 27072 57756 27124
rect 59452 27072 59504 27124
rect 5816 27004 5868 27056
rect 10968 27004 11020 27056
rect 11336 27004 11388 27056
rect 18052 27004 18104 27056
rect 2320 26936 2372 26988
rect 3240 26936 3292 26988
rect 3332 26936 3384 26988
rect 4804 26936 4856 26988
rect 9772 26936 9824 26988
rect 9956 26979 10008 26988
rect 9956 26945 9965 26979
rect 9965 26945 9999 26979
rect 9999 26945 10008 26979
rect 9956 26936 10008 26945
rect 12256 26979 12308 26988
rect 12256 26945 12265 26979
rect 12265 26945 12299 26979
rect 12299 26945 12308 26979
rect 12256 26936 12308 26945
rect 14280 26936 14332 26988
rect 58348 26979 58400 26988
rect 2688 26868 2740 26920
rect 5356 26911 5408 26920
rect 5356 26877 5365 26911
rect 5365 26877 5399 26911
rect 5399 26877 5408 26911
rect 5356 26868 5408 26877
rect 7656 26868 7708 26920
rect 12164 26868 12216 26920
rect 12992 26868 13044 26920
rect 16212 26868 16264 26920
rect 18052 26868 18104 26920
rect 13360 26800 13412 26852
rect 2872 26775 2924 26784
rect 2872 26741 2881 26775
rect 2881 26741 2915 26775
rect 2915 26741 2924 26775
rect 2872 26732 2924 26741
rect 3332 26732 3384 26784
rect 4712 26732 4764 26784
rect 6000 26775 6052 26784
rect 6000 26741 6009 26775
rect 6009 26741 6043 26775
rect 6043 26741 6052 26775
rect 6000 26732 6052 26741
rect 9128 26732 9180 26784
rect 10692 26732 10744 26784
rect 13452 26732 13504 26784
rect 17040 26732 17092 26784
rect 58348 26945 58357 26979
rect 58357 26945 58391 26979
rect 58391 26945 58400 26979
rect 58348 26936 58400 26945
rect 18512 26732 18564 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2136 26528 2188 26580
rect 5632 26460 5684 26512
rect 2320 26435 2372 26444
rect 2320 26401 2329 26435
rect 2329 26401 2363 26435
rect 2363 26401 2372 26435
rect 2320 26392 2372 26401
rect 2504 26435 2556 26444
rect 2504 26401 2513 26435
rect 2513 26401 2547 26435
rect 2547 26401 2556 26435
rect 2504 26392 2556 26401
rect 2780 26392 2832 26444
rect 5356 26392 5408 26444
rect 8392 26528 8444 26580
rect 12348 26528 12400 26580
rect 58348 26528 58400 26580
rect 2688 26324 2740 26376
rect 6368 26460 6420 26512
rect 7656 26460 7708 26512
rect 11428 26460 11480 26512
rect 10416 26392 10468 26444
rect 10876 26367 10928 26376
rect 5540 26256 5592 26308
rect 6368 26256 6420 26308
rect 2688 26188 2740 26240
rect 2964 26231 3016 26240
rect 2964 26197 2973 26231
rect 2973 26197 3007 26231
rect 3007 26197 3016 26231
rect 10876 26333 10885 26367
rect 10885 26333 10919 26367
rect 10919 26333 10928 26367
rect 10876 26324 10928 26333
rect 43720 26460 43772 26512
rect 57612 26503 57664 26512
rect 57612 26469 57621 26503
rect 57621 26469 57655 26503
rect 57655 26469 57664 26503
rect 57612 26460 57664 26469
rect 58072 26460 58124 26512
rect 18236 26392 18288 26444
rect 18512 26324 18564 26376
rect 56508 26324 56560 26376
rect 57520 26324 57572 26376
rect 58348 26367 58400 26376
rect 58348 26333 58357 26367
rect 58357 26333 58391 26367
rect 58391 26333 58400 26367
rect 58348 26324 58400 26333
rect 8392 26256 8444 26308
rect 9772 26256 9824 26308
rect 9956 26299 10008 26308
rect 9956 26265 9965 26299
rect 9965 26265 9999 26299
rect 9999 26265 10008 26299
rect 9956 26256 10008 26265
rect 11152 26256 11204 26308
rect 12164 26256 12216 26308
rect 17960 26256 18012 26308
rect 2964 26188 3016 26197
rect 16580 26231 16632 26240
rect 16580 26197 16589 26231
rect 16589 26197 16623 26231
rect 16623 26197 16632 26231
rect 16580 26188 16632 26197
rect 18512 26188 18564 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 1676 26027 1728 26036
rect 1676 25993 1685 26027
rect 1685 25993 1719 26027
rect 1719 25993 1728 26027
rect 1676 25984 1728 25993
rect 2136 25984 2188 26036
rect 2320 26027 2372 26036
rect 2320 25993 2329 26027
rect 2329 25993 2363 26027
rect 2363 25993 2372 26027
rect 2320 25984 2372 25993
rect 2688 25984 2740 26036
rect 3240 25984 3292 26036
rect 3332 25984 3384 26036
rect 5356 25984 5408 26036
rect 57520 26027 57572 26036
rect 57520 25993 57529 26027
rect 57529 25993 57563 26027
rect 57563 25993 57572 26027
rect 57520 25984 57572 25993
rect 18512 25916 18564 25968
rect 2044 25848 2096 25900
rect 2872 25891 2924 25900
rect 2872 25857 2881 25891
rect 2881 25857 2915 25891
rect 2915 25857 2924 25891
rect 2872 25848 2924 25857
rect 6000 25848 6052 25900
rect 12348 25848 12400 25900
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 18328 25848 18380 25900
rect 58348 25891 58400 25900
rect 58348 25857 58357 25891
rect 58357 25857 58391 25891
rect 58391 25857 58400 25891
rect 58348 25848 58400 25857
rect 19432 25780 19484 25832
rect 6368 25712 6420 25764
rect 9220 25712 9272 25764
rect 14096 25712 14148 25764
rect 3056 25687 3108 25696
rect 3056 25653 3065 25687
rect 3065 25653 3099 25687
rect 3099 25653 3108 25687
rect 3056 25644 3108 25653
rect 3240 25644 3292 25696
rect 4804 25644 4856 25696
rect 6828 25644 6880 25696
rect 10416 25644 10468 25696
rect 14188 25644 14240 25696
rect 16856 25687 16908 25696
rect 16856 25653 16865 25687
rect 16865 25653 16899 25687
rect 16899 25653 16908 25687
rect 16856 25644 16908 25653
rect 18236 25644 18288 25696
rect 18512 25687 18564 25696
rect 18512 25653 18521 25687
rect 18521 25653 18555 25687
rect 18555 25653 18564 25687
rect 18512 25644 18564 25653
rect 19616 25644 19668 25696
rect 55864 25712 55916 25764
rect 20352 25644 20404 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1676 25483 1728 25492
rect 1676 25449 1685 25483
rect 1685 25449 1719 25483
rect 1719 25449 1728 25483
rect 1676 25440 1728 25449
rect 8300 25440 8352 25492
rect 9680 25440 9732 25492
rect 57428 25440 57480 25492
rect 58808 25440 58860 25492
rect 2596 25372 2648 25424
rect 2412 25236 2464 25288
rect 2964 25279 3016 25288
rect 2964 25245 2973 25279
rect 2973 25245 3007 25279
rect 3007 25245 3016 25279
rect 2964 25236 3016 25245
rect 5724 25304 5776 25356
rect 2044 25168 2096 25220
rect 6000 25168 6052 25220
rect 6920 25168 6972 25220
rect 16856 25304 16908 25356
rect 57796 25372 57848 25424
rect 57704 25347 57756 25356
rect 57704 25313 57713 25347
rect 57713 25313 57747 25347
rect 57747 25313 57756 25347
rect 57704 25304 57756 25313
rect 58532 25304 58584 25356
rect 15384 25236 15436 25288
rect 19616 25279 19668 25288
rect 19616 25245 19625 25279
rect 19625 25245 19659 25279
rect 19659 25245 19668 25279
rect 19616 25236 19668 25245
rect 57152 25279 57204 25288
rect 57152 25245 57161 25279
rect 57161 25245 57195 25279
rect 57195 25245 57204 25279
rect 57428 25279 57480 25288
rect 57152 25236 57204 25245
rect 57428 25245 57437 25279
rect 57437 25245 57471 25279
rect 57471 25245 57480 25279
rect 57428 25236 57480 25245
rect 58164 25279 58216 25288
rect 58164 25245 58173 25279
rect 58173 25245 58207 25279
rect 58207 25245 58216 25279
rect 58164 25236 58216 25245
rect 11796 25168 11848 25220
rect 12072 25168 12124 25220
rect 16212 25100 16264 25152
rect 18328 25100 18380 25152
rect 18696 25100 18748 25152
rect 56508 25143 56560 25152
rect 56508 25109 56517 25143
rect 56517 25109 56551 25143
rect 56551 25109 56560 25143
rect 56508 25100 56560 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 4988 24828 5040 24880
rect 14832 24828 14884 24880
rect 3700 24760 3752 24812
rect 5724 24803 5776 24812
rect 5724 24769 5733 24803
rect 5733 24769 5767 24803
rect 5767 24769 5776 24803
rect 5724 24760 5776 24769
rect 6920 24760 6972 24812
rect 8208 24760 8260 24812
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 15384 24760 15436 24769
rect 19616 24760 19668 24812
rect 58348 24803 58400 24812
rect 58348 24769 58357 24803
rect 58357 24769 58391 24803
rect 58391 24769 58400 24803
rect 58348 24760 58400 24769
rect 2504 24692 2556 24744
rect 8392 24692 8444 24744
rect 9772 24735 9824 24744
rect 9772 24701 9781 24735
rect 9781 24701 9815 24735
rect 9815 24701 9824 24735
rect 9772 24692 9824 24701
rect 10048 24735 10100 24744
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 18696 24692 18748 24744
rect 1676 24667 1728 24676
rect 1676 24633 1685 24667
rect 1685 24633 1719 24667
rect 1719 24633 1728 24667
rect 1676 24624 1728 24633
rect 1860 24624 1912 24676
rect 17224 24624 17276 24676
rect 58072 24624 58124 24676
rect 2412 24599 2464 24608
rect 2412 24565 2421 24599
rect 2421 24565 2455 24599
rect 2455 24565 2464 24599
rect 2412 24556 2464 24565
rect 3516 24599 3568 24608
rect 3516 24565 3525 24599
rect 3525 24565 3559 24599
rect 3559 24565 3568 24599
rect 3516 24556 3568 24565
rect 4068 24556 4120 24608
rect 9220 24556 9272 24608
rect 13636 24599 13688 24608
rect 13636 24565 13645 24599
rect 13645 24565 13679 24599
rect 13679 24565 13688 24599
rect 13636 24556 13688 24565
rect 18328 24556 18380 24608
rect 18788 24556 18840 24608
rect 19340 24556 19392 24608
rect 57152 24556 57204 24608
rect 57244 24556 57296 24608
rect 57704 24556 57756 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3516 24352 3568 24404
rect 2780 24259 2832 24268
rect 2780 24225 2789 24259
rect 2789 24225 2823 24259
rect 2823 24225 2832 24259
rect 2780 24216 2832 24225
rect 3424 24216 3476 24268
rect 3700 24284 3752 24336
rect 6092 24284 6144 24336
rect 11980 24352 12032 24404
rect 18052 24352 18104 24404
rect 19616 24395 19668 24404
rect 19616 24361 19625 24395
rect 19625 24361 19659 24395
rect 19659 24361 19668 24395
rect 19616 24352 19668 24361
rect 58348 24352 58400 24404
rect 14924 24284 14976 24336
rect 57060 24284 57112 24336
rect 10048 24216 10100 24268
rect 10692 24259 10744 24268
rect 10692 24225 10701 24259
rect 10701 24225 10735 24259
rect 10735 24225 10744 24259
rect 10692 24216 10744 24225
rect 20260 24259 20312 24268
rect 20260 24225 20269 24259
rect 20269 24225 20303 24259
rect 20303 24225 20312 24259
rect 20260 24216 20312 24225
rect 11796 24148 11848 24200
rect 13912 24148 13964 24200
rect 18788 24191 18840 24200
rect 18788 24157 18797 24191
rect 18797 24157 18831 24191
rect 18831 24157 18840 24191
rect 18788 24148 18840 24157
rect 58348 24191 58400 24200
rect 58348 24157 58357 24191
rect 58357 24157 58391 24191
rect 58391 24157 58400 24191
rect 58348 24148 58400 24157
rect 3700 24080 3752 24132
rect 19340 24080 19392 24132
rect 1676 24055 1728 24064
rect 1676 24021 1685 24055
rect 1685 24021 1719 24055
rect 1719 24021 1728 24055
rect 1676 24012 1728 24021
rect 3424 24055 3476 24064
rect 3424 24021 3433 24055
rect 3433 24021 3467 24055
rect 3467 24021 3476 24055
rect 3424 24012 3476 24021
rect 3516 24012 3568 24064
rect 3976 24012 4028 24064
rect 5172 24012 5224 24064
rect 19984 24055 20036 24064
rect 19984 24021 19993 24055
rect 19993 24021 20027 24055
rect 20027 24021 20036 24055
rect 19984 24012 20036 24021
rect 20260 24012 20312 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 2780 23808 2832 23860
rect 19984 23808 20036 23860
rect 58808 23808 58860 23860
rect 2044 23740 2096 23792
rect 2412 23740 2464 23792
rect 14280 23740 14332 23792
rect 2780 23672 2832 23724
rect 4896 23672 4948 23724
rect 6184 23672 6236 23724
rect 19432 23672 19484 23724
rect 3976 23604 4028 23656
rect 5908 23604 5960 23656
rect 6092 23604 6144 23656
rect 2412 23536 2464 23588
rect 2320 23468 2372 23520
rect 17960 23536 18012 23588
rect 18604 23536 18656 23588
rect 10416 23468 10468 23520
rect 18420 23511 18472 23520
rect 18420 23477 18429 23511
rect 18429 23477 18463 23511
rect 18463 23477 18472 23511
rect 18420 23468 18472 23477
rect 20076 23468 20128 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 16028 23307 16080 23316
rect 16028 23273 16037 23307
rect 16037 23273 16071 23307
rect 16071 23273 16080 23307
rect 16028 23264 16080 23273
rect 19432 23307 19484 23316
rect 4896 23196 4948 23248
rect 16488 23128 16540 23180
rect 19432 23273 19441 23307
rect 19441 23273 19475 23307
rect 19475 23273 19484 23307
rect 19432 23264 19484 23273
rect 58716 23264 58768 23316
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 3424 23060 3476 23112
rect 58348 23103 58400 23112
rect 58348 23069 58357 23103
rect 58357 23069 58391 23103
rect 58391 23069 58400 23103
rect 58348 23060 58400 23069
rect 9956 22992 10008 23044
rect 10876 22992 10928 23044
rect 14832 22992 14884 23044
rect 18420 22992 18472 23044
rect 1676 22967 1728 22976
rect 1676 22933 1685 22967
rect 1685 22933 1719 22967
rect 1719 22933 1728 22967
rect 1676 22924 1728 22933
rect 2780 22924 2832 22976
rect 3976 22924 4028 22976
rect 4804 22924 4856 22976
rect 19984 22924 20036 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2780 22720 2832 22772
rect 3700 22763 3752 22772
rect 3700 22729 3709 22763
rect 3709 22729 3743 22763
rect 3743 22729 3752 22763
rect 3700 22720 3752 22729
rect 8484 22720 8536 22772
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 56140 22720 56192 22772
rect 2596 22652 2648 22704
rect 2136 22559 2188 22568
rect 2136 22525 2145 22559
rect 2145 22525 2179 22559
rect 2179 22525 2188 22559
rect 2136 22516 2188 22525
rect 2596 22380 2648 22432
rect 8392 22652 8444 22704
rect 13912 22652 13964 22704
rect 10048 22627 10100 22636
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 58348 22627 58400 22636
rect 58348 22593 58357 22627
rect 58357 22593 58391 22627
rect 58391 22593 58400 22627
rect 58348 22584 58400 22593
rect 8760 22516 8812 22568
rect 15384 22516 15436 22568
rect 16488 22516 16540 22568
rect 16580 22448 16632 22500
rect 19432 22516 19484 22568
rect 18144 22448 18196 22500
rect 10416 22380 10468 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1676 22219 1728 22228
rect 1676 22185 1685 22219
rect 1685 22185 1719 22219
rect 1719 22185 1728 22219
rect 1676 22176 1728 22185
rect 8576 22176 8628 22228
rect 16304 22176 16356 22228
rect 18144 22176 18196 22228
rect 19432 22176 19484 22228
rect 2136 22040 2188 22092
rect 2688 22040 2740 22092
rect 7104 22040 7156 22092
rect 15384 22040 15436 22092
rect 20076 22040 20128 22092
rect 20628 22040 20680 22092
rect 56508 22040 56560 22092
rect 19156 21972 19208 22024
rect 20168 21972 20220 22024
rect 57980 22015 58032 22024
rect 57980 21981 57989 22015
rect 57989 21981 58023 22015
rect 58023 21981 58032 22015
rect 57980 21972 58032 21981
rect 10692 21904 10744 21956
rect 12348 21836 12400 21888
rect 16212 21904 16264 21956
rect 14832 21836 14884 21888
rect 20628 21836 20680 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 19064 21632 19116 21684
rect 58164 21675 58216 21684
rect 58164 21641 58173 21675
rect 58173 21641 58207 21675
rect 58207 21641 58216 21675
rect 58164 21632 58216 21641
rect 2412 21564 2464 21616
rect 15384 21564 15436 21616
rect 3240 21496 3292 21548
rect 12440 21496 12492 21548
rect 18696 21496 18748 21548
rect 58348 21539 58400 21548
rect 58348 21505 58357 21539
rect 58357 21505 58391 21539
rect 58391 21505 58400 21539
rect 58348 21496 58400 21505
rect 2228 21471 2280 21480
rect 2228 21437 2237 21471
rect 2237 21437 2271 21471
rect 2271 21437 2280 21471
rect 2228 21428 2280 21437
rect 1952 21360 2004 21412
rect 14372 21360 14424 21412
rect 2320 21292 2372 21344
rect 3240 21335 3292 21344
rect 3240 21301 3249 21335
rect 3249 21301 3283 21335
rect 3283 21301 3292 21335
rect 3240 21292 3292 21301
rect 12440 21335 12492 21344
rect 12440 21301 12449 21335
rect 12449 21301 12483 21335
rect 12483 21301 12492 21335
rect 12440 21292 12492 21301
rect 18696 21292 18748 21344
rect 18972 21335 19024 21344
rect 18972 21301 18981 21335
rect 18981 21301 19015 21335
rect 19015 21301 19024 21335
rect 18972 21292 19024 21301
rect 20260 21335 20312 21344
rect 20260 21301 20269 21335
rect 20269 21301 20303 21335
rect 20303 21301 20312 21335
rect 20260 21292 20312 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1676 21131 1728 21140
rect 1676 21097 1685 21131
rect 1685 21097 1719 21131
rect 1719 21097 1728 21131
rect 1676 21088 1728 21097
rect 2228 21088 2280 21140
rect 5816 21088 5868 21140
rect 8300 21131 8352 21140
rect 8300 21097 8321 21131
rect 8321 21097 8352 21131
rect 14372 21131 14424 21140
rect 8300 21088 8352 21097
rect 14372 21097 14381 21131
rect 14381 21097 14415 21131
rect 14415 21097 14424 21131
rect 14372 21088 14424 21097
rect 18880 21088 18932 21140
rect 19064 21088 19116 21140
rect 58256 21088 58308 21140
rect 5724 20995 5776 21004
rect 5724 20961 5733 20995
rect 5733 20961 5767 20995
rect 5767 20961 5776 20995
rect 5724 20952 5776 20961
rect 8300 20952 8352 21004
rect 10048 20952 10100 21004
rect 15384 20952 15436 21004
rect 16120 20995 16172 21004
rect 16120 20961 16129 20995
rect 16129 20961 16163 20995
rect 16163 20961 16172 20995
rect 16120 20952 16172 20961
rect 2044 20884 2096 20936
rect 2320 20927 2372 20936
rect 2320 20893 2329 20927
rect 2329 20893 2363 20927
rect 2363 20893 2372 20927
rect 2320 20884 2372 20893
rect 2412 20884 2464 20936
rect 58348 20927 58400 20936
rect 58348 20893 58357 20927
rect 58357 20893 58391 20927
rect 58391 20893 58400 20927
rect 58348 20884 58400 20893
rect 1952 20816 2004 20868
rect 4988 20816 5040 20868
rect 14832 20816 14884 20868
rect 16948 20816 17000 20868
rect 8392 20748 8444 20800
rect 11888 20791 11940 20800
rect 11888 20757 11897 20791
rect 11897 20757 11931 20791
rect 11931 20757 11940 20791
rect 11888 20748 11940 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 2688 20544 2740 20596
rect 8300 20587 8352 20596
rect 8300 20553 8309 20587
rect 8309 20553 8343 20587
rect 8343 20553 8352 20587
rect 8300 20544 8352 20553
rect 14280 20587 14332 20596
rect 14280 20553 14289 20587
rect 14289 20553 14323 20587
rect 14323 20553 14332 20587
rect 14280 20544 14332 20553
rect 4988 20519 5040 20528
rect 4988 20485 4997 20519
rect 4997 20485 5031 20519
rect 5031 20485 5040 20519
rect 4988 20476 5040 20485
rect 2228 20408 2280 20460
rect 5816 20408 5868 20460
rect 5816 20247 5868 20256
rect 5816 20213 5825 20247
rect 5825 20213 5859 20247
rect 5859 20213 5868 20247
rect 11888 20476 11940 20528
rect 12348 20519 12400 20528
rect 12348 20485 12357 20519
rect 12357 20485 12391 20519
rect 12391 20485 12400 20519
rect 12348 20476 12400 20485
rect 13912 20476 13964 20528
rect 18696 20476 18748 20528
rect 20352 20519 20404 20528
rect 20352 20485 20361 20519
rect 20361 20485 20395 20519
rect 20395 20485 20404 20519
rect 20352 20476 20404 20485
rect 16120 20408 16172 20460
rect 18972 20408 19024 20460
rect 20628 20451 20680 20460
rect 20628 20417 20637 20451
rect 20637 20417 20671 20451
rect 20671 20417 20680 20451
rect 20628 20408 20680 20417
rect 17316 20340 17368 20392
rect 12440 20272 12492 20324
rect 19432 20383 19484 20392
rect 19432 20349 19441 20383
rect 19441 20349 19475 20383
rect 19475 20349 19484 20383
rect 19432 20340 19484 20349
rect 5816 20204 5868 20213
rect 14372 20204 14424 20256
rect 17224 20204 17276 20256
rect 17592 20247 17644 20256
rect 17592 20213 17601 20247
rect 17601 20213 17635 20247
rect 17635 20213 17644 20247
rect 17592 20204 17644 20213
rect 18052 20204 18104 20256
rect 18788 20247 18840 20256
rect 18788 20213 18797 20247
rect 18797 20213 18831 20247
rect 18831 20213 18840 20247
rect 18788 20204 18840 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2688 19864 2740 19916
rect 6184 19932 6236 19984
rect 12624 19975 12676 19984
rect 12624 19941 12633 19975
rect 12633 19941 12667 19975
rect 12667 19941 12676 19975
rect 12624 19932 12676 19941
rect 8300 19864 8352 19916
rect 10048 19864 10100 19916
rect 11244 19864 11296 19916
rect 12348 19864 12400 19916
rect 19340 19864 19392 19916
rect 3884 19796 3936 19848
rect 4988 19796 5040 19848
rect 58348 19839 58400 19848
rect 58348 19805 58357 19839
rect 58357 19805 58391 19839
rect 58391 19805 58400 19839
rect 58348 19796 58400 19805
rect 2136 19728 2188 19780
rect 2412 19660 2464 19712
rect 4988 19660 5040 19712
rect 14372 19660 14424 19712
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 19432 19660 19484 19712
rect 20168 19660 20220 19712
rect 58624 19660 58676 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 1676 19499 1728 19508
rect 1676 19465 1685 19499
rect 1685 19465 1719 19499
rect 1719 19465 1728 19499
rect 1676 19456 1728 19465
rect 10508 19499 10560 19508
rect 10508 19465 10517 19499
rect 10517 19465 10551 19499
rect 10551 19465 10560 19499
rect 10508 19456 10560 19465
rect 10876 19456 10928 19508
rect 13820 19456 13872 19508
rect 8208 19388 8260 19440
rect 13912 19388 13964 19440
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 3148 19252 3200 19304
rect 3884 19252 3936 19304
rect 7656 19252 7708 19304
rect 8300 19320 8352 19372
rect 15384 19320 15436 19372
rect 58440 19456 58492 19508
rect 19340 19320 19392 19372
rect 58348 19363 58400 19372
rect 9036 19295 9088 19304
rect 9036 19261 9045 19295
rect 9045 19261 9079 19295
rect 9079 19261 9088 19295
rect 9036 19252 9088 19261
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 58348 19329 58357 19363
rect 58357 19329 58391 19363
rect 58391 19329 58400 19363
rect 58348 19320 58400 19329
rect 18144 19159 18196 19168
rect 18144 19125 18153 19159
rect 18153 19125 18187 19159
rect 18187 19125 18196 19159
rect 19984 19252 20036 19304
rect 20260 19184 20312 19236
rect 18144 19116 18196 19125
rect 20628 19116 20680 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1676 18955 1728 18964
rect 1676 18921 1685 18955
rect 1685 18921 1719 18955
rect 1719 18921 1728 18955
rect 1676 18912 1728 18921
rect 2504 18955 2556 18964
rect 2504 18921 2513 18955
rect 2513 18921 2547 18955
rect 2547 18921 2556 18955
rect 2504 18912 2556 18921
rect 3332 18912 3384 18964
rect 16948 18955 17000 18964
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 58348 18955 58400 18964
rect 58348 18921 58357 18955
rect 58357 18921 58391 18955
rect 58391 18921 58400 18955
rect 58348 18912 58400 18921
rect 3608 18776 3660 18828
rect 18144 18776 18196 18828
rect 18236 18776 18288 18828
rect 2228 18708 2280 18760
rect 2412 18708 2464 18760
rect 5264 18708 5316 18760
rect 15844 18708 15896 18760
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 18788 18708 18840 18760
rect 20536 18776 20588 18828
rect 6000 18640 6052 18692
rect 11520 18640 11572 18692
rect 18696 18640 18748 18692
rect 20260 18640 20312 18692
rect 6828 18572 6880 18624
rect 8116 18572 8168 18624
rect 17040 18572 17092 18624
rect 19432 18615 19484 18624
rect 19432 18581 19441 18615
rect 19441 18581 19475 18615
rect 19475 18581 19484 18615
rect 19432 18572 19484 18581
rect 19984 18572 20036 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 1860 18368 1912 18420
rect 2412 18411 2464 18420
rect 2412 18377 2421 18411
rect 2421 18377 2455 18411
rect 2455 18377 2464 18411
rect 2412 18368 2464 18377
rect 6644 18411 6696 18420
rect 6644 18377 6653 18411
rect 6653 18377 6687 18411
rect 6687 18377 6696 18411
rect 6644 18368 6696 18377
rect 6736 18368 6788 18420
rect 13820 18368 13872 18420
rect 17132 18368 17184 18420
rect 19340 18368 19392 18420
rect 19524 18368 19576 18420
rect 3332 18300 3384 18352
rect 7656 18300 7708 18352
rect 8116 18343 8168 18352
rect 8116 18309 8125 18343
rect 8125 18309 8159 18343
rect 8159 18309 8168 18343
rect 8116 18300 8168 18309
rect 14464 18300 14516 18352
rect 5540 18232 5592 18284
rect 7104 18232 7156 18284
rect 18144 18232 18196 18284
rect 58348 18275 58400 18284
rect 58348 18241 58357 18275
rect 58357 18241 58391 18275
rect 58391 18241 58400 18275
rect 58348 18232 58400 18241
rect 1952 18164 2004 18216
rect 3608 18164 3660 18216
rect 5908 18164 5960 18216
rect 8668 18164 8720 18216
rect 19340 18164 19392 18216
rect 20536 18164 20588 18216
rect 6736 18096 6788 18148
rect 17316 18139 17368 18148
rect 17316 18105 17325 18139
rect 17325 18105 17359 18139
rect 17359 18105 17368 18139
rect 17316 18096 17368 18105
rect 7104 18028 7156 18080
rect 7656 18028 7708 18080
rect 20260 18028 20312 18080
rect 58808 18028 58860 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1676 17867 1728 17876
rect 1676 17833 1685 17867
rect 1685 17833 1719 17867
rect 1719 17833 1728 17867
rect 1676 17824 1728 17833
rect 1952 17824 2004 17876
rect 9864 17824 9916 17876
rect 11980 17824 12032 17876
rect 17592 17824 17644 17876
rect 18144 17867 18196 17876
rect 18144 17833 18153 17867
rect 18153 17833 18187 17867
rect 18187 17833 18196 17867
rect 18144 17824 18196 17833
rect 19524 17867 19576 17876
rect 19524 17833 19533 17867
rect 19533 17833 19567 17867
rect 19567 17833 19576 17867
rect 19524 17824 19576 17833
rect 20444 17824 20496 17876
rect 11428 17688 11480 17740
rect 15200 17731 15252 17740
rect 15200 17697 15209 17731
rect 15209 17697 15243 17731
rect 15243 17697 15252 17731
rect 15200 17688 15252 17697
rect 18512 17688 18564 17740
rect 19340 17688 19392 17740
rect 2504 17620 2556 17672
rect 2688 17620 2740 17672
rect 13820 17620 13872 17672
rect 17224 17663 17276 17672
rect 17224 17629 17233 17663
rect 17233 17629 17267 17663
rect 17267 17629 17276 17663
rect 17224 17620 17276 17629
rect 7656 17552 7708 17604
rect 9680 17552 9732 17604
rect 13912 17552 13964 17604
rect 15016 17552 15068 17604
rect 17776 17552 17828 17604
rect 2412 17527 2464 17536
rect 2412 17493 2421 17527
rect 2421 17493 2455 17527
rect 2455 17493 2464 17527
rect 2412 17484 2464 17493
rect 14280 17484 14332 17536
rect 17592 17484 17644 17536
rect 19156 17620 19208 17672
rect 58348 17663 58400 17672
rect 58348 17629 58357 17663
rect 58357 17629 58391 17663
rect 58391 17629 58400 17663
rect 58348 17620 58400 17629
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 58256 17484 58308 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 2780 17280 2832 17332
rect 7748 17280 7800 17332
rect 11980 17323 12032 17332
rect 11980 17289 11989 17323
rect 11989 17289 12023 17323
rect 12023 17289 12032 17323
rect 11980 17280 12032 17289
rect 13820 17280 13872 17332
rect 2688 17212 2740 17264
rect 8392 17212 8444 17264
rect 13912 17212 13964 17264
rect 1952 17076 2004 17128
rect 5816 17144 5868 17196
rect 6368 17144 6420 17196
rect 13820 17144 13872 17196
rect 17224 17280 17276 17332
rect 17592 17280 17644 17332
rect 18604 17280 18656 17332
rect 18972 17280 19024 17332
rect 19156 17280 19208 17332
rect 19432 17144 19484 17196
rect 5540 17119 5592 17128
rect 5540 17085 5549 17119
rect 5549 17085 5583 17119
rect 5583 17085 5592 17119
rect 5540 17076 5592 17085
rect 9404 17008 9456 17060
rect 14096 17008 14148 17060
rect 4804 16940 4856 16992
rect 5080 16940 5132 16992
rect 6368 16940 6420 16992
rect 17684 17076 17736 17128
rect 17316 17008 17368 17060
rect 17040 16940 17092 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1952 16736 2004 16788
rect 2688 16736 2740 16788
rect 13084 16736 13136 16788
rect 17316 16736 17368 16788
rect 17776 16779 17828 16788
rect 17776 16745 17785 16779
rect 17785 16745 17819 16779
rect 17819 16745 17828 16779
rect 17776 16736 17828 16745
rect 5080 16600 5132 16652
rect 5908 16643 5960 16652
rect 5908 16609 5917 16643
rect 5917 16609 5951 16643
rect 5951 16609 5960 16643
rect 5908 16600 5960 16609
rect 14096 16600 14148 16652
rect 18512 16600 18564 16652
rect 1860 16575 1912 16584
rect 1860 16541 1869 16575
rect 1869 16541 1903 16575
rect 1903 16541 1912 16575
rect 1860 16532 1912 16541
rect 2320 16532 2372 16584
rect 2688 16532 2740 16584
rect 18788 16532 18840 16584
rect 58348 16575 58400 16584
rect 58348 16541 58357 16575
rect 58357 16541 58391 16575
rect 58391 16541 58400 16575
rect 58348 16532 58400 16541
rect 5540 16464 5592 16516
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 2504 16396 2556 16448
rect 2688 16396 2740 16448
rect 5264 16396 5316 16448
rect 58808 16396 58860 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 2688 16192 2740 16244
rect 6552 16192 6604 16244
rect 6736 16192 6788 16244
rect 10416 16235 10468 16244
rect 2044 16056 2096 16108
rect 4620 15988 4672 16040
rect 10416 16201 10425 16235
rect 10425 16201 10459 16235
rect 10459 16201 10468 16235
rect 10416 16192 10468 16201
rect 17684 16192 17736 16244
rect 18788 16235 18840 16244
rect 18788 16201 18797 16235
rect 18797 16201 18831 16235
rect 18831 16201 18840 16235
rect 18788 16192 18840 16201
rect 16304 16124 16356 16176
rect 10048 16056 10100 16108
rect 12808 16056 12860 16108
rect 19340 16124 19392 16176
rect 20168 16056 20220 16108
rect 58348 16099 58400 16108
rect 58348 16065 58357 16099
rect 58357 16065 58391 16099
rect 58391 16065 58400 16099
rect 58348 16056 58400 16065
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 9680 15988 9732 16040
rect 18604 15988 18656 16040
rect 19432 16031 19484 16040
rect 19432 15997 19441 16031
rect 19441 15997 19475 16031
rect 19475 15997 19484 16031
rect 19432 15988 19484 15997
rect 19984 15988 20036 16040
rect 11520 15920 11572 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 1860 15852 1912 15904
rect 7656 15852 7708 15904
rect 12440 15852 12492 15904
rect 12808 15852 12860 15904
rect 13820 15852 13872 15904
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 14464 15852 14516 15861
rect 19432 15852 19484 15904
rect 20352 15852 20404 15904
rect 20628 15852 20680 15904
rect 57796 15852 57848 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2504 15648 2556 15700
rect 5632 15648 5684 15700
rect 2044 15623 2096 15632
rect 2044 15589 2053 15623
rect 2053 15589 2087 15623
rect 2087 15589 2096 15623
rect 8024 15648 8076 15700
rect 8392 15648 8444 15700
rect 18604 15691 18656 15700
rect 18604 15657 18613 15691
rect 18613 15657 18647 15691
rect 18647 15657 18656 15691
rect 18604 15648 18656 15657
rect 58348 15691 58400 15700
rect 58348 15657 58357 15691
rect 58357 15657 58391 15691
rect 58391 15657 58400 15691
rect 58348 15648 58400 15657
rect 2044 15580 2096 15589
rect 3056 15512 3108 15564
rect 9404 15555 9456 15564
rect 9404 15521 9413 15555
rect 9413 15521 9447 15555
rect 9447 15521 9456 15555
rect 9404 15512 9456 15521
rect 57244 15555 57296 15564
rect 57244 15521 57253 15555
rect 57253 15521 57287 15555
rect 57287 15521 57296 15555
rect 57244 15512 57296 15521
rect 8300 15444 8352 15496
rect 8668 15444 8720 15496
rect 19432 15444 19484 15496
rect 5540 15376 5592 15428
rect 10048 15376 10100 15428
rect 4896 15308 4948 15360
rect 7288 15308 7340 15360
rect 7564 15308 7616 15360
rect 12348 15308 12400 15360
rect 18696 15308 18748 15360
rect 20076 15351 20128 15360
rect 20076 15317 20085 15351
rect 20085 15317 20119 15351
rect 20119 15317 20128 15351
rect 20076 15308 20128 15317
rect 56416 15351 56468 15360
rect 56416 15317 56425 15351
rect 56425 15317 56459 15351
rect 56459 15317 56468 15351
rect 56416 15308 56468 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 12348 15147 12400 15156
rect 12348 15113 12357 15147
rect 12357 15113 12391 15147
rect 12391 15113 12400 15147
rect 12348 15104 12400 15113
rect 13820 15104 13872 15156
rect 18696 15104 18748 15156
rect 19432 15104 19484 15156
rect 2136 15036 2188 15088
rect 2504 15036 2556 15088
rect 15016 15036 15068 15088
rect 3148 14968 3200 15020
rect 2228 14943 2280 14952
rect 2228 14909 2237 14943
rect 2237 14909 2271 14943
rect 2271 14909 2280 14943
rect 2228 14900 2280 14909
rect 14372 14968 14424 15020
rect 13820 14943 13872 14952
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 13820 14900 13872 14909
rect 14464 14900 14516 14952
rect 19892 15036 19944 15088
rect 20168 15036 20220 15088
rect 12808 14832 12860 14884
rect 2688 14807 2740 14816
rect 2688 14773 2697 14807
rect 2697 14773 2731 14807
rect 2731 14773 2740 14807
rect 2688 14764 2740 14773
rect 3148 14807 3200 14816
rect 3148 14773 3157 14807
rect 3157 14773 3191 14807
rect 3191 14773 3200 14807
rect 3148 14764 3200 14773
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 5264 14764 5316 14816
rect 8300 14807 8352 14816
rect 8300 14773 8309 14807
rect 8309 14773 8343 14807
rect 8343 14773 8352 14807
rect 8300 14764 8352 14773
rect 17500 14764 17552 14816
rect 58348 15011 58400 15020
rect 58348 14977 58357 15011
rect 58357 14977 58391 15011
rect 58391 14977 58400 15011
rect 58348 14968 58400 14977
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 20628 14900 20680 14952
rect 19984 14764 20036 14816
rect 20628 14764 20680 14816
rect 57336 14764 57388 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 3792 14560 3844 14612
rect 5172 14560 5224 14612
rect 5264 14560 5316 14612
rect 13268 14560 13320 14612
rect 18512 14560 18564 14612
rect 2596 14492 2648 14544
rect 4620 14492 4672 14544
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 8300 14424 8352 14476
rect 19340 14560 19392 14612
rect 19892 14560 19944 14612
rect 19984 14467 20036 14476
rect 19984 14433 19993 14467
rect 19993 14433 20027 14467
rect 20027 14433 20036 14467
rect 19984 14424 20036 14433
rect 20536 14424 20588 14476
rect 12348 14356 12400 14408
rect 20076 14356 20128 14408
rect 20720 14356 20772 14408
rect 58348 14399 58400 14408
rect 58348 14365 58357 14399
rect 58357 14365 58391 14399
rect 58391 14365 58400 14399
rect 58348 14356 58400 14365
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 5172 14288 5224 14340
rect 9588 14331 9640 14340
rect 9588 14297 9597 14331
rect 9597 14297 9631 14331
rect 9631 14297 9640 14331
rect 9588 14288 9640 14297
rect 8944 14220 8996 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 11612 14288 11664 14340
rect 12624 14220 12676 14272
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 20076 14220 20128 14272
rect 58164 14263 58216 14272
rect 58164 14229 58173 14263
rect 58173 14229 58207 14263
rect 58207 14229 58216 14263
rect 58164 14220 58216 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 5264 14016 5316 14068
rect 16672 14016 16724 14068
rect 17500 14016 17552 14068
rect 20720 14059 20772 14068
rect 2780 13948 2832 14000
rect 3884 13991 3936 14000
rect 3884 13957 3893 13991
rect 3893 13957 3927 13991
rect 3927 13957 3936 13991
rect 3884 13948 3936 13957
rect 12624 13948 12676 14000
rect 20720 14025 20729 14059
rect 20729 14025 20763 14059
rect 20763 14025 20772 14059
rect 20720 14016 20772 14025
rect 57244 14016 57296 14068
rect 57704 14016 57756 14068
rect 58440 14016 58492 14068
rect 58992 14016 59044 14068
rect 2044 13880 2096 13932
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 2688 13880 2740 13932
rect 20076 13880 20128 13932
rect 11060 13812 11112 13864
rect 11612 13812 11664 13864
rect 15016 13855 15068 13864
rect 15016 13821 15025 13855
rect 15025 13821 15059 13855
rect 15059 13821 15068 13855
rect 15016 13812 15068 13821
rect 20352 13812 20404 13864
rect 2320 13676 2372 13728
rect 15752 13676 15804 13728
rect 22100 13812 22152 13864
rect 22652 13744 22704 13796
rect 22100 13676 22152 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 9588 13472 9640 13524
rect 15936 13472 15988 13524
rect 19432 13472 19484 13524
rect 2136 13404 2188 13456
rect 57152 13379 57204 13388
rect 57152 13345 57161 13379
rect 57161 13345 57195 13379
rect 57195 13345 57204 13379
rect 57152 13336 57204 13345
rect 57336 13379 57388 13388
rect 57336 13345 57354 13379
rect 57354 13345 57388 13379
rect 57336 13336 57388 13345
rect 58624 13404 58676 13456
rect 57704 13379 57756 13388
rect 57704 13345 57713 13379
rect 57713 13345 57747 13379
rect 57747 13345 57756 13379
rect 57704 13336 57756 13345
rect 58716 13336 58768 13388
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 58256 13268 58308 13320
rect 16948 13243 17000 13252
rect 16948 13209 16957 13243
rect 16957 13209 16991 13243
rect 16991 13209 17000 13243
rect 16948 13200 17000 13209
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 16028 13132 16080 13184
rect 55680 13132 55732 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 16948 12928 17000 12980
rect 1952 12792 2004 12844
rect 19432 12928 19484 12980
rect 57152 12928 57204 12980
rect 20076 12792 20128 12844
rect 57888 12792 57940 12844
rect 1860 12656 1912 12708
rect 10876 12656 10928 12708
rect 20628 12724 20680 12776
rect 57336 12656 57388 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4988 12384 5040 12436
rect 9220 12427 9272 12436
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 19432 12427 19484 12436
rect 19432 12393 19441 12427
rect 19441 12393 19475 12427
rect 19475 12393 19484 12427
rect 19432 12384 19484 12393
rect 57888 12384 57940 12436
rect 15844 12359 15896 12368
rect 15844 12325 15853 12359
rect 15853 12325 15887 12359
rect 15887 12325 15896 12359
rect 15844 12316 15896 12325
rect 9312 12248 9364 12300
rect 16672 12248 16724 12300
rect 58072 12248 58124 12300
rect 58624 12248 58676 12300
rect 55680 12223 55732 12232
rect 55680 12189 55689 12223
rect 55689 12189 55723 12223
rect 55723 12189 55732 12223
rect 55680 12180 55732 12189
rect 58348 12223 58400 12232
rect 58348 12189 58357 12223
rect 58357 12189 58391 12223
rect 58391 12189 58400 12223
rect 58348 12180 58400 12189
rect 9404 12112 9456 12164
rect 12624 12112 12676 12164
rect 13176 12112 13228 12164
rect 13728 12112 13780 12164
rect 16028 12112 16080 12164
rect 18696 12112 18748 12164
rect 42984 12044 43036 12096
rect 58072 12044 58124 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 5172 11840 5224 11892
rect 2504 11772 2556 11824
rect 6276 11772 6328 11824
rect 11336 11840 11388 11892
rect 13728 11772 13780 11824
rect 15844 11772 15896 11824
rect 19892 11772 19944 11824
rect 9312 11747 9364 11756
rect 1676 11611 1728 11620
rect 1676 11577 1685 11611
rect 1685 11577 1719 11611
rect 1719 11577 1728 11611
rect 1676 11568 1728 11577
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 19432 11704 19484 11756
rect 58348 11747 58400 11756
rect 58348 11713 58357 11747
rect 58357 11713 58391 11747
rect 58391 11713 58400 11747
rect 58348 11704 58400 11713
rect 9128 11636 9180 11688
rect 14464 11636 14516 11688
rect 15016 11636 15068 11688
rect 2688 11568 2740 11620
rect 57244 11568 57296 11620
rect 57428 11568 57480 11620
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 4804 11500 4856 11552
rect 6828 11500 6880 11552
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 20720 11543 20772 11552
rect 20720 11509 20729 11543
rect 20729 11509 20763 11543
rect 20763 11509 20772 11543
rect 20720 11500 20772 11509
rect 56692 11500 56744 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2412 11296 2464 11348
rect 12348 11296 12400 11348
rect 18512 11296 18564 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 57152 11296 57204 11348
rect 57428 11296 57480 11348
rect 58992 11296 59044 11348
rect 6736 11271 6788 11280
rect 2136 11203 2188 11212
rect 2136 11169 2145 11203
rect 2145 11169 2179 11203
rect 2179 11169 2188 11203
rect 2136 11160 2188 11169
rect 2504 11092 2556 11144
rect 6736 11237 6745 11271
rect 6745 11237 6779 11271
rect 6779 11237 6788 11271
rect 6736 11228 6788 11237
rect 5816 11160 5868 11212
rect 6828 11160 6880 11212
rect 16212 11160 16264 11212
rect 4620 11092 4672 11144
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 19984 11160 20036 11212
rect 21088 11160 21140 11212
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 5172 11024 5224 11076
rect 6000 11024 6052 11076
rect 20168 11092 20220 11144
rect 20628 11092 20680 11144
rect 20720 11092 20772 11144
rect 20812 11024 20864 11076
rect 56968 11160 57020 11212
rect 58164 11228 58216 11280
rect 57704 11203 57756 11212
rect 57704 11169 57713 11203
rect 57713 11169 57747 11203
rect 57747 11169 57756 11203
rect 57704 11160 57756 11169
rect 57428 11135 57480 11144
rect 57428 11101 57437 11135
rect 57437 11101 57471 11135
rect 57471 11101 57480 11135
rect 57428 11092 57480 11101
rect 57980 11092 58032 11144
rect 58348 11135 58400 11144
rect 58348 11101 58357 11135
rect 58357 11101 58391 11135
rect 58391 11101 58400 11135
rect 58348 11092 58400 11101
rect 22100 11024 22152 11076
rect 22560 11024 22612 11076
rect 13544 10956 13596 11008
rect 20720 10956 20772 11008
rect 20904 10999 20956 11008
rect 20904 10965 20913 10999
rect 20913 10965 20947 10999
rect 20947 10965 20956 10999
rect 20904 10956 20956 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 14464 10752 14516 10804
rect 5172 10684 5224 10736
rect 10600 10684 10652 10736
rect 13544 10684 13596 10736
rect 13820 10684 13872 10736
rect 16672 10752 16724 10804
rect 19432 10752 19484 10804
rect 56876 10795 56928 10804
rect 56876 10761 56885 10795
rect 56885 10761 56919 10795
rect 56919 10761 56928 10795
rect 56876 10752 56928 10761
rect 56968 10752 57020 10804
rect 57704 10752 57756 10804
rect 2136 10591 2188 10600
rect 2136 10557 2145 10591
rect 2145 10557 2179 10591
rect 2179 10557 2188 10591
rect 2136 10548 2188 10557
rect 2504 10548 2556 10600
rect 3056 10548 3108 10600
rect 5264 10548 5316 10600
rect 6000 10591 6052 10600
rect 6000 10557 6009 10591
rect 6009 10557 6043 10591
rect 6043 10557 6052 10591
rect 6000 10548 6052 10557
rect 18512 10616 18564 10668
rect 2688 10480 2740 10532
rect 2320 10412 2372 10464
rect 9680 10412 9732 10464
rect 12532 10455 12584 10464
rect 12532 10421 12541 10455
rect 12541 10421 12575 10455
rect 12575 10421 12584 10455
rect 19064 10548 19116 10600
rect 12532 10412 12584 10421
rect 18236 10412 18288 10464
rect 18420 10480 18472 10532
rect 20904 10616 20956 10668
rect 58440 10616 58492 10668
rect 57612 10412 57664 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 3332 10208 3384 10260
rect 3976 10208 4028 10260
rect 15108 10208 15160 10260
rect 18512 10251 18564 10260
rect 2044 10140 2096 10192
rect 18512 10217 18521 10251
rect 18521 10217 18555 10251
rect 18555 10217 18564 10251
rect 18512 10208 18564 10217
rect 19064 10208 19116 10260
rect 20628 10208 20680 10260
rect 58256 10208 58308 10260
rect 20168 10140 20220 10192
rect 58440 10140 58492 10192
rect 6000 10072 6052 10124
rect 6920 10072 6972 10124
rect 2412 10004 2464 10056
rect 9036 10072 9088 10124
rect 12532 10072 12584 10124
rect 16764 10115 16816 10124
rect 16764 10081 16773 10115
rect 16773 10081 16807 10115
rect 16807 10081 16816 10115
rect 16764 10072 16816 10081
rect 9312 10004 9364 10056
rect 12164 10004 12216 10056
rect 5172 9936 5224 9988
rect 6000 9936 6052 9988
rect 7288 9979 7340 9988
rect 7288 9945 7297 9979
rect 7297 9945 7331 9979
rect 7331 9945 7340 9979
rect 7288 9936 7340 9945
rect 2688 9868 2740 9920
rect 11060 9868 11112 9920
rect 12164 9911 12216 9920
rect 12164 9877 12173 9911
rect 12173 9877 12207 9911
rect 12207 9877 12216 9911
rect 58164 10047 58216 10056
rect 58164 10013 58173 10047
rect 58173 10013 58207 10047
rect 58207 10013 58216 10047
rect 58164 10004 58216 10013
rect 16028 9936 16080 9988
rect 17868 9936 17920 9988
rect 12164 9868 12216 9877
rect 14648 9868 14700 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 2688 9664 2740 9716
rect 9036 9664 9088 9716
rect 9312 9664 9364 9716
rect 56968 9707 57020 9716
rect 56968 9673 56977 9707
rect 56977 9673 57011 9707
rect 57011 9673 57020 9707
rect 56968 9664 57020 9673
rect 57704 9664 57756 9716
rect 5172 9596 5224 9648
rect 5816 9596 5868 9648
rect 6000 9596 6052 9648
rect 4068 9528 4120 9580
rect 13820 9596 13872 9648
rect 17776 9596 17828 9648
rect 20168 9596 20220 9648
rect 20812 9639 20864 9648
rect 20812 9605 20821 9639
rect 20821 9605 20855 9639
rect 20855 9605 20864 9639
rect 20812 9596 20864 9605
rect 2412 9503 2464 9512
rect 2412 9469 2421 9503
rect 2421 9469 2455 9503
rect 2455 9469 2464 9503
rect 2412 9460 2464 9469
rect 1676 9435 1728 9444
rect 1676 9401 1685 9435
rect 1685 9401 1719 9435
rect 1719 9401 1728 9435
rect 1676 9392 1728 9401
rect 2228 9392 2280 9444
rect 6920 9460 6972 9512
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 14464 9460 14516 9512
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 17868 9392 17920 9444
rect 58164 9571 58216 9580
rect 58164 9537 58173 9571
rect 58173 9537 58207 9571
rect 58207 9537 58216 9571
rect 58164 9528 58216 9537
rect 21088 9503 21140 9512
rect 21088 9469 21097 9503
rect 21097 9469 21131 9503
rect 21131 9469 21140 9503
rect 21088 9460 21140 9469
rect 58348 9435 58400 9444
rect 58348 9401 58357 9435
rect 58357 9401 58391 9435
rect 58391 9401 58400 9435
rect 58348 9392 58400 9401
rect 13544 9324 13596 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 2688 9120 2740 9172
rect 5172 9120 5224 9172
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 2504 9052 2556 9104
rect 8208 9052 8260 9104
rect 4068 8984 4120 9036
rect 12164 9120 12216 9172
rect 13176 9163 13228 9172
rect 13176 9129 13185 9163
rect 13185 9129 13219 9163
rect 13219 9129 13228 9163
rect 13176 9120 13228 9129
rect 14372 9163 14424 9172
rect 14372 9129 14381 9163
rect 14381 9129 14415 9163
rect 14415 9129 14424 9163
rect 14372 9120 14424 9129
rect 20168 9120 20220 9172
rect 57796 9120 57848 9172
rect 9312 8984 9364 9036
rect 20352 8984 20404 9036
rect 22744 8984 22796 9036
rect 56968 8984 57020 9036
rect 57336 9027 57388 9036
rect 57336 8993 57354 9027
rect 57354 8993 57388 9027
rect 57336 8984 57388 8993
rect 57704 9027 57756 9036
rect 57704 8993 57713 9027
rect 57713 8993 57747 9027
rect 57747 8993 57756 9027
rect 57704 8984 57756 8993
rect 2228 8916 2280 8968
rect 6368 8916 6420 8968
rect 12900 8916 12952 8968
rect 14372 8916 14424 8968
rect 20812 8916 20864 8968
rect 58348 8959 58400 8968
rect 10968 8848 11020 8900
rect 13176 8848 13228 8900
rect 22468 8848 22520 8900
rect 58348 8925 58357 8959
rect 58357 8925 58391 8959
rect 58391 8925 58400 8959
rect 58348 8916 58400 8925
rect 58900 8848 58952 8900
rect 20996 8823 21048 8832
rect 20996 8789 21005 8823
rect 21005 8789 21039 8823
rect 21039 8789 21048 8823
rect 20996 8780 21048 8789
rect 22192 8780 22244 8832
rect 22744 8823 22796 8832
rect 22744 8789 22753 8823
rect 22753 8789 22787 8823
rect 22787 8789 22796 8823
rect 22744 8780 22796 8789
rect 56508 8823 56560 8832
rect 56508 8789 56517 8823
rect 56517 8789 56551 8823
rect 56551 8789 56560 8823
rect 56508 8780 56560 8789
rect 56876 8780 56928 8832
rect 58256 8780 58308 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 3424 8576 3476 8628
rect 4068 8576 4120 8628
rect 6368 8576 6420 8628
rect 12900 8576 12952 8628
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 58072 8576 58124 8628
rect 58348 8619 58400 8628
rect 58348 8585 58357 8619
rect 58357 8585 58391 8619
rect 58391 8585 58400 8619
rect 58348 8576 58400 8585
rect 12808 8508 12860 8560
rect 56140 8508 56192 8560
rect 56876 8508 56928 8560
rect 22192 8483 22244 8492
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 22192 8449 22201 8483
rect 22201 8449 22235 8483
rect 22235 8449 22244 8483
rect 22192 8440 22244 8449
rect 56968 8483 57020 8492
rect 56968 8449 56977 8483
rect 56977 8449 57011 8483
rect 57011 8449 57020 8483
rect 56968 8440 57020 8449
rect 58532 8508 58584 8560
rect 58164 8483 58216 8492
rect 58164 8449 58173 8483
rect 58173 8449 58207 8483
rect 58207 8449 58216 8483
rect 58164 8440 58216 8449
rect 3424 8372 3476 8424
rect 57704 8372 57756 8424
rect 2136 8304 2188 8356
rect 2688 8304 2740 8356
rect 5908 8304 5960 8356
rect 53840 8304 53892 8356
rect 15660 8236 15712 8288
rect 20996 8236 21048 8288
rect 22008 8279 22060 8288
rect 22008 8245 22017 8279
rect 22017 8245 22051 8279
rect 22051 8245 22060 8279
rect 22008 8236 22060 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 2228 8032 2280 8084
rect 56968 8032 57020 8084
rect 57704 8075 57756 8084
rect 57704 8041 57713 8075
rect 57713 8041 57747 8075
rect 57747 8041 57756 8075
rect 57704 8032 57756 8041
rect 58256 8032 58308 8084
rect 2688 7964 2740 8016
rect 2504 7896 2556 7948
rect 5908 7939 5960 7948
rect 5908 7905 5917 7939
rect 5917 7905 5951 7939
rect 5951 7905 5960 7939
rect 5908 7896 5960 7905
rect 15660 7896 15712 7948
rect 22008 7896 22060 7948
rect 22560 7939 22612 7948
rect 22560 7905 22569 7939
rect 22569 7905 22603 7939
rect 22603 7905 22612 7939
rect 22560 7896 22612 7905
rect 2320 7828 2372 7880
rect 5356 7760 5408 7812
rect 6000 7760 6052 7812
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 22284 7871 22336 7880
rect 22284 7837 22293 7871
rect 22293 7837 22327 7871
rect 22327 7837 22336 7871
rect 22284 7828 22336 7837
rect 58348 7871 58400 7880
rect 13820 7760 13872 7812
rect 58348 7837 58357 7871
rect 58357 7837 58391 7871
rect 58391 7837 58400 7871
rect 58348 7828 58400 7837
rect 22836 7760 22888 7812
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 2688 7488 2740 7540
rect 2872 7488 2924 7540
rect 3976 7488 4028 7540
rect 9312 7488 9364 7540
rect 10876 7488 10928 7540
rect 9588 7395 9640 7404
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 9588 7352 9640 7361
rect 12808 7352 12860 7404
rect 2136 7327 2188 7336
rect 2136 7293 2145 7327
rect 2145 7293 2179 7327
rect 2179 7293 2188 7327
rect 2136 7284 2188 7293
rect 2504 7284 2556 7336
rect 13912 7420 13964 7472
rect 58348 7488 58400 7540
rect 22744 7420 22796 7472
rect 58164 7420 58216 7472
rect 16856 7352 16908 7404
rect 17868 7352 17920 7404
rect 19984 7352 20036 7404
rect 22284 7352 22336 7404
rect 22836 7395 22888 7404
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 18788 7284 18840 7336
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 56968 7191 57020 7200
rect 56968 7157 56977 7191
rect 56977 7157 57011 7191
rect 57011 7157 57020 7191
rect 56968 7148 57020 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3424 6944 3476 6996
rect 21088 6944 21140 6996
rect 57060 6944 57112 6996
rect 57704 6987 57756 6996
rect 57704 6953 57713 6987
rect 57713 6953 57747 6987
rect 57747 6953 57756 6987
rect 57704 6944 57756 6953
rect 2136 6808 2188 6860
rect 2872 6808 2924 6860
rect 20628 6851 20680 6860
rect 2504 6740 2556 6792
rect 20628 6817 20637 6851
rect 20637 6817 20671 6851
rect 20671 6817 20680 6851
rect 20628 6808 20680 6817
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 19432 6740 19484 6792
rect 22284 6808 22336 6860
rect 57704 6808 57756 6860
rect 5356 6672 5408 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 2780 6604 2832 6613
rect 3240 6604 3292 6656
rect 3516 6604 3568 6656
rect 9404 6672 9456 6724
rect 22192 6740 22244 6792
rect 22928 6783 22980 6792
rect 22928 6749 22937 6783
rect 22937 6749 22971 6783
rect 22971 6749 22980 6783
rect 22928 6740 22980 6749
rect 55404 6740 55456 6792
rect 56048 6740 56100 6792
rect 56876 6740 56928 6792
rect 56968 6740 57020 6792
rect 58348 6783 58400 6792
rect 58348 6749 58357 6783
rect 58357 6749 58391 6783
rect 58391 6749 58400 6783
rect 58348 6740 58400 6749
rect 22100 6672 22152 6724
rect 17776 6604 17828 6656
rect 22284 6604 22336 6656
rect 58164 6647 58216 6656
rect 58164 6613 58173 6647
rect 58173 6613 58207 6647
rect 58207 6613 58216 6647
rect 58164 6604 58216 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 2320 6400 2372 6452
rect 5356 6400 5408 6452
rect 9588 6375 9640 6384
rect 9588 6341 9597 6375
rect 9597 6341 9631 6375
rect 9631 6341 9640 6375
rect 9588 6332 9640 6341
rect 2228 6264 2280 6316
rect 2780 6264 2832 6316
rect 14740 6400 14792 6452
rect 19248 6443 19300 6452
rect 19248 6409 19257 6443
rect 19257 6409 19291 6443
rect 19291 6409 19300 6443
rect 19248 6400 19300 6409
rect 19432 6400 19484 6452
rect 13452 6375 13504 6384
rect 13452 6341 13461 6375
rect 13461 6341 13495 6375
rect 13495 6341 13504 6375
rect 13452 6332 13504 6341
rect 13912 6332 13964 6384
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 2872 6060 2924 6112
rect 13452 6196 13504 6248
rect 13544 6196 13596 6248
rect 19248 6264 19300 6316
rect 58164 6400 58216 6452
rect 56692 6307 56744 6316
rect 56692 6273 56726 6307
rect 56726 6273 56744 6307
rect 56876 6307 56928 6316
rect 56692 6264 56744 6273
rect 56876 6273 56885 6307
rect 56885 6273 56919 6307
rect 56919 6273 56928 6307
rect 56876 6264 56928 6273
rect 58348 6307 58400 6316
rect 58348 6273 58357 6307
rect 58357 6273 58391 6307
rect 58391 6273 58400 6307
rect 58348 6264 58400 6273
rect 14924 6239 14976 6248
rect 14924 6205 14933 6239
rect 14933 6205 14967 6239
rect 14967 6205 14976 6239
rect 14924 6196 14976 6205
rect 18696 6196 18748 6248
rect 20628 6196 20680 6248
rect 55864 6239 55916 6248
rect 55864 6205 55873 6239
rect 55873 6205 55907 6239
rect 55907 6205 55916 6239
rect 55864 6196 55916 6205
rect 58808 6196 58860 6248
rect 8576 6060 8628 6112
rect 9496 6060 9548 6112
rect 22192 6060 22244 6112
rect 57060 6060 57112 6112
rect 57244 6060 57296 6112
rect 58164 6103 58216 6112
rect 58164 6069 58173 6103
rect 58173 6069 58207 6103
rect 58207 6069 58216 6103
rect 58164 6060 58216 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1676 5899 1728 5908
rect 1676 5865 1685 5899
rect 1685 5865 1719 5899
rect 1719 5865 1728 5899
rect 1676 5856 1728 5865
rect 13084 5856 13136 5908
rect 18788 5899 18840 5908
rect 18788 5865 18797 5899
rect 18797 5865 18831 5899
rect 18831 5865 18840 5899
rect 18788 5856 18840 5865
rect 19984 5856 20036 5908
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 22100 5720 22152 5772
rect 58164 5856 58216 5908
rect 57060 5788 57112 5840
rect 57428 5763 57480 5772
rect 57428 5729 57437 5763
rect 57437 5729 57471 5763
rect 57471 5729 57480 5763
rect 57428 5720 57480 5729
rect 57612 5720 57664 5772
rect 2504 5652 2556 5704
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 20260 5652 20312 5704
rect 56692 5695 56744 5704
rect 56692 5661 56701 5695
rect 56701 5661 56735 5695
rect 56735 5661 56744 5695
rect 56692 5652 56744 5661
rect 57704 5695 57756 5704
rect 57704 5661 57713 5695
rect 57713 5661 57747 5695
rect 57747 5661 57756 5695
rect 57704 5652 57756 5661
rect 9404 5584 9456 5636
rect 57704 5516 57756 5568
rect 58256 5516 58308 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 12808 5312 12860 5364
rect 19432 5312 19484 5364
rect 20260 5312 20312 5364
rect 57060 5312 57112 5364
rect 57520 5355 57572 5364
rect 57520 5321 57529 5355
rect 57529 5321 57563 5355
rect 57563 5321 57572 5355
rect 57520 5312 57572 5321
rect 58716 5312 58768 5364
rect 9404 5244 9456 5296
rect 2412 5176 2464 5228
rect 10324 5151 10376 5160
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 1676 5083 1728 5092
rect 1676 5049 1685 5083
rect 1685 5049 1719 5083
rect 1719 5049 1728 5083
rect 1676 5040 1728 5049
rect 58348 5219 58400 5228
rect 58348 5185 58357 5219
rect 58357 5185 58391 5219
rect 58391 5185 58400 5219
rect 58348 5176 58400 5185
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 16856 5108 16908 5160
rect 20720 5040 20772 5092
rect 7656 4972 7708 5024
rect 8576 5015 8628 5024
rect 8576 4981 8585 5015
rect 8585 4981 8619 5015
rect 8619 4981 8628 5015
rect 8576 4972 8628 4981
rect 9496 4972 9548 5024
rect 10324 4972 10376 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 5448 4768 5500 4820
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 8576 4768 8628 4820
rect 18972 4700 19024 4752
rect 9496 4632 9548 4684
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 18144 4632 18196 4684
rect 18880 4675 18932 4684
rect 18880 4641 18889 4675
rect 18889 4641 18923 4675
rect 18923 4641 18932 4675
rect 18880 4632 18932 4641
rect 57796 4768 57848 4820
rect 57980 4768 58032 4820
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 22100 4564 22152 4616
rect 57520 4607 57572 4616
rect 57520 4573 57529 4607
rect 57529 4573 57563 4607
rect 57563 4573 57572 4607
rect 57520 4564 57572 4573
rect 58348 4607 58400 4616
rect 58348 4573 58357 4607
rect 58357 4573 58391 4607
rect 58391 4573 58400 4607
rect 58348 4564 58400 4573
rect 8300 4496 8352 4548
rect 9404 4496 9456 4548
rect 14740 4496 14792 4548
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 1676 4428 1728 4437
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 20076 4471 20128 4480
rect 20076 4437 20085 4471
rect 20085 4437 20119 4471
rect 20119 4437 20128 4471
rect 20076 4428 20128 4437
rect 22376 4428 22428 4480
rect 22652 4428 22704 4480
rect 56324 4428 56376 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 3240 4156 3292 4208
rect 4620 4156 4672 4208
rect 13912 4156 13964 4208
rect 14740 4156 14792 4208
rect 18972 4224 19024 4276
rect 9036 4088 9088 4140
rect 16856 4156 16908 4208
rect 2412 4020 2464 4072
rect 6368 4020 6420 4072
rect 11704 4020 11756 4072
rect 18880 4088 18932 4140
rect 20628 4088 20680 4140
rect 22192 4088 22244 4140
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 22744 4088 22796 4140
rect 55956 4088 56008 4140
rect 56600 4131 56652 4140
rect 56600 4097 56609 4131
rect 56609 4097 56643 4131
rect 56643 4097 56652 4131
rect 56600 4088 56652 4097
rect 57152 4088 57204 4140
rect 15936 4020 15988 4072
rect 18052 4020 18104 4072
rect 19800 4063 19852 4072
rect 19800 4029 19809 4063
rect 19809 4029 19843 4063
rect 19843 4029 19852 4063
rect 19800 4020 19852 4029
rect 56508 4020 56560 4072
rect 2780 3952 2832 4004
rect 9496 3952 9548 4004
rect 2228 3884 2280 3936
rect 3240 3927 3292 3936
rect 3240 3893 3249 3927
rect 3249 3893 3283 3927
rect 3283 3893 3292 3927
rect 3240 3884 3292 3893
rect 12256 3927 12308 3936
rect 12256 3893 12265 3927
rect 12265 3893 12299 3927
rect 12299 3893 12308 3927
rect 12256 3884 12308 3893
rect 50160 3952 50212 4004
rect 16672 3884 16724 3936
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 19340 3884 19392 3936
rect 20352 3884 20404 3936
rect 20720 3884 20772 3936
rect 57428 3884 57480 3936
rect 58072 3927 58124 3936
rect 58072 3893 58081 3927
rect 58081 3893 58115 3927
rect 58115 3893 58124 3927
rect 58072 3884 58124 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 10692 3680 10744 3732
rect 13360 3723 13412 3732
rect 1860 3612 1912 3664
rect 2780 3544 2832 3596
rect 3424 3544 3476 3596
rect 11612 3544 11664 3596
rect 13360 3689 13369 3723
rect 13369 3689 13403 3723
rect 13403 3689 13412 3723
rect 13360 3680 13412 3689
rect 18880 3723 18932 3732
rect 13268 3612 13320 3664
rect 18880 3689 18889 3723
rect 18889 3689 18923 3723
rect 18923 3689 18932 3723
rect 18880 3680 18932 3689
rect 22744 3723 22796 3732
rect 22744 3689 22753 3723
rect 22753 3689 22787 3723
rect 22787 3689 22796 3723
rect 22744 3680 22796 3689
rect 20352 3612 20404 3664
rect 20720 3612 20772 3664
rect 21364 3612 21416 3664
rect 15660 3544 15712 3596
rect 16856 3544 16908 3596
rect 19800 3544 19852 3596
rect 22100 3587 22152 3596
rect 2964 3408 3016 3460
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 5172 3408 5224 3460
rect 8300 3476 8352 3528
rect 14740 3476 14792 3528
rect 6368 3408 6420 3460
rect 8024 3408 8076 3460
rect 7288 3383 7340 3392
rect 7288 3349 7297 3383
rect 7297 3349 7331 3383
rect 7331 3349 7340 3383
rect 7288 3340 7340 3349
rect 8944 3340 8996 3392
rect 12164 3408 12216 3460
rect 15844 3340 15896 3392
rect 15936 3340 15988 3392
rect 20260 3408 20312 3460
rect 20812 3476 20864 3528
rect 22100 3553 22109 3587
rect 22109 3553 22143 3587
rect 22143 3553 22152 3587
rect 22100 3544 22152 3553
rect 22468 3476 22520 3528
rect 22560 3476 22612 3528
rect 53840 3612 53892 3664
rect 44824 3544 44876 3596
rect 58624 3544 58676 3596
rect 48504 3519 48556 3528
rect 21088 3408 21140 3460
rect 48504 3485 48513 3519
rect 48513 3485 48547 3519
rect 48547 3485 48556 3519
rect 48504 3476 48556 3485
rect 53104 3519 53156 3528
rect 53104 3485 53113 3519
rect 53113 3485 53147 3519
rect 53147 3485 53156 3519
rect 53104 3476 53156 3485
rect 54668 3476 54720 3528
rect 55956 3476 56008 3528
rect 56600 3476 56652 3528
rect 57244 3476 57296 3528
rect 57612 3519 57664 3528
rect 57612 3485 57621 3519
rect 57621 3485 57655 3519
rect 57655 3485 57664 3519
rect 57612 3476 57664 3485
rect 55588 3408 55640 3460
rect 20720 3340 20772 3392
rect 22100 3340 22152 3392
rect 38936 3383 38988 3392
rect 38936 3349 38945 3383
rect 38945 3349 38979 3383
rect 38979 3349 38988 3383
rect 38936 3340 38988 3349
rect 45744 3340 45796 3392
rect 48320 3383 48372 3392
rect 48320 3349 48329 3383
rect 48329 3349 48363 3383
rect 48363 3349 48372 3383
rect 48320 3340 48372 3349
rect 52920 3383 52972 3392
rect 52920 3349 52929 3383
rect 52929 3349 52963 3383
rect 52963 3349 52972 3383
rect 52920 3340 52972 3349
rect 54392 3383 54444 3392
rect 54392 3349 54401 3383
rect 54401 3349 54435 3383
rect 54435 3349 54444 3383
rect 54392 3340 54444 3349
rect 55496 3383 55548 3392
rect 55496 3349 55505 3383
rect 55505 3349 55539 3383
rect 55539 3349 55548 3383
rect 55496 3340 55548 3349
rect 55772 3340 55824 3392
rect 56968 3383 57020 3392
rect 56968 3349 56977 3383
rect 56977 3349 57011 3383
rect 57011 3349 57020 3383
rect 56968 3340 57020 3349
rect 57796 3383 57848 3392
rect 57796 3349 57805 3383
rect 57805 3349 57839 3383
rect 57839 3349 57848 3383
rect 57796 3340 57848 3349
rect 58348 3383 58400 3392
rect 58348 3349 58357 3383
rect 58357 3349 58391 3383
rect 58391 3349 58400 3383
rect 58348 3340 58400 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 2412 3136 2464 3188
rect 2780 3068 2832 3120
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 4896 3136 4948 3188
rect 5172 3136 5224 3188
rect 6368 3136 6420 3188
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 11704 3179 11756 3188
rect 11704 3145 11713 3179
rect 11713 3145 11747 3179
rect 11747 3145 11756 3179
rect 11704 3136 11756 3145
rect 9496 3111 9548 3120
rect 9496 3077 9505 3111
rect 9505 3077 9539 3111
rect 9539 3077 9548 3111
rect 9496 3068 9548 3077
rect 12164 3068 12216 3120
rect 2964 3000 3016 3009
rect 5908 3000 5960 3052
rect 8392 3000 8444 3052
rect 10324 3000 10376 3052
rect 14740 3068 14792 3120
rect 22560 3179 22612 3188
rect 22560 3145 22569 3179
rect 22569 3145 22603 3179
rect 22603 3145 22612 3179
rect 22560 3136 22612 3145
rect 23940 3136 23992 3188
rect 28724 3179 28776 3188
rect 15844 3068 15896 3120
rect 21364 3111 21416 3120
rect 21364 3077 21373 3111
rect 21373 3077 21407 3111
rect 21407 3077 21416 3111
rect 21364 3068 21416 3077
rect 13912 3000 13964 3052
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 18052 3000 18104 3052
rect 18972 3000 19024 3052
rect 19340 3043 19392 3052
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 20444 3000 20496 3052
rect 20628 3000 20680 3052
rect 22376 3043 22428 3052
rect 22376 3009 22385 3043
rect 22385 3009 22419 3043
rect 22419 3009 22428 3043
rect 22376 3000 22428 3009
rect 28724 3145 28733 3179
rect 28733 3145 28767 3179
rect 28767 3145 28776 3179
rect 28724 3136 28776 3145
rect 29828 3179 29880 3188
rect 29828 3145 29837 3179
rect 29837 3145 29871 3179
rect 29871 3145 29880 3179
rect 29828 3136 29880 3145
rect 30932 3179 30984 3188
rect 30932 3145 30941 3179
rect 30941 3145 30975 3179
rect 30975 3145 30984 3179
rect 30932 3136 30984 3145
rect 33140 3179 33192 3188
rect 33140 3145 33149 3179
rect 33149 3145 33183 3179
rect 33183 3145 33192 3179
rect 33140 3136 33192 3145
rect 42984 3179 43036 3188
rect 42984 3145 42993 3179
rect 42993 3145 43027 3179
rect 43027 3145 43036 3179
rect 42984 3136 43036 3145
rect 43720 3179 43772 3188
rect 43720 3145 43729 3179
rect 43729 3145 43763 3179
rect 43763 3145 43772 3179
rect 43720 3136 43772 3145
rect 44824 3179 44876 3188
rect 44824 3145 44833 3179
rect 44833 3145 44867 3179
rect 44867 3145 44876 3179
rect 44824 3136 44876 3145
rect 51448 3179 51500 3188
rect 51448 3145 51457 3179
rect 51457 3145 51491 3179
rect 51491 3145 51500 3179
rect 51448 3136 51500 3145
rect 54668 3179 54720 3188
rect 54668 3145 54677 3179
rect 54677 3145 54711 3179
rect 54711 3145 54720 3179
rect 54668 3136 54720 3145
rect 55864 3179 55916 3188
rect 55864 3145 55873 3179
rect 55873 3145 55907 3179
rect 55907 3145 55916 3179
rect 55864 3136 55916 3145
rect 56692 3136 56744 3188
rect 30288 3068 30340 3120
rect 32312 3111 32364 3120
rect 32312 3077 32321 3111
rect 32321 3077 32355 3111
rect 32355 3077 32364 3111
rect 32312 3068 32364 3077
rect 37740 3068 37792 3120
rect 1952 2796 2004 2848
rect 17776 2932 17828 2984
rect 40316 2932 40368 2984
rect 50160 2932 50212 2984
rect 50620 2932 50672 2984
rect 54484 2932 54536 2984
rect 56048 3043 56100 3052
rect 56048 3009 56057 3043
rect 56057 3009 56091 3043
rect 56091 3009 56100 3043
rect 56048 3000 56100 3009
rect 58348 3068 58400 3120
rect 57336 3043 57388 3052
rect 57336 3009 57345 3043
rect 57345 3009 57379 3043
rect 57379 3009 57388 3043
rect 57336 3000 57388 3009
rect 58256 3043 58308 3052
rect 58256 3009 58265 3043
rect 58265 3009 58299 3043
rect 58299 3009 58308 3043
rect 58256 3000 58308 3009
rect 38660 2907 38712 2916
rect 38660 2873 38669 2907
rect 38669 2873 38703 2907
rect 38703 2873 38712 2907
rect 38660 2864 38712 2873
rect 56968 2864 57020 2916
rect 7840 2796 7892 2848
rect 10048 2796 10100 2848
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 13820 2796 13872 2848
rect 18880 2796 18932 2848
rect 23296 2796 23348 2848
rect 24400 2839 24452 2848
rect 24400 2805 24409 2839
rect 24409 2805 24443 2839
rect 24443 2805 24452 2839
rect 24400 2796 24452 2805
rect 25504 2839 25556 2848
rect 25504 2805 25513 2839
rect 25513 2805 25547 2839
rect 25547 2805 25556 2839
rect 25504 2796 25556 2805
rect 27712 2796 27764 2848
rect 35992 2839 36044 2848
rect 35992 2805 36001 2839
rect 36001 2805 36035 2839
rect 36035 2805 36044 2839
rect 35992 2796 36044 2805
rect 55956 2796 56008 2848
rect 57152 2839 57204 2848
rect 57152 2805 57161 2839
rect 57161 2805 57195 2839
rect 57195 2805 57204 2839
rect 57152 2796 57204 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4620 2592 4672 2644
rect 4804 2635 4856 2644
rect 4804 2601 4813 2635
rect 4813 2601 4847 2635
rect 4847 2601 4856 2635
rect 4804 2592 4856 2601
rect 14648 2635 14700 2644
rect 14648 2601 14657 2635
rect 14657 2601 14691 2635
rect 14691 2601 14700 2635
rect 14648 2592 14700 2601
rect 18696 2592 18748 2644
rect 22468 2635 22520 2644
rect 22468 2601 22477 2635
rect 22477 2601 22511 2635
rect 22511 2601 22520 2635
rect 22468 2592 22520 2601
rect 28908 2592 28960 2644
rect 4896 2524 4948 2576
rect 18236 2524 18288 2576
rect 39672 2524 39724 2576
rect 3976 2456 4028 2508
rect 2320 2388 2372 2440
rect 4528 2388 4580 2440
rect 18880 2499 18932 2508
rect 18880 2465 18889 2499
rect 18889 2465 18923 2499
rect 18923 2465 18932 2499
rect 18880 2456 18932 2465
rect 21088 2456 21140 2508
rect 22652 2456 22704 2508
rect 29736 2456 29788 2508
rect 55404 2592 55456 2644
rect 57612 2592 57664 2644
rect 56140 2524 56192 2576
rect 5632 2388 5684 2440
rect 6920 2388 6972 2440
rect 7288 2388 7340 2440
rect 12164 2388 12216 2440
rect 12440 2388 12492 2440
rect 13360 2388 13412 2440
rect 13820 2388 13872 2440
rect 14464 2388 14516 2440
rect 15568 2388 15620 2440
rect 19432 2388 19484 2440
rect 20996 2388 21048 2440
rect 4068 2252 4120 2304
rect 7840 2320 7892 2372
rect 8944 2320 8996 2372
rect 10048 2320 10100 2372
rect 11152 2320 11204 2372
rect 5908 2295 5960 2304
rect 5908 2261 5917 2295
rect 5917 2261 5951 2295
rect 5951 2261 5960 2295
rect 5908 2252 5960 2261
rect 8116 2295 8168 2304
rect 8116 2261 8125 2295
rect 8125 2261 8159 2295
rect 8159 2261 8168 2295
rect 8116 2252 8168 2261
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 16672 2320 16724 2372
rect 22192 2320 22244 2372
rect 23296 2388 23348 2440
rect 25504 2388 25556 2440
rect 28724 2388 28776 2440
rect 29828 2388 29880 2440
rect 30932 2388 30984 2440
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 33140 2388 33192 2440
rect 24400 2320 24452 2372
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 26608 2295 26660 2304
rect 26608 2261 26617 2295
rect 26617 2261 26651 2295
rect 26651 2261 26660 2295
rect 35992 2388 36044 2440
rect 37740 2431 37792 2440
rect 37740 2397 37749 2431
rect 37749 2397 37783 2431
rect 37783 2397 37792 2431
rect 37740 2388 37792 2397
rect 38660 2388 38712 2440
rect 38936 2431 38988 2440
rect 38936 2397 38945 2431
rect 38945 2397 38979 2431
rect 38979 2397 38988 2431
rect 38936 2388 38988 2397
rect 40316 2431 40368 2440
rect 40316 2397 40325 2431
rect 40325 2397 40359 2431
rect 40359 2397 40368 2431
rect 40316 2388 40368 2397
rect 42984 2388 43036 2440
rect 43720 2388 43772 2440
rect 44824 2388 44876 2440
rect 45744 2431 45796 2440
rect 45744 2397 45753 2431
rect 45753 2397 45787 2431
rect 45787 2397 45796 2431
rect 45744 2388 45796 2397
rect 57152 2456 57204 2508
rect 48320 2388 48372 2440
rect 49056 2431 49108 2440
rect 49056 2397 49065 2431
rect 49065 2397 49099 2431
rect 49099 2397 49108 2431
rect 49056 2388 49108 2397
rect 50620 2431 50672 2440
rect 50620 2397 50629 2431
rect 50629 2397 50663 2431
rect 50663 2397 50672 2431
rect 50620 2388 50672 2397
rect 51448 2388 51500 2440
rect 52920 2388 52972 2440
rect 54392 2388 54444 2440
rect 55496 2388 55548 2440
rect 55772 2431 55824 2440
rect 55772 2397 55781 2431
rect 55781 2397 55815 2431
rect 55815 2397 55824 2431
rect 55772 2388 55824 2397
rect 55956 2388 56008 2440
rect 56416 2388 56468 2440
rect 56232 2320 56284 2372
rect 56324 2320 56376 2372
rect 57796 2388 57848 2440
rect 26608 2252 26660 2261
rect 28816 2252 28868 2304
rect 29920 2252 29972 2304
rect 31024 2252 31076 2304
rect 32128 2252 32180 2304
rect 33232 2252 33284 2304
rect 34336 2295 34388 2304
rect 34336 2261 34345 2295
rect 34345 2261 34379 2295
rect 34379 2261 34388 2295
rect 34336 2252 34388 2261
rect 36544 2252 36596 2304
rect 37648 2252 37700 2304
rect 38752 2252 38804 2304
rect 39856 2252 39908 2304
rect 40960 2252 41012 2304
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 42064 2252 42116 2304
rect 43168 2252 43220 2304
rect 44272 2252 44324 2304
rect 45376 2252 45428 2304
rect 46480 2252 46532 2304
rect 47584 2252 47636 2304
rect 48688 2252 48740 2304
rect 49792 2252 49844 2304
rect 50896 2252 50948 2304
rect 52000 2252 52052 2304
rect 53104 2252 53156 2304
rect 54208 2252 54260 2304
rect 55312 2252 55364 2304
rect 57520 2252 57572 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 4804 2048 4856 2100
rect 22376 2048 22428 2100
rect 41880 2048 41932 2100
rect 58072 2048 58124 2100
rect 3240 1980 3292 2032
rect 8116 1980 8168 2032
rect 5908 1912 5960 1964
rect 20628 1912 20680 1964
rect 3332 1844 3384 1896
rect 12164 1844 12216 1896
rect 6184 1776 6236 1828
rect 13636 1776 13688 1828
rect 3516 1708 3568 1760
rect 10968 1708 11020 1760
<< metal2 >>
rect 1858 59200 1914 60000
rect 3054 59200 3110 60000
rect 4250 59200 4306 60000
rect 5446 59200 5502 60000
rect 6642 59200 6698 60000
rect 7838 59200 7894 60000
rect 9034 59200 9090 60000
rect 10230 59200 10286 60000
rect 11426 59200 11482 60000
rect 12622 59200 12678 60000
rect 13818 59200 13874 60000
rect 15014 59200 15070 60000
rect 16210 59200 16266 60000
rect 17406 59200 17462 60000
rect 18602 59200 18658 60000
rect 19798 59200 19854 60000
rect 20994 59200 21050 60000
rect 22190 59200 22246 60000
rect 23386 59200 23442 60000
rect 24582 59200 24638 60000
rect 25778 59200 25834 60000
rect 26974 59200 27030 60000
rect 28170 59200 28226 60000
rect 29366 59200 29422 60000
rect 30562 59200 30618 60000
rect 31758 59200 31814 60000
rect 32954 59200 33010 60000
rect 34150 59200 34206 60000
rect 35346 59200 35402 60000
rect 36542 59200 36598 60000
rect 37738 59200 37794 60000
rect 38934 59200 38990 60000
rect 40130 59200 40186 60000
rect 41326 59200 41382 60000
rect 42522 59200 42578 60000
rect 43718 59200 43774 60000
rect 44914 59200 44970 60000
rect 46110 59200 46166 60000
rect 47306 59200 47362 60000
rect 48502 59200 48558 60000
rect 49698 59200 49754 60000
rect 50894 59200 50950 60000
rect 52090 59200 52146 60000
rect 53286 59200 53342 60000
rect 54482 59200 54538 60000
rect 55678 59200 55734 60000
rect 56874 59200 56930 60000
rect 58070 59200 58126 60000
rect 1872 57458 1900 59200
rect 3068 57458 3096 59200
rect 4264 57458 4292 59200
rect 1860 57452 1912 57458
rect 1860 57394 1912 57400
rect 3056 57452 3108 57458
rect 3056 57394 3108 57400
rect 4252 57452 4304 57458
rect 4252 57394 4304 57400
rect 4620 57452 4672 57458
rect 5460 57440 5488 59200
rect 5540 57452 5592 57458
rect 5460 57412 5540 57440
rect 4620 57394 4672 57400
rect 5540 57394 5592 57400
rect 1872 57050 1900 57394
rect 3068 57050 3096 57394
rect 3148 57384 3200 57390
rect 3148 57326 3200 57332
rect 1860 57044 1912 57050
rect 1860 56986 1912 56992
rect 3056 57044 3108 57050
rect 3056 56986 3108 56992
rect 3160 55729 3188 57326
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4632 57050 4660 57394
rect 5724 57384 5776 57390
rect 5724 57326 5776 57332
rect 5448 57248 5500 57254
rect 5448 57190 5500 57196
rect 4620 57044 4672 57050
rect 4620 56986 4672 56992
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 1674 55720 1730 55729
rect 1674 55655 1730 55664
rect 3146 55720 3202 55729
rect 3146 55655 3202 55664
rect 1688 55622 1716 55655
rect 1676 55616 1728 55622
rect 1676 55558 1728 55564
rect 2320 55616 2372 55622
rect 2320 55558 2372 55564
rect 1676 55072 1728 55078
rect 1676 55014 1728 55020
rect 1688 54913 1716 55014
rect 1674 54904 1730 54913
rect 1674 54839 1730 54848
rect 1674 54088 1730 54097
rect 1674 54023 1676 54032
rect 1728 54023 1730 54032
rect 1676 53994 1728 54000
rect 1676 53440 1728 53446
rect 1676 53382 1728 53388
rect 1688 53281 1716 53382
rect 1674 53272 1730 53281
rect 1674 53207 1730 53216
rect 1676 52624 1728 52630
rect 1676 52566 1728 52572
rect 1688 52465 1716 52566
rect 1674 52456 1730 52465
rect 1674 52391 1730 52400
rect 1676 51808 1728 51814
rect 1676 51750 1728 51756
rect 1688 51649 1716 51750
rect 1674 51640 1730 51649
rect 1674 51575 1730 51584
rect 1674 50824 1730 50833
rect 1674 50759 1676 50768
rect 1728 50759 1730 50768
rect 1676 50730 1728 50736
rect 1952 50312 2004 50318
rect 1952 50254 2004 50260
rect 1676 50176 1728 50182
rect 1676 50118 1728 50124
rect 1688 50017 1716 50118
rect 1674 50008 1730 50017
rect 1674 49943 1730 49952
rect 1674 49192 1730 49201
rect 1674 49127 1730 49136
rect 1688 49094 1716 49127
rect 1676 49088 1728 49094
rect 1676 49030 1728 49036
rect 1676 48544 1728 48550
rect 1676 48486 1728 48492
rect 1688 48385 1716 48486
rect 1674 48376 1730 48385
rect 1674 48311 1730 48320
rect 1674 47560 1730 47569
rect 1674 47495 1676 47504
rect 1728 47495 1730 47504
rect 1676 47466 1728 47472
rect 1676 46912 1728 46918
rect 1676 46854 1728 46860
rect 1688 46753 1716 46854
rect 1674 46744 1730 46753
rect 1674 46679 1730 46688
rect 1674 45928 1730 45937
rect 1674 45863 1730 45872
rect 1688 45830 1716 45863
rect 1676 45824 1728 45830
rect 1676 45766 1728 45772
rect 1676 45280 1728 45286
rect 1676 45222 1728 45228
rect 1688 45121 1716 45222
rect 1674 45112 1730 45121
rect 1674 45047 1730 45056
rect 1674 44296 1730 44305
rect 1674 44231 1676 44240
rect 1728 44231 1730 44240
rect 1676 44202 1728 44208
rect 1676 43648 1728 43654
rect 1676 43590 1728 43596
rect 1688 43489 1716 43590
rect 1674 43480 1730 43489
rect 1674 43415 1730 43424
rect 1674 42664 1730 42673
rect 1674 42599 1730 42608
rect 1688 42566 1716 42599
rect 1676 42560 1728 42566
rect 1676 42502 1728 42508
rect 1676 42016 1728 42022
rect 1676 41958 1728 41964
rect 1688 41857 1716 41958
rect 1674 41848 1730 41857
rect 1674 41783 1730 41792
rect 1674 41032 1730 41041
rect 1674 40967 1676 40976
rect 1728 40967 1730 40976
rect 1676 40938 1728 40944
rect 1676 40384 1728 40390
rect 1676 40326 1728 40332
rect 1688 40225 1716 40326
rect 1674 40216 1730 40225
rect 1674 40151 1730 40160
rect 1674 39400 1730 39409
rect 1674 39335 1730 39344
rect 1688 39302 1716 39335
rect 1676 39296 1728 39302
rect 1676 39238 1728 39244
rect 1676 38752 1728 38758
rect 1676 38694 1728 38700
rect 1688 38593 1716 38694
rect 1674 38584 1730 38593
rect 1674 38519 1730 38528
rect 1674 37768 1730 37777
rect 1674 37703 1676 37712
rect 1728 37703 1730 37712
rect 1676 37674 1728 37680
rect 1676 37120 1728 37126
rect 1676 37062 1728 37068
rect 1688 36961 1716 37062
rect 1674 36952 1730 36961
rect 1674 36887 1730 36896
rect 1674 36136 1730 36145
rect 1674 36071 1730 36080
rect 1688 36038 1716 36071
rect 1676 36032 1728 36038
rect 1676 35974 1728 35980
rect 1676 35488 1728 35494
rect 1676 35430 1728 35436
rect 1688 35329 1716 35430
rect 1674 35320 1730 35329
rect 1674 35255 1730 35264
rect 1674 34504 1730 34513
rect 1674 34439 1676 34448
rect 1728 34439 1730 34448
rect 1676 34410 1728 34416
rect 1676 33856 1728 33862
rect 1676 33798 1728 33804
rect 1688 33697 1716 33798
rect 1674 33688 1730 33697
rect 1674 33623 1730 33632
rect 1674 32872 1730 32881
rect 1674 32807 1730 32816
rect 1688 32774 1716 32807
rect 1676 32768 1728 32774
rect 1676 32710 1728 32716
rect 1676 32224 1728 32230
rect 1676 32166 1728 32172
rect 1688 32065 1716 32166
rect 1674 32056 1730 32065
rect 1674 31991 1730 32000
rect 1964 31634 1992 50254
rect 2044 48748 2096 48754
rect 2044 48690 2096 48696
rect 2056 48550 2084 48690
rect 2044 48544 2096 48550
rect 2044 48486 2096 48492
rect 2056 31770 2084 48486
rect 2136 46980 2188 46986
rect 2136 46922 2188 46928
rect 2148 35894 2176 46922
rect 2332 45554 2360 55558
rect 2412 55276 2464 55282
rect 2412 55218 2464 55224
rect 2424 53106 2452 55218
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 2872 53984 2924 53990
rect 2872 53926 2924 53932
rect 2504 53440 2556 53446
rect 2504 53382 2556 53388
rect 2412 53100 2464 53106
rect 2412 53042 2464 53048
rect 2516 51066 2544 53382
rect 2780 52488 2832 52494
rect 2780 52430 2832 52436
rect 2504 51060 2556 51066
rect 2504 51002 2556 51008
rect 2596 50720 2648 50726
rect 2596 50662 2648 50668
rect 2332 45526 2452 45554
rect 2424 44878 2452 45526
rect 2412 44872 2464 44878
rect 2412 44814 2464 44820
rect 2412 37664 2464 37670
rect 2412 37606 2464 37612
rect 2424 37466 2452 37606
rect 2412 37460 2464 37466
rect 2412 37402 2464 37408
rect 2412 37120 2464 37126
rect 2412 37062 2464 37068
rect 2424 36922 2452 37062
rect 2412 36916 2464 36922
rect 2412 36858 2464 36864
rect 2148 35866 2360 35894
rect 2056 31742 2176 31770
rect 1964 31606 2084 31634
rect 1674 31240 1730 31249
rect 1674 31175 1676 31184
rect 1728 31175 1730 31184
rect 1676 31146 1728 31152
rect 1676 30592 1728 30598
rect 1676 30534 1728 30540
rect 1688 30433 1716 30534
rect 1674 30424 1730 30433
rect 1674 30359 1730 30368
rect 1674 29608 1730 29617
rect 1674 29543 1730 29552
rect 1688 29510 1716 29543
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1676 29028 1728 29034
rect 1676 28970 1728 28976
rect 1688 28801 1716 28970
rect 1674 28792 1730 28801
rect 1674 28727 1730 28736
rect 1952 28416 2004 28422
rect 1952 28358 2004 28364
rect 1674 27976 1730 27985
rect 1674 27911 1676 27920
rect 1728 27911 1730 27920
rect 1676 27882 1728 27888
rect 1964 27470 1992 28358
rect 2056 27470 2084 31606
rect 1952 27464 2004 27470
rect 1952 27406 2004 27412
rect 2044 27464 2096 27470
rect 2044 27406 2096 27412
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1688 27169 1716 27270
rect 1674 27160 1730 27169
rect 1674 27095 1730 27104
rect 1674 26344 1730 26353
rect 1674 26279 1730 26288
rect 1688 26042 1716 26279
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 1674 25528 1730 25537
rect 1674 25463 1676 25472
rect 1728 25463 1730 25472
rect 1676 25434 1728 25440
rect 1674 24712 1730 24721
rect 1674 24647 1676 24656
rect 1728 24647 1730 24656
rect 1860 24676 1912 24682
rect 1676 24618 1728 24624
rect 1860 24618 1912 24624
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1688 23905 1716 24006
rect 1674 23896 1730 23905
rect 1674 23831 1730 23840
rect 1674 23080 1730 23089
rect 1674 23015 1730 23024
rect 1688 22982 1716 23015
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1674 22264 1730 22273
rect 1674 22199 1676 22208
rect 1728 22199 1730 22208
rect 1676 22170 1728 22176
rect 1674 21448 1730 21457
rect 1674 21383 1730 21392
rect 1688 21146 1716 21383
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 1674 20632 1730 20641
rect 1674 20567 1676 20576
rect 1728 20567 1730 20576
rect 1676 20538 1728 20544
rect 1674 19816 1730 19825
rect 1674 19751 1730 19760
rect 1688 19514 1716 19751
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1872 19378 1900 24618
rect 1964 21418 1992 27406
rect 2148 26586 2176 31742
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 2240 31142 2268 31282
rect 2228 31136 2280 31142
rect 2228 31078 2280 31084
rect 2136 26580 2188 26586
rect 2136 26522 2188 26528
rect 2136 26036 2188 26042
rect 2136 25978 2188 25984
rect 2044 25900 2096 25906
rect 2044 25842 2096 25848
rect 2056 25226 2084 25842
rect 2044 25220 2096 25226
rect 2044 25162 2096 25168
rect 2044 23792 2096 23798
rect 2044 23734 2096 23740
rect 1952 21412 2004 21418
rect 1952 21354 2004 21360
rect 2056 20942 2084 23734
rect 2148 22574 2176 25978
rect 2136 22568 2188 22574
rect 2136 22510 2188 22516
rect 2148 22098 2176 22510
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 2240 21570 2268 31078
rect 2332 27130 2360 35866
rect 2504 33992 2556 33998
rect 2504 33934 2556 33940
rect 2412 30592 2464 30598
rect 2412 30534 2464 30540
rect 2320 27124 2372 27130
rect 2320 27066 2372 27072
rect 2320 26988 2372 26994
rect 2320 26930 2372 26936
rect 2332 26450 2360 26930
rect 2320 26444 2372 26450
rect 2320 26386 2372 26392
rect 2332 26042 2360 26386
rect 2320 26036 2372 26042
rect 2320 25978 2372 25984
rect 2424 25378 2452 30534
rect 2516 26450 2544 33934
rect 2504 26444 2556 26450
rect 2504 26386 2556 26392
rect 2608 25430 2636 50662
rect 2792 50386 2820 52430
rect 2780 50380 2832 50386
rect 2780 50322 2832 50328
rect 2884 47598 2912 53926
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 5460 53446 5488 57190
rect 5736 53990 5764 57326
rect 6656 56914 6684 59200
rect 7852 57458 7880 59200
rect 9048 57458 9076 59200
rect 10244 57458 10272 59200
rect 11440 57594 11468 59200
rect 11428 57588 11480 57594
rect 11428 57530 11480 57536
rect 11440 57458 11468 57530
rect 12636 57458 12664 59200
rect 13832 57594 13860 59200
rect 13820 57588 13872 57594
rect 13820 57530 13872 57536
rect 13832 57458 13860 57530
rect 15028 57458 15056 59200
rect 16224 57594 16252 59200
rect 16212 57588 16264 57594
rect 16212 57530 16264 57536
rect 16224 57458 16252 57530
rect 17420 57458 17448 59200
rect 18616 57458 18644 59200
rect 19812 57882 19840 59200
rect 19812 57854 20024 57882
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 19996 57458 20024 57854
rect 20720 57588 20772 57594
rect 20720 57530 20772 57536
rect 7840 57452 7892 57458
rect 7840 57394 7892 57400
rect 8484 57452 8536 57458
rect 8484 57394 8536 57400
rect 9036 57452 9088 57458
rect 9036 57394 9088 57400
rect 10232 57452 10284 57458
rect 10232 57394 10284 57400
rect 11428 57452 11480 57458
rect 11428 57394 11480 57400
rect 12624 57452 12676 57458
rect 12624 57394 12676 57400
rect 13820 57452 13872 57458
rect 13820 57394 13872 57400
rect 15016 57452 15068 57458
rect 15016 57394 15068 57400
rect 16212 57452 16264 57458
rect 16212 57394 16264 57400
rect 17408 57452 17460 57458
rect 17408 57394 17460 57400
rect 18604 57452 18656 57458
rect 18604 57394 18656 57400
rect 19984 57452 20036 57458
rect 19984 57394 20036 57400
rect 8300 57384 8352 57390
rect 8300 57326 8352 57332
rect 6644 56908 6696 56914
rect 6644 56850 6696 56856
rect 7012 56840 7064 56846
rect 7012 56782 7064 56788
rect 7024 55350 7052 56782
rect 8312 55826 8340 57326
rect 8496 57050 8524 57394
rect 9048 57050 9076 57394
rect 9312 57248 9364 57254
rect 9312 57190 9364 57196
rect 10508 57248 10560 57254
rect 10508 57190 10560 57196
rect 11888 57248 11940 57254
rect 11888 57190 11940 57196
rect 8484 57044 8536 57050
rect 8484 56986 8536 56992
rect 9036 57044 9088 57050
rect 9036 56986 9088 56992
rect 9324 56982 9352 57190
rect 9312 56976 9364 56982
rect 9312 56918 9364 56924
rect 10520 56914 10548 57190
rect 10508 56908 10560 56914
rect 10508 56850 10560 56856
rect 11900 56846 11928 57190
rect 12636 57050 12664 57394
rect 12900 57248 12952 57254
rect 12900 57190 12952 57196
rect 14464 57248 14516 57254
rect 14464 57190 14516 57196
rect 12624 57044 12676 57050
rect 12624 56986 12676 56992
rect 11888 56840 11940 56846
rect 11888 56782 11940 56788
rect 12912 56778 12940 57190
rect 12900 56772 12952 56778
rect 12900 56714 12952 56720
rect 14476 56710 14504 57190
rect 15028 57050 15056 57394
rect 17420 57050 17448 57394
rect 18880 57248 18932 57254
rect 18880 57190 18932 57196
rect 15016 57044 15068 57050
rect 15016 56986 15068 56992
rect 17408 57044 17460 57050
rect 17408 56986 17460 56992
rect 17224 56976 17276 56982
rect 17224 56918 17276 56924
rect 14464 56704 14516 56710
rect 14464 56646 14516 56652
rect 17236 56506 17264 56918
rect 17960 56908 18012 56914
rect 17960 56850 18012 56856
rect 17224 56500 17276 56506
rect 17224 56442 17276 56448
rect 17972 56438 18000 56850
rect 17960 56432 18012 56438
rect 17960 56374 18012 56380
rect 8300 55820 8352 55826
rect 8300 55762 8352 55768
rect 7012 55344 7064 55350
rect 7012 55286 7064 55292
rect 18892 54262 18920 57190
rect 19996 57050 20024 57394
rect 20536 57384 20588 57390
rect 20536 57326 20588 57332
rect 20076 57248 20128 57254
rect 20076 57190 20128 57196
rect 19984 57044 20036 57050
rect 19984 56986 20036 56992
rect 20088 56914 20116 57190
rect 20076 56908 20128 56914
rect 20076 56850 20128 56856
rect 19340 56840 19392 56846
rect 19340 56782 19392 56788
rect 19352 54670 19380 56782
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 20548 55758 20576 57326
rect 20732 56302 20760 57530
rect 20904 57520 20956 57526
rect 20904 57462 20956 57468
rect 20812 56772 20864 56778
rect 20812 56714 20864 56720
rect 20720 56296 20772 56302
rect 20720 56238 20772 56244
rect 20536 55752 20588 55758
rect 20536 55694 20588 55700
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 20824 55282 20852 56714
rect 20916 55962 20944 57462
rect 21008 57458 21036 59200
rect 22204 57458 22232 59200
rect 23400 57458 23428 59200
rect 24596 57458 24624 59200
rect 25792 57594 25820 59200
rect 26988 57594 27016 59200
rect 25780 57588 25832 57594
rect 25780 57530 25832 57536
rect 26976 57588 27028 57594
rect 26976 57530 27028 57536
rect 28184 57458 28212 59200
rect 29380 57594 29408 59200
rect 29368 57588 29420 57594
rect 29368 57530 29420 57536
rect 30576 57458 30604 59200
rect 31772 57458 31800 59200
rect 32968 57458 32996 59200
rect 34164 57594 34192 59200
rect 34152 57588 34204 57594
rect 34152 57530 34204 57536
rect 35360 57458 35388 59200
rect 36556 57458 36584 59200
rect 37752 57458 37780 59200
rect 38752 57588 38804 57594
rect 38752 57530 38804 57536
rect 20996 57452 21048 57458
rect 20996 57394 21048 57400
rect 22192 57452 22244 57458
rect 22192 57394 22244 57400
rect 23388 57452 23440 57458
rect 23388 57394 23440 57400
rect 24584 57452 24636 57458
rect 24584 57394 24636 57400
rect 28172 57452 28224 57458
rect 28172 57394 28224 57400
rect 30564 57452 30616 57458
rect 30564 57394 30616 57400
rect 31760 57452 31812 57458
rect 31760 57394 31812 57400
rect 32128 57452 32180 57458
rect 32128 57394 32180 57400
rect 32956 57452 33008 57458
rect 32956 57394 33008 57400
rect 35348 57452 35400 57458
rect 35348 57394 35400 57400
rect 36544 57452 36596 57458
rect 36544 57394 36596 57400
rect 37740 57452 37792 57458
rect 37740 57394 37792 57400
rect 21272 57248 21324 57254
rect 21272 57190 21324 57196
rect 21284 56846 21312 57190
rect 22204 57050 22232 57394
rect 24596 57050 24624 57394
rect 24952 57384 25004 57390
rect 24952 57326 25004 57332
rect 24860 57248 24912 57254
rect 24860 57190 24912 57196
rect 22192 57044 22244 57050
rect 22192 56986 22244 56992
rect 24584 57044 24636 57050
rect 24584 56986 24636 56992
rect 21272 56840 21324 56846
rect 21272 56782 21324 56788
rect 21180 56772 21232 56778
rect 21180 56714 21232 56720
rect 21192 56370 21220 56714
rect 24214 56400 24270 56409
rect 21180 56364 21232 56370
rect 21180 56306 21232 56312
rect 21916 56364 21968 56370
rect 21916 56306 21968 56312
rect 23756 56364 23808 56370
rect 24872 56370 24900 57190
rect 24964 56506 24992 57326
rect 25044 57316 25096 57322
rect 25044 57258 25096 57264
rect 24952 56500 25004 56506
rect 24952 56442 25004 56448
rect 24214 56335 24216 56344
rect 23756 56306 23808 56312
rect 24268 56335 24270 56344
rect 24860 56364 24912 56370
rect 24216 56306 24268 56312
rect 24860 56306 24912 56312
rect 20904 55956 20956 55962
rect 20904 55898 20956 55904
rect 21928 55622 21956 56306
rect 23388 56160 23440 56166
rect 23388 56102 23440 56108
rect 23572 56160 23624 56166
rect 23572 56102 23624 56108
rect 23400 55758 23428 56102
rect 23584 55758 23612 56102
rect 23664 55956 23716 55962
rect 23664 55898 23716 55904
rect 23676 55758 23704 55898
rect 23388 55752 23440 55758
rect 23388 55694 23440 55700
rect 23572 55752 23624 55758
rect 23572 55694 23624 55700
rect 23664 55752 23716 55758
rect 23664 55694 23716 55700
rect 21916 55616 21968 55622
rect 21916 55558 21968 55564
rect 21928 55282 21956 55558
rect 20812 55276 20864 55282
rect 20812 55218 20864 55224
rect 21916 55276 21968 55282
rect 21916 55218 21968 55224
rect 19340 54664 19392 54670
rect 19340 54606 19392 54612
rect 21928 54602 21956 55218
rect 21916 54596 21968 54602
rect 21916 54538 21968 54544
rect 23768 54534 23796 56306
rect 24584 56296 24636 56302
rect 24584 56238 24636 56244
rect 24596 55962 24624 56238
rect 24584 55956 24636 55962
rect 24584 55898 24636 55904
rect 23940 55888 23992 55894
rect 23940 55830 23992 55836
rect 22928 54528 22980 54534
rect 22928 54470 22980 54476
rect 23756 54528 23808 54534
rect 23756 54470 23808 54476
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 18880 54256 18932 54262
rect 18880 54198 18932 54204
rect 5724 53984 5776 53990
rect 5724 53926 5776 53932
rect 22940 53582 22968 54470
rect 22928 53576 22980 53582
rect 22928 53518 22980 53524
rect 5448 53440 5500 53446
rect 5448 53382 5500 53388
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 10600 53100 10652 53106
rect 10600 53042 10652 53048
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4804 51808 4856 51814
rect 4804 51750 4856 51756
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 3608 51060 3660 51066
rect 3608 51002 3660 51008
rect 2872 47592 2924 47598
rect 2872 47534 2924 47540
rect 3056 45824 3108 45830
rect 3056 45766 3108 45772
rect 2780 38752 2832 38758
rect 2780 38694 2832 38700
rect 2792 37806 2820 38694
rect 2780 37800 2832 37806
rect 2780 37742 2832 37748
rect 2688 32768 2740 32774
rect 2688 32710 2740 32716
rect 2700 26926 2728 32710
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 2792 27538 2820 27814
rect 3068 27538 3096 45766
rect 3424 28008 3476 28014
rect 3424 27950 3476 27956
rect 3436 27878 3464 27950
rect 3424 27872 3476 27878
rect 3424 27814 3476 27820
rect 2780 27532 2832 27538
rect 2780 27474 2832 27480
rect 3056 27532 3108 27538
rect 3056 27474 3108 27480
rect 2688 26920 2740 26926
rect 2688 26862 2740 26868
rect 2700 26382 2728 26862
rect 2792 26450 2820 27474
rect 3240 27396 3292 27402
rect 3240 27338 3292 27344
rect 3252 26994 3280 27338
rect 3332 27328 3384 27334
rect 3332 27270 3384 27276
rect 3344 26994 3372 27270
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 3252 26874 3280 26930
rect 3252 26846 3372 26874
rect 3344 26790 3372 26846
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 3332 26784 3384 26790
rect 3332 26726 3384 26732
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2688 26376 2740 26382
rect 2688 26318 2740 26324
rect 2688 26240 2740 26246
rect 2688 26182 2740 26188
rect 2700 26042 2728 26182
rect 2688 26036 2740 26042
rect 2688 25978 2740 25984
rect 2596 25424 2648 25430
rect 2424 25350 2544 25378
rect 2596 25366 2648 25372
rect 2412 25288 2464 25294
rect 2412 25230 2464 25236
rect 2424 24614 2452 25230
rect 2516 24834 2544 25350
rect 2516 24806 2636 24834
rect 2504 24744 2556 24750
rect 2504 24686 2556 24692
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2424 23798 2452 24550
rect 2412 23792 2464 23798
rect 2412 23734 2464 23740
rect 2412 23588 2464 23594
rect 2412 23530 2464 23536
rect 2320 23520 2372 23526
rect 2320 23462 2372 23468
rect 2332 23118 2360 23462
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2424 21622 2452 23530
rect 2148 21542 2268 21570
rect 2412 21616 2464 21622
rect 2412 21558 2464 21564
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 1952 20868 2004 20874
rect 1952 20810 2004 20816
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1674 19000 1730 19009
rect 1674 18935 1676 18944
rect 1728 18935 1730 18944
rect 1676 18906 1728 18912
rect 1872 18426 1900 19314
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 1964 18222 1992 20810
rect 1952 18216 2004 18222
rect 1674 18184 1730 18193
rect 1952 18158 2004 18164
rect 1674 18119 1730 18128
rect 1688 17882 1716 18119
rect 1964 17882 1992 18158
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1964 17134 1992 17818
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1964 16794 1992 17070
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1860 16584 1912 16590
rect 1674 16552 1730 16561
rect 2056 16574 2084 20878
rect 2148 19786 2176 21542
rect 2228 21480 2280 21486
rect 2228 21422 2280 21428
rect 2240 21146 2268 21422
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2240 20466 2268 21082
rect 2332 20942 2360 21286
rect 2424 20942 2452 21558
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 2412 20936 2464 20942
rect 2412 20878 2464 20884
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2136 19780 2188 19786
rect 2136 19722 2188 19728
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2424 18850 2452 19654
rect 2516 18970 2544 24686
rect 2608 22710 2636 24806
rect 2792 24274 2820 26386
rect 2884 25906 2912 26726
rect 2964 26240 3016 26246
rect 2964 26182 3016 26188
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2976 25294 3004 26182
rect 3344 26042 3372 26726
rect 3240 26036 3292 26042
rect 3240 25978 3292 25984
rect 3332 26036 3384 26042
rect 3332 25978 3384 25984
rect 3252 25702 3280 25978
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 2964 25288 3016 25294
rect 2964 25230 3016 25236
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2792 23866 2820 24210
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2792 22982 2820 23666
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2596 22704 2648 22710
rect 2596 22646 2648 22652
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2332 18822 2452 18850
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 1860 16526 1912 16532
rect 1964 16546 2084 16574
rect 1674 16487 1730 16496
rect 1688 16454 1716 16487
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1872 15910 1900 16526
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1674 14920 1730 14929
rect 1674 14855 1730 14864
rect 1688 14618 1716 14855
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1860 13320 1912 13326
rect 1674 13288 1730 13297
rect 1860 13262 1912 13268
rect 1674 13223 1730 13232
rect 1688 13190 1716 13223
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1872 12714 1900 13262
rect 1964 13002 1992 16546
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2056 15638 2084 16050
rect 2044 15632 2096 15638
rect 2044 15574 2096 15580
rect 2240 15450 2268 18702
rect 2332 16590 2360 18822
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2424 18426 2452 18702
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2424 17377 2452 17478
rect 2410 17368 2466 17377
rect 2410 17303 2466 17312
rect 2320 16584 2372 16590
rect 2516 16574 2544 17614
rect 2320 16526 2372 16532
rect 2424 16546 2544 16574
rect 2056 15422 2268 15450
rect 2056 13938 2084 15422
rect 2424 15314 2452 16546
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 15706 2544 16390
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2240 15286 2452 15314
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2148 13870 2176 15030
rect 2240 14958 2268 15286
rect 2516 15094 2544 15642
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2148 13462 2176 13806
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 2240 13138 2268 14894
rect 2608 14550 2636 22374
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2700 20602 2728 22034
rect 2688 20596 2740 20602
rect 2688 20538 2740 20544
rect 2700 19922 2728 20538
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2700 17270 2728 17614
rect 2792 17338 2820 22714
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2688 17264 2740 17270
rect 2688 17206 2740 17212
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2700 16590 2728 16730
rect 2688 16584 2740 16590
rect 2792 16574 2820 17274
rect 2792 16546 3004 16574
rect 2688 16526 2740 16532
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2700 16250 2728 16390
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2424 14113 2452 14214
rect 2410 14104 2466 14113
rect 2410 14039 2466 14048
rect 2700 13938 2728 14758
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13326 2360 13670
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2240 13110 2360 13138
rect 1964 12974 2084 13002
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12481 1716 12582
rect 1674 12472 1730 12481
rect 1674 12407 1730 12416
rect 1964 12102 1992 12786
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1674 11656 1730 11665
rect 1674 11591 1676 11600
rect 1728 11591 1730 11600
rect 1676 11562 1728 11568
rect 1674 10840 1730 10849
rect 1674 10775 1730 10784
rect 1688 10266 1716 10775
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1674 10024 1730 10033
rect 1674 9959 1730 9968
rect 1688 9450 1716 9959
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1674 9208 1730 9217
rect 1674 9143 1676 9152
rect 1728 9143 1730 9152
rect 1676 9114 1728 9120
rect 1674 8392 1730 8401
rect 1674 8327 1730 8336
rect 1688 8090 1716 8327
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1674 6760 1730 6769
rect 1674 6695 1730 6704
rect 1688 6458 1716 6695
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1674 5944 1730 5953
rect 1674 5879 1676 5888
rect 1728 5879 1730 5888
rect 1676 5850 1728 5856
rect 1674 5128 1730 5137
rect 1674 5063 1676 5072
rect 1728 5063 1730 5072
rect 1676 5034 1728 5040
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1688 4321 1716 4422
rect 1674 4312 1730 4321
rect 1674 4247 1730 4256
rect 1872 3670 1900 4558
rect 1860 3664 1912 3670
rect 1860 3606 1912 3612
rect 1964 2854 1992 12038
rect 2056 10198 2084 12974
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2148 10606 2176 11154
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2044 10192 2096 10198
rect 2044 10134 2096 10140
rect 2240 9450 2268 11018
rect 2332 10470 2360 13110
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 11354 2452 11494
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2516 11150 2544 11766
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2424 9518 2452 9998
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2240 8974 2268 9386
rect 2516 9110 2544 10542
rect 2700 10538 2728 11562
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2700 9926 2728 10474
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 9722 2728 9862
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2700 9178 2728 9658
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2148 7342 2176 8298
rect 2240 8090 2268 8366
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2148 6866 2176 7278
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2240 6322 2268 8026
rect 2516 7954 2544 9046
rect 2700 8362 2728 9114
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2700 8022 2728 8298
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2332 6662 2360 7822
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7585 2452 7686
rect 2410 7576 2466 7585
rect 2792 7562 2820 13942
rect 2700 7546 2912 7562
rect 2410 7511 2466 7520
rect 2688 7540 2924 7546
rect 2740 7534 2872 7540
rect 2688 7482 2740 7488
rect 2872 7482 2924 7488
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2516 6798 2544 7278
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 6458 2360 6598
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2516 5710 2544 6734
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 6322 2820 6598
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2884 6118 2912 6802
rect 2872 6112 2924 6118
rect 2792 6060 2872 6066
rect 2792 6054 2924 6060
rect 2792 6038 2912 6054
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2424 4078 2452 5170
rect 2792 4486 2820 6038
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3058 2268 3878
rect 2424 3194 2452 4014
rect 2792 4010 2820 4422
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2792 3602 2820 3946
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2792 3126 2820 3538
rect 2976 3466 3004 16546
rect 3068 15570 3096 25638
rect 3252 21554 3280 25638
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3252 21350 3280 21490
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3160 15026 3188 19246
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3160 14822 3188 14962
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3068 10266 3096 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3160 4298 3188 14758
rect 3252 6662 3280 21286
rect 3344 18970 3372 25978
rect 3516 24608 3568 24614
rect 3516 24550 3568 24556
rect 3528 24410 3556 24550
rect 3516 24404 3568 24410
rect 3516 24346 3568 24352
rect 3424 24268 3476 24274
rect 3424 24210 3476 24216
rect 3436 24154 3464 24210
rect 3436 24126 3556 24154
rect 3528 24070 3556 24126
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3436 23118 3464 24006
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3344 18358 3372 18906
rect 3620 18834 3648 51002
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4712 47456 4764 47462
rect 4712 47398 4764 47404
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 3976 43648 4028 43654
rect 3976 43590 4028 43596
rect 3792 28756 3844 28762
rect 3792 28698 3844 28704
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3712 24342 3740 24754
rect 3700 24336 3752 24342
rect 3700 24278 3752 24284
rect 3700 24132 3752 24138
rect 3700 24074 3752 24080
rect 3712 22778 3740 24074
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3332 18352 3384 18358
rect 3332 18294 3384 18300
rect 3344 16574 3372 18294
rect 3620 18222 3648 18770
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3804 16574 3832 28698
rect 3884 27464 3936 27470
rect 3884 27406 3936 27412
rect 3896 19854 3924 27406
rect 3988 24070 4016 43590
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4620 37800 4672 37806
rect 4620 37742 4672 37748
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 4080 28014 4108 28358
rect 4068 28008 4120 28014
rect 4068 27950 4120 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27532 4120 27538
rect 4068 27474 4120 27480
rect 4080 24614 4108 27474
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3988 22982 4016 23598
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3896 19310 3924 19790
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3344 16546 3464 16574
rect 3804 16546 3924 16574
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3160 4270 3280 4298
rect 3252 4214 3280 4270
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3252 3942 3280 4150
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2976 3058 3004 3402
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2332 800 2360 2382
rect 3252 2038 3280 3878
rect 3240 2032 3292 2038
rect 3240 1974 3292 1980
rect 3344 1902 3372 10202
rect 3436 8634 3464 16546
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3804 14618 3832 14758
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3896 14006 3924 16546
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3988 10266 4016 22918
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16266 4660 37742
rect 4724 28218 4752 47398
rect 4816 35894 4844 51750
rect 9588 45280 9640 45286
rect 9588 45222 9640 45228
rect 6184 44192 6236 44198
rect 6184 44134 6236 44140
rect 4816 35866 4936 35894
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4724 16561 4752 26726
rect 4816 25702 4844 26930
rect 4804 25696 4856 25702
rect 4804 25638 4856 25644
rect 4908 23730 4936 35866
rect 5908 29028 5960 29034
rect 5908 28970 5960 28976
rect 5920 28626 5948 28970
rect 5908 28620 5960 28626
rect 5908 28562 5960 28568
rect 5264 27940 5316 27946
rect 5264 27882 5316 27888
rect 5172 27872 5224 27878
rect 5172 27814 5224 27820
rect 5184 27470 5212 27814
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 4988 24880 5040 24886
rect 4988 24822 5040 24828
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4896 23248 4948 23254
rect 4896 23190 4948 23196
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4816 16998 4844 22918
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4710 16552 4766 16561
rect 4710 16487 4766 16496
rect 4632 16238 4844 16266
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14550 4660 15982
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4816 11558 4844 16238
rect 4908 15366 4936 23190
rect 5000 20874 5028 24822
rect 5172 24064 5224 24070
rect 5172 24006 5224 24012
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 5000 20534 5028 20810
rect 4988 20528 5040 20534
rect 4988 20470 5040 20476
rect 5000 19854 5028 20470
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 5000 18442 5028 19654
rect 5184 18578 5212 24006
rect 5276 18766 5304 27882
rect 5920 27690 5948 28562
rect 6000 28552 6052 28558
rect 6000 28494 6052 28500
rect 6012 28082 6040 28494
rect 6196 28218 6224 44134
rect 7564 40928 7616 40934
rect 7564 40870 7616 40876
rect 6276 40384 6328 40390
rect 6276 40326 6328 40332
rect 6288 35222 6316 40326
rect 6276 35216 6328 35222
rect 6276 35158 6328 35164
rect 6920 34536 6972 34542
rect 6920 34478 6972 34484
rect 6828 28960 6880 28966
rect 6828 28902 6880 28908
rect 6840 28558 6868 28902
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6932 28490 6960 34478
rect 6920 28484 6972 28490
rect 6920 28426 6972 28432
rect 7104 28484 7156 28490
rect 7104 28426 7156 28432
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6460 28144 6512 28150
rect 6460 28086 6512 28092
rect 6000 28076 6052 28082
rect 6000 28018 6052 28024
rect 5828 27662 5948 27690
rect 6012 27674 6040 28018
rect 6000 27668 6052 27674
rect 5356 27464 5408 27470
rect 5356 27406 5408 27412
rect 5368 26926 5396 27406
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 5356 26920 5408 26926
rect 5356 26862 5408 26868
rect 5368 26450 5396 26862
rect 5356 26444 5408 26450
rect 5356 26386 5408 26392
rect 5368 26042 5396 26386
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 5184 18550 5304 18578
rect 5000 18414 5212 18442
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16658 5120 16934
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 4986 16552 5042 16561
rect 4986 16487 5042 16496
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 5000 12442 5028 16487
rect 5184 14618 5212 18414
rect 5276 16454 5304 18550
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5276 14618 5304 14758
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5184 11898 5212 14282
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4816 11234 4844 11494
rect 4632 11206 4844 11234
rect 4632 11150 4660 11206
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 5184 11082 5212 11834
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5184 10742 5212 11018
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 5184 9994 5212 10678
rect 5276 10606 5304 14010
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5172 9988 5224 9994
rect 5172 9930 5224 9936
rect 5184 9654 5212 9930
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4080 9042 4108 9522
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5184 9178 5212 9590
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3436 8430 3464 8570
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3436 7002 3464 7142
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 3436 800 3464 3538
rect 3528 1766 3556 6598
rect 3988 2514 4016 7482
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4080 2310 4108 8570
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5368 6730 5396 7754
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5368 6458 5396 6666
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 5460 4826 5488 27270
rect 5828 27062 5856 27662
rect 6000 27610 6052 27616
rect 6012 27554 6040 27610
rect 5920 27526 6040 27554
rect 5816 27056 5868 27062
rect 5816 26998 5868 27004
rect 5632 26512 5684 26518
rect 5632 26454 5684 26460
rect 5540 26308 5592 26314
rect 5540 26250 5592 26256
rect 5552 21434 5580 26250
rect 5644 25514 5672 26454
rect 5644 25486 5856 25514
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 5736 24818 5764 25298
rect 5724 24812 5776 24818
rect 5724 24754 5776 24760
rect 5552 21406 5672 21434
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5552 17134 5580 18226
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5552 16522 5580 17070
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5552 15434 5580 16458
rect 5644 15706 5672 21406
rect 5736 21010 5764 24754
rect 5828 21146 5856 25486
rect 5920 23662 5948 27526
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 6012 25906 6040 26726
rect 6368 26512 6420 26518
rect 6368 26454 6420 26460
rect 6380 26314 6408 26454
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6000 25900 6052 25906
rect 6000 25842 6052 25848
rect 6380 25770 6408 26250
rect 6368 25764 6420 25770
rect 6368 25706 6420 25712
rect 6000 25220 6052 25226
rect 6000 25162 6052 25168
rect 5908 23656 5960 23662
rect 5908 23598 5960 23604
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5724 21004 5776 21010
rect 5724 20946 5776 20952
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5828 20262 5856 20402
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5828 17202 5856 20198
rect 6012 18698 6040 25162
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6104 23662 6132 24278
rect 6184 23724 6236 23730
rect 6184 23666 6236 23672
rect 6092 23656 6144 23662
rect 6092 23598 6144 23604
rect 6196 19990 6224 23666
rect 6380 22794 6408 25706
rect 6288 22766 6408 22794
rect 6184 19984 6236 19990
rect 6184 19926 6236 19932
rect 6000 18692 6052 18698
rect 6000 18634 6052 18640
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5920 16658 5948 18158
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 6288 11830 6316 22766
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6380 16998 6408 17138
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5828 9654 5856 11154
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 6012 10606 6040 11018
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6012 10130 6040 10542
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 6012 9654 6040 9930
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5920 7954 5948 8298
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6012 6254 6040 7754
rect 6288 6914 6316 11766
rect 6380 9178 6408 16934
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6380 8974 6408 9114
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6380 8634 6408 8910
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6196 6886 6316 6914
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6012 5114 6040 6190
rect 5920 5086 6040 5114
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 4150
rect 5920 3534 5948 5086
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5184 3194 5212 3402
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 3516 1760 3568 1766
rect 3516 1702 3568 1708
rect 4540 800 4568 2382
rect 4816 2106 4844 2586
rect 4908 2582 4936 3130
rect 5920 3058 5948 3470
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 5644 800 5672 2382
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5920 1970 5948 2246
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 6196 1834 6224 6886
rect 6380 4078 6408 8570
rect 6472 4690 6500 28086
rect 6840 28082 6868 28358
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6656 18426 6684 27066
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6840 18630 6868 25638
rect 6920 25220 6972 25226
rect 6920 25162 6972 25168
rect 6932 24818 6960 25162
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 7116 22098 7144 28426
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6748 18154 6776 18362
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 7116 18086 7144 18226
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6564 14482 6592 16186
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6748 11286 6776 16186
rect 7576 15366 7604 40870
rect 7656 39296 7708 39302
rect 7656 39238 7708 39244
rect 7668 35894 7696 39238
rect 8484 36168 8536 36174
rect 8484 36110 8536 36116
rect 7668 35866 7788 35894
rect 7656 28960 7708 28966
rect 7656 28902 7708 28908
rect 7668 28558 7696 28902
rect 7656 28552 7708 28558
rect 7656 28494 7708 28500
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7668 26518 7696 26862
rect 7656 26512 7708 26518
rect 7656 26454 7708 26460
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 18358 7696 19246
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7668 18086 7696 18294
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7668 17610 7696 18022
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7760 17338 7788 35866
rect 8496 29306 8524 36110
rect 9220 29572 9272 29578
rect 9220 29514 9272 29520
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 7932 28756 7984 28762
rect 7852 28716 7932 28744
rect 7852 28014 7880 28716
rect 7932 28698 7984 28704
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 7840 28008 7892 28014
rect 7840 27950 7892 27956
rect 8128 27606 8156 28018
rect 8116 27600 8168 27606
rect 8116 27542 8168 27548
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8404 26314 8432 26522
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 8300 25492 8352 25498
rect 8300 25434 8352 25440
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8220 19446 8248 24754
rect 8312 21146 8340 25434
rect 8404 24750 8432 26250
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8496 22778 8524 29242
rect 8760 28688 8812 28694
rect 8760 28630 8812 28636
rect 8576 27872 8628 27878
rect 8576 27814 8628 27820
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8312 20602 8340 20946
rect 8404 20806 8432 22646
rect 8588 22234 8616 27814
rect 8772 22574 8800 28630
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9140 27470 9168 28358
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9036 27328 9088 27334
rect 9036 27270 9088 27276
rect 8760 22568 8812 22574
rect 8760 22510 8812 22516
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8312 19922 8340 20538
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8312 19378 8340 19858
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 9048 19310 9076 27270
rect 9128 26784 9180 26790
rect 9128 26726 9180 26732
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 8128 18358 8156 18566
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6840 11218 6868 11494
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 9518 6960 10066
rect 7300 9994 7328 15302
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 7668 5030 7696 15846
rect 8404 15706 8432 17206
rect 8680 16046 8708 18158
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6380 3466 6408 4014
rect 8036 3466 8064 15642
rect 8680 15502 8708 15982
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8312 14822 8340 15438
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8312 14482 8340 14758
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9110 8248 9318
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8956 6914 8984 14214
rect 9140 11694 9168 26726
rect 9232 25770 9260 29514
rect 9600 28626 9628 45222
rect 9772 29572 9824 29578
rect 9772 29514 9824 29520
rect 9784 29102 9812 29514
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 9956 29028 10008 29034
rect 9956 28970 10008 28976
rect 9772 28688 9824 28694
rect 9772 28630 9824 28636
rect 9588 28620 9640 28626
rect 9588 28562 9640 28568
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 9508 28150 9536 28494
rect 9496 28144 9548 28150
rect 9496 28086 9548 28092
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9220 25764 9272 25770
rect 9220 25706 9272 25712
rect 9692 25498 9720 27814
rect 9784 26994 9812 28630
rect 9864 27396 9916 27402
rect 9864 27338 9916 27344
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9784 24750 9812 26250
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9232 12442 9260 24550
rect 9876 17882 9904 27338
rect 9968 26994 9996 28970
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10416 27600 10468 27606
rect 10416 27542 10468 27548
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 10428 26450 10456 27542
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 9956 26308 10008 26314
rect 9956 26250 10008 26256
rect 9968 23050 9996 26250
rect 10428 25702 10456 26386
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10060 24274 10088 24686
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 10060 22642 10088 24210
rect 10428 23526 10456 25638
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10060 21010 10088 22578
rect 10416 22432 10468 22438
rect 10416 22374 10468 22380
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 10060 19922 10088 20946
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9416 15570 9444 17002
rect 9692 16046 9720 17546
rect 10428 16250 10456 22374
rect 10520 19514 10548 28494
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 10060 15434 10088 16050
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9600 13530 9628 14282
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9324 11762 9352 12242
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9048 9722 9076 10066
rect 9324 10062 9352 11698
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9324 9722 9352 9998
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9324 9042 9352 9658
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9324 7546 9352 8978
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 8956 6886 9076 6914
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8588 6118 8616 6734
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4826 8616 4966
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8312 3534 8340 4490
rect 9048 4146 9076 6886
rect 9416 6730 9444 12106
rect 10612 10742 10640 53042
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19064 50380 19116 50386
rect 19064 50322 19116 50328
rect 10784 49224 10836 49230
rect 10784 49166 10836 49172
rect 10796 29306 10824 49166
rect 15200 47592 15252 47598
rect 15200 47534 15252 47540
rect 14464 42220 14516 42226
rect 14464 42162 14516 42168
rect 13636 37460 13688 37466
rect 13636 37402 13688 37408
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 11060 30252 11112 30258
rect 11060 30194 11112 30200
rect 11072 30054 11100 30194
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11428 30048 11480 30054
rect 11428 29990 11480 29996
rect 10784 29300 10836 29306
rect 10784 29242 10836 29248
rect 10968 29028 11020 29034
rect 10968 28970 11020 28976
rect 10980 28626 11008 28970
rect 10968 28620 11020 28626
rect 10968 28562 11020 28568
rect 10980 27878 11008 28562
rect 11072 28150 11100 29990
rect 11152 29708 11204 29714
rect 11152 29650 11204 29656
rect 11164 29170 11192 29650
rect 11440 29646 11468 29990
rect 11428 29640 11480 29646
rect 11428 29582 11480 29588
rect 11244 29504 11296 29510
rect 11244 29446 11296 29452
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11164 28422 11192 29106
rect 11152 28416 11204 28422
rect 11152 28358 11204 28364
rect 11060 28144 11112 28150
rect 11060 28086 11112 28092
rect 10968 27872 11020 27878
rect 10968 27814 11020 27820
rect 10784 27396 10836 27402
rect 10784 27338 10836 27344
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 10704 24274 10732 26726
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10796 21978 10824 27338
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 10888 26382 10916 27270
rect 10980 27062 11008 27814
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11072 27334 11100 27406
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 11072 27130 11100 27270
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 11164 26314 11192 28358
rect 11152 26308 11204 26314
rect 11152 26250 11204 26256
rect 10876 23044 10928 23050
rect 10876 22986 10928 22992
rect 10704 21962 10824 21978
rect 10692 21956 10824 21962
rect 10744 21950 10824 21956
rect 10692 21898 10744 21904
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 9518 9720 10406
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9416 5642 9444 6666
rect 9600 6390 9628 7346
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5710 9536 6054
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9416 5302 9444 5578
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9416 4554 9444 5238
rect 9508 5030 9536 5646
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10336 5030 10364 5102
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 9508 4690 9536 4966
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 8300 3528 8352 3534
rect 8352 3476 8432 3482
rect 8300 3470 8432 3476
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 8024 3460 8076 3466
rect 8312 3454 8432 3470
rect 8024 3402 8076 3408
rect 6380 3194 6408 3402
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 7300 2446 7328 3334
rect 8036 3194 8064 3402
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8404 3058 8432 3454
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 6920 2440 6972 2446
rect 6748 2400 6920 2428
rect 6184 1828 6236 1834
rect 6184 1770 6236 1776
rect 6748 800 6776 2400
rect 6920 2382 6972 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7852 2378 7880 2790
rect 8956 2378 8984 3334
rect 9508 3126 9536 3946
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 10336 3058 10364 4966
rect 10704 3738 10732 21898
rect 10888 19514 10916 22986
rect 11256 19922 11284 29446
rect 11716 28558 11744 35634
rect 12440 32428 12492 32434
rect 12440 32370 12492 32376
rect 12452 30326 12480 32370
rect 12440 30320 12492 30326
rect 12440 30262 12492 30268
rect 12624 30320 12676 30326
rect 12624 30262 12676 30268
rect 12348 30184 12400 30190
rect 12348 30126 12400 30132
rect 12360 29510 12388 30126
rect 12348 29504 12400 29510
rect 12348 29446 12400 29452
rect 11980 29300 12032 29306
rect 11980 29242 12032 29248
rect 11704 28552 11756 28558
rect 11704 28494 11756 28500
rect 11716 28150 11744 28494
rect 11428 28144 11480 28150
rect 11428 28086 11480 28092
rect 11704 28144 11756 28150
rect 11704 28086 11756 28092
rect 11336 27532 11388 27538
rect 11336 27474 11388 27480
rect 11348 27062 11376 27474
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 11440 26874 11468 28086
rect 11348 26846 11468 26874
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13870 11100 14214
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 7546 10916 12650
rect 11348 11898 11376 26846
rect 11428 26512 11480 26518
rect 11428 26454 11480 26460
rect 11440 17746 11468 26454
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11808 24206 11836 25162
rect 11992 24410 12020 29242
rect 12360 28626 12388 29446
rect 12348 28620 12400 28626
rect 12348 28562 12400 28568
rect 12164 28416 12216 28422
rect 12164 28358 12216 28364
rect 12072 28212 12124 28218
rect 12072 28154 12124 28160
rect 12084 25226 12112 28154
rect 12176 26926 12204 28358
rect 12360 28218 12388 28562
rect 12348 28212 12400 28218
rect 12348 28154 12400 28160
rect 12256 27328 12308 27334
rect 12256 27270 12308 27276
rect 12268 26994 12296 27270
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 12164 26920 12216 26926
rect 12164 26862 12216 26868
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 12072 25220 12124 25226
rect 12072 25162 12124 25168
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 11900 20534 11928 20742
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11532 15978 11560 18634
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11992 17338 12020 17818
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 8922 11100 9862
rect 10980 8906 11100 8922
rect 10968 8900 11100 8906
rect 11020 8894 11100 8900
rect 10968 8842 11020 8848
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 11532 5778 11560 15914
rect 11612 14340 11664 14346
rect 11612 14282 11664 14288
rect 11624 13870 11652 14282
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 11624 3602 11652 13806
rect 12176 10062 12204 26250
rect 12360 25906 12388 26522
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12360 20534 12388 21830
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12452 21350 12480 21490
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12348 20528 12400 20534
rect 12348 20470 12400 20476
rect 12360 19922 12388 20470
rect 12452 20330 12480 21286
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12452 15910 12480 20266
rect 12636 19990 12664 30262
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13556 27606 13584 27814
rect 13544 27600 13596 27606
rect 13544 27542 13596 27548
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 13004 26926 13032 27270
rect 12992 26920 13044 26926
rect 12992 26862 13044 26868
rect 13360 26852 13412 26858
rect 13360 26794 13412 26800
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 15910 12848 16050
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12360 15162 12388 15302
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12360 14414 12388 15098
rect 12820 14890 12848 15846
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12820 14278 12848 14826
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12636 14006 12664 14214
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12636 12170 12664 13942
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11354 12388 11494
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 10130 12572 10406
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12176 9178 12204 9862
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12820 8566 12848 14214
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12912 8634 12940 8910
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12820 7410 12848 8502
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12820 5370 12848 7346
rect 13096 5914 13124 16730
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13188 9178 13216 12106
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13188 8906 13216 9114
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11716 3194 11744 4014
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 12176 3126 12204 3402
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 10060 2378 10088 2790
rect 11164 2378 11192 2790
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 7852 800 7880 2314
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8128 2038 8156 2246
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 8956 800 8984 2314
rect 10060 800 10088 2314
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 1766 11008 2246
rect 10968 1760 11020 1766
rect 10968 1702 11020 1708
rect 11164 800 11192 2314
rect 12176 1902 12204 2382
rect 12268 2258 12296 3878
rect 13280 3670 13308 14554
rect 13372 3738 13400 26794
rect 13452 26784 13504 26790
rect 13452 26726 13504 26732
rect 13464 6390 13492 26726
rect 13648 24614 13676 37402
rect 14476 30326 14504 42162
rect 14464 30320 14516 30326
rect 14464 30262 14516 30268
rect 15016 29232 15068 29238
rect 15016 29174 15068 29180
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14924 27328 14976 27334
rect 14924 27270 14976 27276
rect 14292 26994 14320 27270
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 14096 25764 14148 25770
rect 14096 25706 14148 25712
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13924 22710 13952 24142
rect 13912 22704 13964 22710
rect 13912 22646 13964 22652
rect 13924 20534 13952 22646
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13832 18426 13860 19450
rect 13924 19446 13952 20470
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 17338 13860 17614
rect 13924 17610 13952 19382
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13832 17202 13860 17274
rect 13924 17270 13952 17546
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13832 15910 13860 17138
rect 14108 17066 14136 25706
rect 14188 25696 14240 25702
rect 14188 25638 14240 25644
rect 14200 19310 14228 25638
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 14292 20602 14320 23734
rect 14844 23050 14872 24822
rect 14936 24342 14964 27270
rect 15028 26234 15056 29174
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15120 27130 15148 27474
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15028 26206 15148 26234
rect 14924 24336 14976 24342
rect 14924 24278 14976 24284
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14844 21894 14872 22986
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14372 21412 14424 21418
rect 14372 21354 14424 21360
rect 14384 21146 14412 21354
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14292 17542 14320 20538
rect 14384 20346 14412 21082
rect 14844 20874 14872 21830
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14384 20318 14504 20346
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14384 19718 14412 20198
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14476 18358 14504 20318
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14096 17060 14148 17066
rect 14096 17002 14148 17008
rect 14108 16658 14136 17002
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13832 14958 13860 15098
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 14384 14278 14412 14962
rect 14476 14958 14504 15846
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11830 13768 12106
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13556 10742 13584 10950
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13832 9654 13860 10678
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13464 6254 13492 6326
rect 13556 6254 13584 9318
rect 13832 7818 13860 9590
rect 14384 9178 14412 14214
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 10810 14504 11630
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14476 9518 14504 10746
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14384 8974 14412 9114
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14476 8634 14504 9454
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13832 7562 13860 7754
rect 13832 7534 13952 7562
rect 13924 7478 13952 7534
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13924 6390 13952 7414
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13924 4214 13952 6326
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13924 3058 13952 4150
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13832 2446 13860 2790
rect 14660 2650 14688 9862
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14752 5166 14780 6394
rect 14936 6254 14964 24278
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15028 15094 15056 17546
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 11694 15056 13806
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15120 10266 15148 26206
rect 15212 17746 15240 47534
rect 17408 44872 17460 44878
rect 17408 44814 17460 44820
rect 15936 42696 15988 42702
rect 15936 42638 15988 42644
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15396 24818 15424 25230
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 22574 15424 24754
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15396 22098 15424 22510
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15396 21622 15424 22034
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15396 21010 15424 21558
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15396 19378 15424 20946
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15672 8294 15700 30262
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15764 13734 15792 27814
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15856 12374 15884 18702
rect 15948 13530 15976 42638
rect 16580 36916 16632 36922
rect 16580 36858 16632 36864
rect 16028 35216 16080 35222
rect 16028 35158 16080 35164
rect 16040 23322 16068 35158
rect 16592 28762 16620 36858
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16592 28150 16620 28698
rect 16580 28144 16632 28150
rect 16632 28092 16712 28098
rect 16580 28086 16712 28092
rect 16592 28070 16712 28086
rect 16212 26920 16264 26926
rect 16212 26862 16264 26868
rect 16224 25158 16252 26862
rect 16580 26240 16632 26246
rect 16580 26182 16632 26188
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16500 22574 16528 23122
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16592 22506 16620 26182
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 16132 20466 16160 20946
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 15856 11830 15884 12310
rect 16040 12170 16068 13126
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 16040 9994 16068 12106
rect 16224 11218 16252 21898
rect 16316 16182 16344 22170
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16684 14074 16712 28070
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17236 27402 17264 28018
rect 17224 27396 17276 27402
rect 17224 27338 17276 27344
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 17052 25906 17080 26726
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16868 25362 16896 25638
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 17224 24676 17276 24682
rect 17224 24618 17276 24624
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 16960 18970 16988 20810
rect 17236 20262 17264 24618
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17052 16998 17080 18566
rect 17144 18426 17172 18702
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 17328 18154 17356 20334
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17236 17338 17264 17614
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17328 16794 17356 17002
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17420 16574 17448 44814
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 18064 27062 18092 27270
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18052 27056 18104 27062
rect 18052 26998 18104 27004
rect 18064 26926 18092 26998
rect 18052 26920 18104 26926
rect 18052 26862 18104 26868
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17972 23594 18000 26250
rect 18064 24410 18092 26862
rect 18248 26450 18276 27066
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 18248 25702 18276 26386
rect 18524 26382 18552 26726
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 18524 26246 18552 26318
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18524 25974 18552 26182
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18052 24404 18104 24410
rect 18052 24346 18104 24352
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 18144 22500 18196 22506
rect 18144 22442 18196 22448
rect 18156 22234 18184 22442
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17604 17882 17632 20198
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 17338 17632 17478
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17420 16546 17540 16574
rect 17512 14822 17540 16546
rect 17696 16250 17724 17070
rect 17788 16794 17816 17546
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 18064 16574 18092 20198
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18834 18184 19110
rect 18248 18834 18276 25638
rect 18340 25158 18368 25842
rect 18524 25702 18552 25910
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18340 24614 18368 25094
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18432 23050 18460 23462
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18524 22930 18552 25638
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18708 24750 18736 25094
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18800 24206 18828 24550
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 18432 22902 18552 22930
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18156 17882 18184 18226
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18064 16546 18184 16574
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17512 14074 17540 14758
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16684 12306 16712 13262
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16960 12986 16988 13194
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16684 10810 16712 12242
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16684 10690 16712 10746
rect 16684 10662 16804 10690
rect 16776 10130 16804 10662
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15672 7954 15700 8230
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 16868 5166 16896 7346
rect 17788 6662 17816 9590
rect 17880 9450 17908 9930
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7410 17908 7822
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 4690 16896 5102
rect 18156 4690 18184 16546
rect 18432 10538 18460 22902
rect 18616 22778 18644 23530
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 19076 21690 19104 50322
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18708 21350 18736 21490
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18708 20534 18736 21286
rect 18880 21140 18932 21146
rect 18880 21082 18932 21088
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 18708 19718 18736 20470
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 18698 18736 19654
rect 18800 18766 18828 20198
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18524 17218 18552 17682
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 17338 18644 17478
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18524 17190 18644 17218
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18524 14618 18552 16594
rect 18616 16046 18644 17190
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18800 16250 18828 16526
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18616 15706 18644 15982
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 15162 18736 15302
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18708 11354 18736 12106
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18524 10674 18552 11290
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14752 4214 14780 4490
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14752 3534 14780 4150
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 3126 14780 3470
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 15580 2446 15608 4422
rect 16868 4214 16896 4626
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15672 3058 15700 3538
rect 15948 3398 15976 4014
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15856 3126 15884 3334
rect 15844 3120 15896 3126
rect 15844 3062 15896 3068
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 12452 2258 12480 2382
rect 12268 2230 12480 2258
rect 12164 1896 12216 1902
rect 12164 1838 12216 1844
rect 12268 800 12296 2230
rect 13372 800 13400 2382
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13648 1834 13676 2246
rect 13636 1828 13688 1834
rect 13636 1770 13688 1776
rect 14476 800 14504 2382
rect 15580 800 15608 2382
rect 16684 2378 16712 3878
rect 16868 3602 16896 4150
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18064 3942 18092 4014
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 18064 3058 18092 3878
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 16684 800 16712 2314
rect 17788 800 17816 2926
rect 18248 2582 18276 10406
rect 18524 10266 18552 10610
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18708 2650 18736 6190
rect 18800 5914 18828 7278
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18892 4690 18920 21082
rect 18984 20466 19012 21286
rect 19076 21146 19104 21626
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19168 17678 19196 21966
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19168 17338 19196 17614
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 18984 4758 19012 17274
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19076 10266 19104 10542
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19260 6458 19288 27338
rect 19444 25838 19472 27814
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 19628 25294 19656 25638
rect 19616 25288 19668 25294
rect 19616 25230 19668 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19352 24138 19380 24550
rect 19628 24410 19656 24754
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 20260 24268 20312 24274
rect 20260 24210 20312 24216
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19352 19922 19380 24074
rect 20272 24070 20300 24210
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23866 20024 24006
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19444 23322 19472 23666
rect 19996 23610 20024 23802
rect 19996 23582 20208 23610
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 20088 23186 20116 23462
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19444 22234 19472 22510
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19444 19718 19472 20334
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19352 18426 19380 19314
rect 19996 19310 20024 22918
rect 20088 22098 20116 23122
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 20180 22030 20208 23582
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20272 21350 20300 24006
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19352 17746 19380 18158
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19444 17202 19472 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19536 17882 19564 18362
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19352 14618 19380 16118
rect 19996 16046 20024 18566
rect 20180 16574 20208 19654
rect 20272 19242 20300 21286
rect 20364 20534 20392 25638
rect 20628 22092 20680 22098
rect 20628 22034 20680 22040
rect 20640 21894 20668 22034
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20640 20466 20668 21830
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20260 19236 20312 19242
rect 20260 19178 20312 19184
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20272 18086 20300 18634
rect 20548 18222 20576 18770
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20088 16546 20208 16574
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19444 15910 19472 15982
rect 19432 15904 19484 15910
rect 20088 15858 20116 16546
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 19432 15846 19484 15852
rect 19996 15830 20116 15858
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19444 15162 19472 15438
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19904 14618 19932 15030
rect 19996 14822 20024 15830
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 20088 14958 20116 15302
rect 20180 15094 20208 16050
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19444 12986 19472 13466
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19444 12442 19472 12922
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19892 11824 19944 11830
rect 19892 11766 19944 11772
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19444 10810 19472 11698
rect 19904 11218 19932 11766
rect 19996 11218 20024 14418
rect 20088 14414 20116 14894
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 13938 20116 14214
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20088 12850 20116 13874
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 20180 11150 20208 15030
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 20168 10192 20220 10198
rect 20168 10134 20220 10140
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 20180 9654 20208 10134
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20180 9178 20208 9590
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19444 6458 19472 6734
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19260 6322 19288 6394
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19996 5914 20024 7346
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 20272 5710 20300 18022
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20364 13870 20392 15846
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 9042 20392 12582
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20272 5370 20300 5646
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18984 4282 19012 4694
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18892 3738 18920 4082
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18984 3058 19012 4218
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19352 3058 19380 3878
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18236 2576 18288 2582
rect 18236 2518 18288 2524
rect 18892 2514 18920 2790
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18892 800 18920 2450
rect 19444 2446 19472 5306
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19812 3602 19840 4014
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20088 3058 20116 4422
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20364 3670 20392 3878
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 20260 3460 20312 3466
rect 20456 3448 20484 17818
rect 20548 14482 20576 18158
rect 20640 15910 20668 19110
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14822 20668 14894
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20640 12782 20668 14758
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20732 14074 20760 14350
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22112 13734 22140 13806
rect 22652 13796 22704 13802
rect 22652 13738 22704 13744
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20732 11150 20760 11494
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20640 10554 20668 11086
rect 20732 11014 20760 11086
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20640 10526 20760 10554
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20640 6866 20668 10202
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20640 6254 20668 6802
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20732 5250 20760 10526
rect 20824 9654 20852 11018
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20916 10674 20944 10950
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20824 8974 20852 9590
rect 21100 9518 21128 11154
rect 22112 11082 22140 13670
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21008 8294 21036 8774
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 21100 7002 21128 9454
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22204 8498 22232 8774
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22020 7954 22048 8230
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22296 7410 22324 7822
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 22296 6866 22324 7346
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22112 5778 22140 6666
rect 22204 6118 22232 6734
rect 22296 6662 22324 6802
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 20732 5222 20852 5250
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20312 3420 20484 3448
rect 20260 3402 20312 3408
rect 20456 3058 20484 3420
rect 20640 3058 20668 4082
rect 20732 3942 20760 5034
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20732 3398 20760 3606
rect 20824 3534 20852 5222
rect 22112 4622 22140 5714
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20088 2774 20116 2994
rect 19996 2746 20116 2774
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2746
rect 20640 1970 20668 2994
rect 21100 2666 21128 3402
rect 21376 3126 21404 3606
rect 22112 3602 22140 4558
rect 22204 4146 22232 6054
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22112 3398 22140 3538
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 22296 3040 22324 6598
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22388 4146 22416 4422
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22480 3534 22508 8842
rect 22572 7954 22600 11018
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22664 4486 22692 13738
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22756 8838 22784 8978
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22756 7478 22784 8774
rect 22836 7812 22888 7818
rect 22836 7754 22888 7760
rect 22744 7472 22796 7478
rect 22744 7414 22796 7420
rect 22848 7410 22876 7754
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22848 6914 22876 7346
rect 22848 6886 22968 6914
rect 22940 6798 22968 6886
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22376 3052 22428 3058
rect 22296 3012 22376 3040
rect 22376 2994 22428 3000
rect 21008 2638 21128 2666
rect 21008 2446 21036 2638
rect 21088 2508 21140 2514
rect 21088 2450 21140 2456
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 20628 1964 20680 1970
rect 20628 1906 20680 1912
rect 21100 800 21128 2450
rect 22192 2372 22244 2378
rect 22192 2314 22244 2320
rect 22204 800 22232 2314
rect 22388 2106 22416 2994
rect 22480 2650 22508 3470
rect 22572 3194 22600 3470
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22664 2514 22692 4422
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22756 3738 22784 4082
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 23952 3194 23980 55830
rect 25056 55826 25084 57258
rect 25872 57248 25924 57254
rect 25872 57190 25924 57196
rect 26148 57248 26200 57254
rect 26148 57190 26200 57196
rect 25320 56432 25372 56438
rect 25320 56374 25372 56380
rect 25778 56400 25834 56409
rect 25228 56364 25280 56370
rect 25228 56306 25280 56312
rect 25136 56160 25188 56166
rect 25136 56102 25188 56108
rect 25044 55820 25096 55826
rect 25044 55762 25096 55768
rect 25148 55758 25176 56102
rect 25240 55894 25268 56306
rect 25332 56166 25360 56374
rect 25778 56335 25780 56344
rect 25832 56335 25834 56344
rect 25780 56306 25832 56312
rect 25320 56160 25372 56166
rect 25320 56102 25372 56108
rect 25792 55894 25820 56306
rect 25228 55888 25280 55894
rect 25228 55830 25280 55836
rect 25412 55888 25464 55894
rect 25412 55830 25464 55836
rect 25780 55888 25832 55894
rect 25780 55830 25832 55836
rect 24676 55752 24728 55758
rect 24676 55694 24728 55700
rect 25136 55752 25188 55758
rect 25136 55694 25188 55700
rect 24400 54528 24452 54534
rect 24400 54470 24452 54476
rect 24412 54194 24440 54470
rect 24400 54188 24452 54194
rect 24400 54130 24452 54136
rect 24688 54126 24716 55694
rect 25240 55622 25268 55830
rect 25228 55616 25280 55622
rect 25228 55558 25280 55564
rect 25424 54194 25452 55830
rect 25780 55752 25832 55758
rect 25780 55694 25832 55700
rect 25792 55418 25820 55694
rect 25780 55412 25832 55418
rect 25780 55354 25832 55360
rect 25792 54874 25820 55354
rect 25780 54868 25832 54874
rect 25780 54810 25832 54816
rect 25792 54754 25820 54810
rect 25700 54726 25820 54754
rect 25700 54194 25728 54726
rect 25884 54194 25912 57190
rect 25964 55616 26016 55622
rect 25964 55558 26016 55564
rect 25976 54670 26004 55558
rect 26056 55276 26108 55282
rect 26056 55218 26108 55224
rect 25964 54664 26016 54670
rect 25964 54606 26016 54612
rect 25976 54262 26004 54606
rect 25964 54256 26016 54262
rect 25964 54198 26016 54204
rect 26068 54194 26096 55218
rect 26160 54670 26188 57190
rect 28184 57050 28212 57394
rect 30380 57384 30432 57390
rect 30380 57326 30432 57332
rect 28356 57248 28408 57254
rect 28356 57190 28408 57196
rect 29736 57248 29788 57254
rect 29736 57190 29788 57196
rect 28172 57044 28224 57050
rect 28172 56986 28224 56992
rect 26240 56908 26292 56914
rect 26240 56850 26292 56856
rect 26148 54664 26200 54670
rect 26148 54606 26200 54612
rect 26252 54602 26280 56850
rect 27436 56500 27488 56506
rect 27436 56442 27488 56448
rect 27448 56409 27476 56442
rect 26422 56400 26478 56409
rect 26422 56335 26424 56344
rect 26476 56335 26478 56344
rect 27434 56400 27490 56409
rect 27434 56335 27490 56344
rect 27528 56364 27580 56370
rect 26424 56306 26476 56312
rect 26884 56296 26936 56302
rect 26884 56238 26936 56244
rect 27344 56296 27396 56302
rect 27344 56238 27396 56244
rect 26896 56001 26924 56238
rect 26882 55992 26938 56001
rect 26882 55927 26938 55936
rect 26608 55888 26660 55894
rect 26608 55830 26660 55836
rect 26620 55282 26648 55830
rect 27356 55758 27384 56238
rect 26976 55752 27028 55758
rect 26974 55720 26976 55729
rect 27344 55752 27396 55758
rect 27028 55720 27030 55729
rect 27344 55694 27396 55700
rect 26974 55655 27030 55664
rect 26608 55276 26660 55282
rect 26608 55218 26660 55224
rect 26620 54670 26648 55218
rect 26608 54664 26660 54670
rect 26608 54606 26660 54612
rect 27448 54602 27476 56335
rect 27528 56306 27580 56312
rect 27540 55593 27568 56306
rect 28368 55826 28396 57190
rect 29184 56976 29236 56982
rect 29184 56918 29236 56924
rect 28998 56400 29054 56409
rect 28954 56370 28998 56376
rect 28816 56364 28868 56370
rect 29006 56335 29054 56344
rect 29006 56324 29040 56335
rect 28954 56312 29006 56318
rect 28816 56306 28868 56312
rect 28540 56296 28592 56302
rect 28540 56238 28592 56244
rect 28630 56264 28686 56273
rect 28356 55820 28408 55826
rect 28356 55762 28408 55768
rect 28448 55752 28500 55758
rect 28354 55720 28410 55729
rect 28448 55694 28500 55700
rect 28354 55655 28356 55664
rect 28408 55655 28410 55664
rect 28356 55626 28408 55632
rect 27526 55584 27582 55593
rect 27526 55519 27582 55528
rect 26240 54596 26292 54602
rect 26240 54538 26292 54544
rect 27436 54596 27488 54602
rect 27436 54538 27488 54544
rect 27344 54528 27396 54534
rect 27344 54470 27396 54476
rect 27356 54262 27384 54470
rect 27344 54256 27396 54262
rect 27344 54198 27396 54204
rect 27540 54194 27568 55519
rect 28460 55418 28488 55694
rect 28448 55412 28500 55418
rect 28448 55354 28500 55360
rect 28552 55282 28580 56238
rect 28630 56199 28632 56208
rect 28684 56199 28686 56208
rect 28632 56170 28684 56176
rect 28724 56160 28776 56166
rect 28724 56102 28776 56108
rect 28540 55276 28592 55282
rect 28540 55218 28592 55224
rect 25412 54188 25464 54194
rect 25412 54130 25464 54136
rect 25688 54188 25740 54194
rect 25688 54130 25740 54136
rect 25872 54188 25924 54194
rect 25872 54130 25924 54136
rect 26056 54188 26108 54194
rect 26056 54130 26108 54136
rect 27528 54188 27580 54194
rect 27528 54130 27580 54136
rect 24676 54120 24728 54126
rect 24676 54062 24728 54068
rect 24688 53650 24716 54062
rect 24768 53984 24820 53990
rect 24768 53926 24820 53932
rect 24676 53644 24728 53650
rect 24676 53586 24728 53592
rect 24780 53582 24808 53926
rect 24768 53576 24820 53582
rect 24768 53518 24820 53524
rect 28736 3194 28764 56102
rect 28828 55962 28856 56306
rect 28906 55992 28962 56001
rect 28816 55956 28868 55962
rect 28906 55927 28908 55936
rect 28816 55898 28868 55904
rect 28960 55927 28962 55936
rect 28908 55898 28960 55904
rect 29196 55758 29224 56918
rect 29748 56914 29776 57190
rect 29736 56908 29788 56914
rect 29736 56850 29788 56856
rect 29368 56840 29420 56846
rect 29368 56782 29420 56788
rect 29828 56840 29880 56846
rect 29828 56782 29880 56788
rect 29380 56438 29408 56782
rect 29460 56772 29512 56778
rect 29460 56714 29512 56720
rect 29368 56432 29420 56438
rect 29368 56374 29420 56380
rect 29184 55752 29236 55758
rect 29184 55694 29236 55700
rect 29472 55690 29500 56714
rect 29460 55684 29512 55690
rect 29460 55626 29512 55632
rect 28816 55616 28868 55622
rect 28814 55584 28816 55593
rect 28868 55584 28870 55593
rect 28814 55519 28870 55528
rect 29000 55412 29052 55418
rect 29000 55354 29052 55360
rect 29012 53242 29040 55354
rect 29472 53990 29500 55626
rect 29840 55418 29868 56782
rect 30196 56704 30248 56710
rect 30196 56646 30248 56652
rect 30208 56370 30236 56646
rect 30392 56370 30420 57326
rect 32140 57050 32168 57394
rect 32312 57248 32364 57254
rect 32312 57190 32364 57196
rect 32956 57248 33008 57254
rect 32956 57190 33008 57196
rect 33232 57248 33284 57254
rect 33232 57190 33284 57196
rect 34704 57248 34756 57254
rect 34704 57190 34756 57196
rect 32128 57044 32180 57050
rect 32128 56986 32180 56992
rect 30472 56500 30524 56506
rect 30472 56442 30524 56448
rect 31392 56500 31444 56506
rect 31392 56442 31444 56448
rect 30484 56370 30512 56442
rect 31024 56432 31076 56438
rect 31024 56374 31076 56380
rect 30196 56364 30248 56370
rect 30196 56306 30248 56312
rect 30380 56364 30432 56370
rect 30380 56306 30432 56312
rect 30472 56364 30524 56370
rect 30472 56306 30524 56312
rect 30656 56364 30708 56370
rect 30656 56306 30708 56312
rect 29920 56160 29972 56166
rect 29920 56102 29972 56108
rect 29932 55758 29960 56102
rect 30288 55888 30340 55894
rect 30288 55830 30340 55836
rect 29920 55752 29972 55758
rect 29920 55694 29972 55700
rect 30012 55684 30064 55690
rect 30012 55626 30064 55632
rect 29828 55412 29880 55418
rect 29828 55354 29880 55360
rect 30024 55350 30052 55626
rect 30012 55344 30064 55350
rect 30012 55286 30064 55292
rect 29736 54120 29788 54126
rect 29736 54062 29788 54068
rect 29460 53984 29512 53990
rect 29460 53926 29512 53932
rect 29748 53582 29776 54062
rect 29920 53984 29972 53990
rect 29920 53926 29972 53932
rect 29828 53712 29880 53718
rect 29828 53654 29880 53660
rect 29736 53576 29788 53582
rect 29736 53518 29788 53524
rect 29000 53236 29052 53242
rect 29000 53178 29052 53184
rect 29748 53038 29776 53518
rect 29736 53032 29788 53038
rect 29736 52974 29788 52980
rect 28816 52896 28868 52902
rect 28816 52838 28868 52844
rect 28828 16574 28856 52838
rect 29748 52698 29776 52974
rect 29736 52692 29788 52698
rect 29736 52634 29788 52640
rect 28828 16546 28948 16574
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 23308 2446 23336 2790
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 23308 800 23336 2382
rect 24412 2378 24440 2790
rect 25516 2446 25544 2790
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 24400 2372 24452 2378
rect 24400 2314 24452 2320
rect 24412 800 24440 2314
rect 25516 800 25544 2382
rect 26608 2304 26660 2310
rect 26608 2246 26660 2252
rect 26620 800 26648 2246
rect 27724 800 27752 2790
rect 28736 2446 28764 3130
rect 28920 2650 28948 16546
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 29748 2514 29776 52634
rect 29840 3194 29868 53654
rect 29932 53582 29960 53926
rect 29920 53576 29972 53582
rect 29920 53518 29972 53524
rect 29932 53106 29960 53518
rect 29920 53100 29972 53106
rect 29920 53042 29972 53048
rect 29828 3188 29880 3194
rect 29828 3130 29880 3136
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 29840 2446 29868 3130
rect 30300 3126 30328 55830
rect 30484 53718 30512 56306
rect 30668 55729 30696 56306
rect 30840 56296 30892 56302
rect 30840 56238 30892 56244
rect 30654 55720 30710 55729
rect 30654 55655 30710 55664
rect 30564 54188 30616 54194
rect 30564 54130 30616 54136
rect 30472 53712 30524 53718
rect 30472 53654 30524 53660
rect 30576 53582 30604 54130
rect 30852 53786 30880 56238
rect 31036 55894 31064 56374
rect 31208 56364 31260 56370
rect 31208 56306 31260 56312
rect 31024 55888 31076 55894
rect 31024 55830 31076 55836
rect 31220 55826 31248 56306
rect 31208 55820 31260 55826
rect 31208 55762 31260 55768
rect 31404 54738 31432 56442
rect 32324 56438 32352 57190
rect 32312 56432 32364 56438
rect 32312 56374 32364 56380
rect 31668 56364 31720 56370
rect 32772 56364 32824 56370
rect 31720 56324 31800 56352
rect 31668 56306 31720 56312
rect 31772 55690 31800 56324
rect 32824 56324 32904 56352
rect 32772 56306 32824 56312
rect 32586 56264 32642 56273
rect 32586 56199 32642 56208
rect 32600 56166 32628 56199
rect 32588 56160 32640 56166
rect 32588 56102 32640 56108
rect 32876 55758 32904 56324
rect 32968 55758 32996 57190
rect 33048 56364 33100 56370
rect 33048 56306 33100 56312
rect 33060 56166 33088 56306
rect 33140 56228 33192 56234
rect 33140 56170 33192 56176
rect 33048 56160 33100 56166
rect 33048 56102 33100 56108
rect 32864 55752 32916 55758
rect 32864 55694 32916 55700
rect 32956 55752 33008 55758
rect 32956 55694 33008 55700
rect 31760 55684 31812 55690
rect 31760 55626 31812 55632
rect 31392 54732 31444 54738
rect 31392 54674 31444 54680
rect 30932 54324 30984 54330
rect 30932 54266 30984 54272
rect 30840 53780 30892 53786
rect 30840 53722 30892 53728
rect 30564 53576 30616 53582
rect 30564 53518 30616 53524
rect 30944 3194 30972 54266
rect 31772 53786 31800 55626
rect 32404 55072 32456 55078
rect 32404 55014 32456 55020
rect 32416 54670 32444 55014
rect 32876 54874 32904 55694
rect 32864 54868 32916 54874
rect 32864 54810 32916 54816
rect 32496 54800 32548 54806
rect 32496 54742 32548 54748
rect 32404 54664 32456 54670
rect 32404 54606 32456 54612
rect 31852 54528 31904 54534
rect 31852 54470 31904 54476
rect 31864 54330 31892 54470
rect 31852 54324 31904 54330
rect 31852 54266 31904 54272
rect 31864 54126 31892 54266
rect 32312 54256 32364 54262
rect 32312 54198 32364 54204
rect 32324 54126 32352 54198
rect 32416 54126 32444 54606
rect 32508 54330 32536 54742
rect 32772 54528 32824 54534
rect 32772 54470 32824 54476
rect 32496 54324 32548 54330
rect 32496 54266 32548 54272
rect 32588 54256 32640 54262
rect 32588 54198 32640 54204
rect 31852 54120 31904 54126
rect 31852 54062 31904 54068
rect 32312 54120 32364 54126
rect 32312 54062 32364 54068
rect 32404 54120 32456 54126
rect 32404 54062 32456 54068
rect 32312 53984 32364 53990
rect 32312 53926 32364 53932
rect 31760 53780 31812 53786
rect 31760 53722 31812 53728
rect 32324 53582 32352 53926
rect 32312 53576 32364 53582
rect 32312 53518 32364 53524
rect 32324 53106 32352 53518
rect 32416 53174 32444 54062
rect 32600 53718 32628 54198
rect 32680 54188 32732 54194
rect 32680 54130 32732 54136
rect 32588 53712 32640 53718
rect 32588 53654 32640 53660
rect 32600 53582 32628 53654
rect 32692 53582 32720 54130
rect 32784 53650 32812 54470
rect 32772 53644 32824 53650
rect 32772 53586 32824 53592
rect 32588 53576 32640 53582
rect 32588 53518 32640 53524
rect 32680 53576 32732 53582
rect 32680 53518 32732 53524
rect 32600 53446 32628 53518
rect 32588 53440 32640 53446
rect 32588 53382 32640 53388
rect 32784 53242 32812 53586
rect 32772 53236 32824 53242
rect 32772 53178 32824 53184
rect 32404 53168 32456 53174
rect 32404 53110 32456 53116
rect 32312 53100 32364 53106
rect 32312 53042 32364 53048
rect 33152 3194 33180 56170
rect 33244 54602 33272 57190
rect 34716 56438 34744 57190
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 35360 57050 35388 57394
rect 36452 57316 36504 57322
rect 36452 57258 36504 57264
rect 35808 57248 35860 57254
rect 35808 57190 35860 57196
rect 35900 57248 35952 57254
rect 35900 57190 35952 57196
rect 35348 57044 35400 57050
rect 35348 56986 35400 56992
rect 34980 56500 35032 56506
rect 34980 56442 35032 56448
rect 34520 56432 34572 56438
rect 34520 56374 34572 56380
rect 34704 56432 34756 56438
rect 34704 56374 34756 56380
rect 33324 56364 33376 56370
rect 33324 56306 33376 56312
rect 33336 56234 33364 56306
rect 33324 56228 33376 56234
rect 33324 56170 33376 56176
rect 33336 55758 33364 56170
rect 33324 55752 33376 55758
rect 33324 55694 33376 55700
rect 34532 55418 34560 56374
rect 34992 56370 35020 56442
rect 35820 56438 35848 57190
rect 35808 56432 35860 56438
rect 35162 56400 35218 56409
rect 34612 56364 34664 56370
rect 34612 56306 34664 56312
rect 34980 56364 35032 56370
rect 34980 56306 35032 56312
rect 35072 56364 35124 56370
rect 35162 56335 35218 56344
rect 35530 56400 35586 56409
rect 35808 56374 35860 56380
rect 35530 56335 35532 56344
rect 35072 56306 35124 56312
rect 34624 55758 34652 56306
rect 35084 56234 35112 56306
rect 35176 56234 35204 56335
rect 35584 56335 35586 56344
rect 35716 56364 35768 56370
rect 35532 56306 35584 56312
rect 35716 56306 35768 56312
rect 35072 56228 35124 56234
rect 35072 56170 35124 56176
rect 35164 56228 35216 56234
rect 35164 56170 35216 56176
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34612 55752 34664 55758
rect 34612 55694 34664 55700
rect 34520 55412 34572 55418
rect 34520 55354 34572 55360
rect 34624 54874 34652 55694
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34612 54868 34664 54874
rect 34612 54810 34664 54816
rect 34624 54670 34652 54810
rect 35544 54754 35572 56306
rect 35624 56228 35676 56234
rect 35624 56170 35676 56176
rect 35636 55690 35664 56170
rect 35728 55758 35756 56306
rect 35912 55758 35940 57190
rect 35992 56704 36044 56710
rect 35992 56646 36044 56652
rect 36004 56506 36032 56646
rect 35992 56500 36044 56506
rect 35992 56442 36044 56448
rect 36174 56400 36230 56409
rect 36084 56364 36136 56370
rect 36230 56344 36308 56352
rect 36174 56335 36176 56344
rect 36084 56306 36136 56312
rect 36228 56324 36308 56344
rect 36176 56306 36228 56312
rect 36096 55962 36124 56306
rect 36084 55956 36136 55962
rect 36084 55898 36136 55904
rect 36280 55758 36308 56324
rect 35716 55752 35768 55758
rect 35716 55694 35768 55700
rect 35900 55752 35952 55758
rect 35900 55694 35952 55700
rect 36268 55752 36320 55758
rect 36268 55694 36320 55700
rect 35624 55684 35676 55690
rect 35624 55626 35676 55632
rect 35624 55208 35676 55214
rect 35624 55150 35676 55156
rect 34704 54732 34756 54738
rect 34704 54674 34756 54680
rect 35360 54726 35572 54754
rect 34612 54664 34664 54670
rect 34612 54606 34664 54612
rect 33232 54596 33284 54602
rect 33232 54538 33284 54544
rect 34716 54194 34744 54674
rect 34888 54528 34940 54534
rect 34888 54470 34940 54476
rect 34704 54188 34756 54194
rect 34704 54130 34756 54136
rect 34900 54058 34928 54470
rect 35360 54330 35388 54726
rect 35544 54670 35572 54726
rect 35440 54664 35492 54670
rect 35440 54606 35492 54612
rect 35532 54664 35584 54670
rect 35532 54606 35584 54612
rect 35452 54330 35480 54606
rect 35636 54602 35664 55150
rect 35624 54596 35676 54602
rect 35624 54538 35676 54544
rect 35348 54324 35400 54330
rect 35348 54266 35400 54272
rect 35440 54324 35492 54330
rect 35440 54266 35492 54272
rect 35348 54188 35400 54194
rect 35348 54130 35400 54136
rect 34888 54052 34940 54058
rect 34888 53994 34940 54000
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 35360 53514 35388 54130
rect 36464 54058 36492 57258
rect 36556 57050 36584 57394
rect 38384 57384 38436 57390
rect 38384 57326 38436 57332
rect 37648 57248 37700 57254
rect 37648 57190 37700 57196
rect 36544 57044 36596 57050
rect 36544 56986 36596 56992
rect 37660 56370 37688 57190
rect 37832 56976 37884 56982
rect 37832 56918 37884 56924
rect 37844 56438 37872 56918
rect 38016 56500 38068 56506
rect 38016 56442 38068 56448
rect 37832 56432 37884 56438
rect 37832 56374 37884 56380
rect 38028 56370 38056 56442
rect 37648 56364 37700 56370
rect 37648 56306 37700 56312
rect 37740 56364 37792 56370
rect 37740 56306 37792 56312
rect 38016 56364 38068 56370
rect 38016 56306 38068 56312
rect 37556 56160 37608 56166
rect 37556 56102 37608 56108
rect 37568 55894 37596 56102
rect 37556 55888 37608 55894
rect 37556 55830 37608 55836
rect 37752 55758 37780 56306
rect 38292 55888 38344 55894
rect 38292 55830 38344 55836
rect 37740 55752 37792 55758
rect 37740 55694 37792 55700
rect 37464 55684 37516 55690
rect 37464 55626 37516 55632
rect 37476 54874 37504 55626
rect 38304 55418 38332 55830
rect 38292 55412 38344 55418
rect 38292 55354 38344 55360
rect 37464 54868 37516 54874
rect 37464 54810 37516 54816
rect 38396 54738 38424 57326
rect 38660 57248 38712 57254
rect 38660 57190 38712 57196
rect 38672 56370 38700 57190
rect 38764 56846 38792 57530
rect 38844 57520 38896 57526
rect 38844 57462 38896 57468
rect 38752 56840 38804 56846
rect 38752 56782 38804 56788
rect 38752 56704 38804 56710
rect 38752 56646 38804 56652
rect 38764 56370 38792 56646
rect 38660 56364 38712 56370
rect 38660 56306 38712 56312
rect 38752 56364 38804 56370
rect 38752 56306 38804 56312
rect 38660 56160 38712 56166
rect 38660 56102 38712 56108
rect 38672 55978 38700 56102
rect 38626 55962 38700 55978
rect 38614 55956 38700 55962
rect 38666 55950 38700 55956
rect 38614 55898 38666 55904
rect 38764 55865 38792 56306
rect 38750 55856 38806 55865
rect 38672 55800 38750 55808
rect 38856 55826 38884 57462
rect 38948 57458 38976 59200
rect 40144 57458 40172 59200
rect 41340 57458 41368 59200
rect 42536 57882 42564 59200
rect 42536 57854 42840 57882
rect 42708 57588 42760 57594
rect 42708 57530 42760 57536
rect 38936 57452 38988 57458
rect 38936 57394 38988 57400
rect 40132 57452 40184 57458
rect 40132 57394 40184 57400
rect 41328 57452 41380 57458
rect 41328 57394 41380 57400
rect 38948 57050 38976 57394
rect 41340 57050 41368 57394
rect 38936 57044 38988 57050
rect 38936 56986 38988 56992
rect 41328 57044 41380 57050
rect 41328 56986 41380 56992
rect 39120 56840 39172 56846
rect 39028 56818 39080 56824
rect 38948 56766 39028 56794
rect 39120 56782 39172 56788
rect 38948 56370 38976 56766
rect 39028 56760 39080 56766
rect 39132 56692 39160 56782
rect 39040 56664 39160 56692
rect 39040 56370 39068 56664
rect 42720 56438 42748 57530
rect 42812 57458 42840 57854
rect 43732 57458 43760 59200
rect 44928 57458 44956 59200
rect 46124 57458 46152 59200
rect 47320 57458 47348 59200
rect 48516 57458 48544 59200
rect 49712 57458 49740 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50908 57474 50936 59200
rect 50908 57458 51120 57474
rect 52104 57458 52132 59200
rect 53300 57458 53328 59200
rect 54496 57458 54524 59200
rect 55692 57458 55720 59200
rect 56888 57458 56916 59200
rect 57518 58984 57574 58993
rect 57518 58919 57574 58928
rect 42800 57452 42852 57458
rect 42800 57394 42852 57400
rect 43720 57452 43772 57458
rect 43720 57394 43772 57400
rect 44916 57452 44968 57458
rect 44916 57394 44968 57400
rect 46112 57452 46164 57458
rect 46112 57394 46164 57400
rect 47308 57452 47360 57458
rect 47308 57394 47360 57400
rect 48504 57452 48556 57458
rect 48504 57394 48556 57400
rect 49700 57452 49752 57458
rect 49700 57394 49752 57400
rect 50344 57452 50396 57458
rect 50908 57452 51132 57458
rect 50908 57446 51080 57452
rect 50344 57394 50396 57400
rect 51080 57394 51132 57400
rect 52092 57452 52144 57458
rect 52092 57394 52144 57400
rect 53288 57452 53340 57458
rect 53288 57394 53340 57400
rect 54484 57452 54536 57458
rect 54484 57394 54536 57400
rect 55680 57452 55732 57458
rect 55680 57394 55732 57400
rect 56876 57452 56928 57458
rect 56876 57394 56928 57400
rect 44548 57384 44600 57390
rect 44548 57326 44600 57332
rect 42800 57316 42852 57322
rect 42800 57258 42852 57264
rect 42708 56432 42760 56438
rect 42708 56374 42760 56380
rect 38936 56364 38988 56370
rect 38936 56306 38988 56312
rect 39028 56364 39080 56370
rect 39028 56306 39080 56312
rect 40776 56364 40828 56370
rect 40960 56364 41012 56370
rect 40828 56324 40908 56352
rect 40776 56306 40828 56312
rect 38672 55791 38806 55800
rect 38844 55820 38896 55826
rect 38672 55780 38792 55791
rect 38476 55752 38528 55758
rect 38672 55740 38700 55780
rect 38844 55762 38896 55768
rect 38528 55712 38700 55740
rect 38752 55730 38804 55736
rect 38750 55720 38752 55729
rect 38804 55720 38806 55729
rect 38476 55694 38528 55700
rect 37556 54732 37608 54738
rect 37556 54674 37608 54680
rect 38384 54732 38436 54738
rect 38384 54674 38436 54680
rect 37568 54602 37596 54674
rect 37924 54664 37976 54670
rect 37924 54606 37976 54612
rect 38016 54664 38068 54670
rect 38016 54606 38068 54612
rect 37556 54596 37608 54602
rect 37556 54538 37608 54544
rect 36544 54188 36596 54194
rect 36544 54130 36596 54136
rect 36820 54188 36872 54194
rect 36820 54130 36872 54136
rect 36452 54052 36504 54058
rect 36452 53994 36504 54000
rect 36556 53718 36584 54130
rect 36832 53990 36860 54130
rect 36820 53984 36872 53990
rect 36820 53926 36872 53932
rect 37568 53786 37596 54538
rect 37936 54534 37964 54606
rect 37924 54528 37976 54534
rect 37924 54470 37976 54476
rect 37936 54262 37964 54470
rect 38028 54330 38056 54606
rect 38016 54324 38068 54330
rect 38016 54266 38068 54272
rect 37924 54256 37976 54262
rect 37924 54198 37976 54204
rect 38488 53786 38516 55694
rect 38750 55655 38806 55664
rect 38844 55684 38896 55690
rect 38948 55672 38976 56306
rect 39040 55690 39068 56306
rect 40500 56296 40552 56302
rect 40500 56238 40552 56244
rect 40512 55758 40540 56238
rect 40500 55752 40552 55758
rect 40500 55694 40552 55700
rect 40880 55740 40908 56324
rect 40960 56306 41012 56312
rect 41236 56364 41288 56370
rect 41236 56306 41288 56312
rect 42616 56364 42668 56370
rect 42616 56306 42668 56312
rect 40972 55962 41000 56306
rect 41144 56160 41196 56166
rect 41144 56102 41196 56108
rect 40960 55956 41012 55962
rect 40960 55898 41012 55904
rect 41156 55894 41184 56102
rect 41144 55888 41196 55894
rect 41144 55830 41196 55836
rect 41052 55752 41104 55758
rect 40880 55712 41052 55740
rect 38896 55644 38976 55672
rect 38844 55626 38896 55632
rect 38752 55276 38804 55282
rect 38752 55218 38804 55224
rect 38660 54664 38712 54670
rect 38764 54618 38792 55218
rect 38712 54612 38792 54618
rect 38660 54606 38792 54612
rect 38672 54590 38792 54606
rect 38672 54262 38700 54590
rect 38948 54534 38976 55644
rect 39028 55684 39080 55690
rect 39028 55626 39080 55632
rect 38936 54528 38988 54534
rect 38936 54470 38988 54476
rect 39040 54330 39068 55626
rect 40316 55344 40368 55350
rect 40316 55286 40368 55292
rect 39580 55276 39632 55282
rect 39580 55218 39632 55224
rect 39592 54602 39620 55218
rect 39580 54596 39632 54602
rect 39580 54538 39632 54544
rect 39028 54324 39080 54330
rect 39028 54266 39080 54272
rect 38660 54256 38712 54262
rect 38660 54198 38712 54204
rect 37556 53780 37608 53786
rect 37556 53722 37608 53728
rect 38476 53780 38528 53786
rect 38476 53722 38528 53728
rect 36544 53712 36596 53718
rect 36544 53654 36596 53660
rect 37568 53514 37596 53722
rect 38672 53582 38700 54198
rect 39592 54126 39620 54538
rect 39672 54528 39724 54534
rect 39672 54470 39724 54476
rect 39684 54194 39712 54470
rect 40328 54330 40356 55286
rect 40880 55282 40908 55712
rect 41052 55694 41104 55700
rect 41248 55350 41276 56306
rect 41512 55956 41564 55962
rect 41512 55898 41564 55904
rect 41524 55690 41552 55898
rect 42628 55758 42656 56306
rect 41788 55752 41840 55758
rect 41788 55694 41840 55700
rect 42616 55752 42668 55758
rect 42616 55694 42668 55700
rect 41512 55684 41564 55690
rect 41512 55626 41564 55632
rect 41236 55344 41288 55350
rect 41236 55286 41288 55292
rect 40868 55276 40920 55282
rect 40868 55218 40920 55224
rect 40880 54330 40908 55218
rect 41524 55214 41552 55626
rect 41800 55350 41828 55694
rect 41788 55344 41840 55350
rect 41788 55286 41840 55292
rect 42628 55282 42656 55694
rect 42812 55690 42840 57258
rect 43352 56840 43404 56846
rect 43352 56782 43404 56788
rect 43904 56840 43956 56846
rect 43904 56782 43956 56788
rect 42984 56432 43036 56438
rect 42984 56374 43036 56380
rect 42800 55684 42852 55690
rect 42800 55626 42852 55632
rect 42996 55282 43024 56374
rect 43364 56370 43392 56782
rect 43628 56772 43680 56778
rect 43628 56714 43680 56720
rect 43640 56438 43668 56714
rect 43628 56432 43680 56438
rect 43628 56374 43680 56380
rect 43352 56364 43404 56370
rect 43352 56306 43404 56312
rect 43168 56160 43220 56166
rect 43168 56102 43220 56108
rect 43180 55622 43208 56102
rect 43640 55758 43668 56374
rect 43916 56370 43944 56782
rect 43904 56364 43956 56370
rect 43904 56306 43956 56312
rect 43916 55758 43944 56306
rect 43628 55752 43680 55758
rect 43628 55694 43680 55700
rect 43904 55752 43956 55758
rect 43904 55694 43956 55700
rect 43168 55616 43220 55622
rect 43168 55558 43220 55564
rect 43916 55418 43944 55694
rect 43352 55412 43404 55418
rect 43352 55354 43404 55360
rect 43904 55412 43956 55418
rect 43904 55354 43956 55360
rect 43364 55282 43392 55354
rect 44560 55282 44588 57326
rect 44640 57316 44692 57322
rect 44640 57258 44692 57264
rect 44652 56506 44680 57258
rect 44928 57050 44956 57394
rect 47320 57050 47348 57394
rect 48596 57248 48648 57254
rect 48596 57190 48648 57196
rect 48688 57248 48740 57254
rect 48688 57190 48740 57196
rect 44916 57044 44968 57050
rect 44916 56986 44968 56992
rect 47308 57044 47360 57050
rect 47308 56986 47360 56992
rect 48608 56982 48636 57190
rect 44732 56976 44784 56982
rect 44732 56918 44784 56924
rect 48596 56976 48648 56982
rect 48596 56918 48648 56924
rect 44640 56500 44692 56506
rect 44640 56442 44692 56448
rect 44744 55690 44772 56918
rect 48700 56914 48728 57190
rect 50356 57050 50384 57394
rect 52104 57050 52132 57394
rect 52184 57248 52236 57254
rect 52184 57190 52236 57196
rect 53380 57248 53432 57254
rect 53380 57190 53432 57196
rect 50344 57044 50396 57050
rect 50344 56986 50396 56992
rect 52092 57044 52144 57050
rect 52092 56986 52144 56992
rect 48688 56908 48740 56914
rect 48688 56850 48740 56856
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 52196 55826 52224 57190
rect 53392 56234 53420 57190
rect 54496 57050 54524 57394
rect 54576 57248 54628 57254
rect 54576 57190 54628 57196
rect 55772 57248 55824 57254
rect 55772 57190 55824 57196
rect 54484 57044 54536 57050
rect 54484 56986 54536 56992
rect 53380 56228 53432 56234
rect 53380 56170 53432 56176
rect 52184 55820 52236 55826
rect 52184 55762 52236 55768
rect 44732 55684 44784 55690
rect 44732 55626 44784 55632
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 54588 55350 54616 57190
rect 55784 55690 55812 57190
rect 56888 57050 56916 57394
rect 57058 57352 57114 57361
rect 57058 57287 57114 57296
rect 56968 57248 57020 57254
rect 56968 57190 57020 57196
rect 56876 57044 56928 57050
rect 56876 56986 56928 56992
rect 56980 56778 57008 57190
rect 57072 56846 57100 57287
rect 57532 56846 57560 58919
rect 58084 57458 58112 59200
rect 58438 58168 58494 58177
rect 58438 58103 58494 58112
rect 58072 57452 58124 57458
rect 58072 57394 58124 57400
rect 57060 56840 57112 56846
rect 57060 56782 57112 56788
rect 57520 56840 57572 56846
rect 57520 56782 57572 56788
rect 56968 56772 57020 56778
rect 56968 56714 57020 56720
rect 56876 56704 56928 56710
rect 56876 56646 56928 56652
rect 55772 55684 55824 55690
rect 55772 55626 55824 55632
rect 56692 55412 56744 55418
rect 56692 55354 56744 55360
rect 54576 55344 54628 55350
rect 54576 55286 54628 55292
rect 42616 55276 42668 55282
rect 42616 55218 42668 55224
rect 42984 55276 43036 55282
rect 42984 55218 43036 55224
rect 43352 55276 43404 55282
rect 43352 55218 43404 55224
rect 44548 55276 44600 55282
rect 44548 55218 44600 55224
rect 41512 55208 41564 55214
rect 41512 55150 41564 55156
rect 40316 54324 40368 54330
rect 40316 54266 40368 54272
rect 40868 54324 40920 54330
rect 40868 54266 40920 54272
rect 39672 54188 39724 54194
rect 39672 54130 39724 54136
rect 39580 54120 39632 54126
rect 39580 54062 39632 54068
rect 39592 53990 39620 54062
rect 39684 54058 39712 54130
rect 39672 54052 39724 54058
rect 39672 53994 39724 54000
rect 39580 53984 39632 53990
rect 39580 53926 39632 53932
rect 39592 53718 39620 53926
rect 39684 53786 39712 53994
rect 41524 53786 41552 55150
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 39672 53780 39724 53786
rect 39672 53722 39724 53728
rect 41512 53780 41564 53786
rect 41512 53722 41564 53728
rect 39580 53712 39632 53718
rect 39580 53654 39632 53660
rect 38660 53576 38712 53582
rect 38660 53518 38712 53524
rect 35348 53508 35400 53514
rect 35348 53450 35400 53456
rect 37556 53508 37608 53514
rect 37556 53450 37608 53456
rect 39592 53242 39620 53654
rect 39580 53236 39632 53242
rect 39580 53178 39632 53184
rect 39684 52902 39712 53722
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 39672 52896 39724 52902
rect 39672 52838 39724 52844
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 38936 3392 38988 3398
rect 38936 3334 38988 3340
rect 30932 3188 30984 3194
rect 30932 3130 30984 3136
rect 33140 3188 33192 3194
rect 33140 3130 33192 3136
rect 30288 3120 30340 3126
rect 30288 3062 30340 3068
rect 30944 2446 30972 3130
rect 32312 3120 32364 3126
rect 32312 3062 32364 3068
rect 32324 2446 32352 3062
rect 33152 2446 33180 3130
rect 37740 3120 37792 3126
rect 37740 3062 37792 3068
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 36004 2446 36032 2790
rect 37752 2446 37780 3062
rect 38660 2916 38712 2922
rect 38660 2858 38712 2864
rect 38672 2446 38700 2858
rect 38948 2446 38976 3334
rect 39684 2582 39712 52838
rect 55496 52488 55548 52494
rect 55496 52430 55548 52436
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 55404 38956 55456 38962
rect 55404 38898 55456 38904
rect 55416 38758 55444 38898
rect 55404 38752 55456 38758
rect 55404 38694 55456 38700
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 54852 37936 54904 37942
rect 54852 37878 54904 37884
rect 54576 37664 54628 37670
rect 54576 37606 54628 37612
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 53104 36304 53156 36310
rect 53104 36246 53156 36252
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 52368 35012 52420 35018
rect 52368 34954 52420 34960
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 52380 34610 52408 34954
rect 52368 34604 52420 34610
rect 52368 34546 52420 34552
rect 51448 34536 51500 34542
rect 51448 34478 51500 34484
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 48504 33040 48556 33046
rect 48504 32982 48556 32988
rect 43720 26512 43772 26518
rect 43720 26454 43772 26460
rect 42984 12096 43036 12102
rect 42984 12038 43036 12044
rect 42996 3194 43024 12038
rect 43732 3194 43760 26454
rect 44824 3596 44876 3602
rect 44824 3538 44876 3544
rect 44836 3194 44864 3538
rect 48516 3534 48544 32982
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 49056 31272 49108 31278
rect 49056 31214 49108 31220
rect 48504 3528 48556 3534
rect 48504 3470 48556 3476
rect 45744 3392 45796 3398
rect 45744 3334 45796 3340
rect 48320 3392 48372 3398
rect 48320 3334 48372 3340
rect 42984 3188 43036 3194
rect 42984 3130 43036 3136
rect 43720 3188 43772 3194
rect 43720 3130 43772 3136
rect 44824 3188 44876 3194
rect 44824 3130 44876 3136
rect 40316 2984 40368 2990
rect 40316 2926 40368 2932
rect 39672 2576 39724 2582
rect 39672 2518 39724 2524
rect 40328 2446 40356 2926
rect 42996 2446 43024 3130
rect 43732 2446 43760 3130
rect 44836 2446 44864 3130
rect 45756 2446 45784 3334
rect 48332 2446 48360 3334
rect 49068 2446 49096 31214
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50160 4004 50212 4010
rect 50160 3946 50212 3952
rect 50172 2990 50200 3946
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 51460 3194 51488 34478
rect 53116 3534 53144 36246
rect 54588 35894 54616 37606
rect 54588 35866 54708 35894
rect 54392 34400 54444 34406
rect 54392 34342 54444 34348
rect 54404 33522 54432 34342
rect 54392 33516 54444 33522
rect 54392 33458 54444 33464
rect 54484 31816 54536 31822
rect 54484 31758 54536 31764
rect 54496 31346 54524 31758
rect 54484 31340 54536 31346
rect 54484 31282 54536 31288
rect 53840 8356 53892 8362
rect 53840 8298 53892 8304
rect 53852 3670 53880 8298
rect 53840 3664 53892 3670
rect 53840 3606 53892 3612
rect 54680 3534 54708 35866
rect 54760 33448 54812 33454
rect 54760 33390 54812 33396
rect 53104 3528 53156 3534
rect 53104 3470 53156 3476
rect 54668 3528 54720 3534
rect 54668 3470 54720 3476
rect 52920 3392 52972 3398
rect 52920 3334 52972 3340
rect 54392 3392 54444 3398
rect 54392 3334 54444 3340
rect 51448 3188 51500 3194
rect 51448 3130 51500 3136
rect 50160 2984 50212 2990
rect 50160 2926 50212 2932
rect 50620 2984 50672 2990
rect 50620 2926 50672 2932
rect 50632 2446 50660 2926
rect 51460 2446 51488 3130
rect 52932 2446 52960 3334
rect 54404 2446 54432 3334
rect 54680 3194 54708 3470
rect 54668 3188 54720 3194
rect 54668 3130 54720 3136
rect 54484 2984 54536 2990
rect 54772 2972 54800 33390
rect 54864 27946 54892 37878
rect 55416 37874 55444 38694
rect 55508 37942 55536 52430
rect 56416 39840 56468 39846
rect 56416 39782 56468 39788
rect 56428 39506 56456 39782
rect 56048 39500 56100 39506
rect 56048 39442 56100 39448
rect 56416 39500 56468 39506
rect 56416 39442 56468 39448
rect 56060 38894 56088 39442
rect 56140 39296 56192 39302
rect 56140 39238 56192 39244
rect 56600 39296 56652 39302
rect 56600 39238 56652 39244
rect 56152 38962 56180 39238
rect 56140 38956 56192 38962
rect 56140 38898 56192 38904
rect 56048 38888 56100 38894
rect 56048 38830 56100 38836
rect 55956 38752 56008 38758
rect 55956 38694 56008 38700
rect 55496 37936 55548 37942
rect 55864 37936 55916 37942
rect 55548 37896 55864 37924
rect 55496 37878 55548 37884
rect 55864 37878 55916 37884
rect 55404 37868 55456 37874
rect 55404 37810 55456 37816
rect 55416 36106 55444 37810
rect 55404 36100 55456 36106
rect 55404 36042 55456 36048
rect 55772 35148 55824 35154
rect 55772 35090 55824 35096
rect 55784 34950 55812 35090
rect 55036 34944 55088 34950
rect 55036 34886 55088 34892
rect 55772 34944 55824 34950
rect 55772 34886 55824 34892
rect 55048 34542 55076 34886
rect 55312 34740 55364 34746
rect 55312 34682 55364 34688
rect 55324 34610 55352 34682
rect 55312 34604 55364 34610
rect 55312 34546 55364 34552
rect 55036 34536 55088 34542
rect 55036 34478 55088 34484
rect 55588 34468 55640 34474
rect 55588 34410 55640 34416
rect 55600 34202 55628 34410
rect 55588 34196 55640 34202
rect 55588 34138 55640 34144
rect 55784 32774 55812 34886
rect 55864 34536 55916 34542
rect 55864 34478 55916 34484
rect 55772 32768 55824 32774
rect 55772 32710 55824 32716
rect 55784 32570 55812 32710
rect 55772 32564 55824 32570
rect 55772 32506 55824 32512
rect 55784 31958 55812 32506
rect 55772 31952 55824 31958
rect 55772 31894 55824 31900
rect 55588 29504 55640 29510
rect 55588 29446 55640 29452
rect 54852 27940 54904 27946
rect 54852 27882 54904 27888
rect 55404 6792 55456 6798
rect 55404 6734 55456 6740
rect 54536 2944 54800 2972
rect 54484 2926 54536 2932
rect 55416 2650 55444 6734
rect 55600 3466 55628 29446
rect 55876 25770 55904 34478
rect 55864 25764 55916 25770
rect 55864 25706 55916 25712
rect 55680 13184 55732 13190
rect 55680 13126 55732 13132
rect 55692 12238 55720 13126
rect 55680 12232 55732 12238
rect 55680 12174 55732 12180
rect 55864 6248 55916 6254
rect 55864 6190 55916 6196
rect 55588 3460 55640 3466
rect 55588 3402 55640 3408
rect 55496 3392 55548 3398
rect 55496 3334 55548 3340
rect 55772 3392 55824 3398
rect 55772 3334 55824 3340
rect 55404 2644 55456 2650
rect 55404 2586 55456 2592
rect 55508 2446 55536 3334
rect 55784 2446 55812 3334
rect 55876 3194 55904 6190
rect 55968 4146 55996 38694
rect 56060 38214 56088 38830
rect 56048 38208 56100 38214
rect 56048 38150 56100 38156
rect 56060 37806 56088 38150
rect 56048 37800 56100 37806
rect 56048 37742 56100 37748
rect 56508 37800 56560 37806
rect 56508 37742 56560 37748
rect 56060 37466 56088 37742
rect 56048 37460 56100 37466
rect 56048 37402 56100 37408
rect 56520 36582 56548 37742
rect 56508 36576 56560 36582
rect 56508 36518 56560 36524
rect 56520 36242 56548 36518
rect 56508 36236 56560 36242
rect 56508 36178 56560 36184
rect 56324 36100 56376 36106
rect 56324 36042 56376 36048
rect 56336 35154 56364 36042
rect 56520 35894 56548 36178
rect 56428 35866 56548 35894
rect 56428 35494 56456 35866
rect 56416 35488 56468 35494
rect 56416 35430 56468 35436
rect 56324 35148 56376 35154
rect 56324 35090 56376 35096
rect 56428 34406 56456 35430
rect 56416 34400 56468 34406
rect 56416 34342 56468 34348
rect 56428 32910 56456 34342
rect 56416 32904 56468 32910
rect 56416 32846 56468 32852
rect 56428 32230 56456 32846
rect 56416 32224 56468 32230
rect 56416 32166 56468 32172
rect 56232 31952 56284 31958
rect 56232 31894 56284 31900
rect 56140 29572 56192 29578
rect 56140 29514 56192 29520
rect 56152 22778 56180 29514
rect 56140 22772 56192 22778
rect 56140 22714 56192 22720
rect 56244 16574 56272 31894
rect 56428 31142 56456 32166
rect 56416 31136 56468 31142
rect 56416 31078 56468 31084
rect 56152 16546 56272 16574
rect 56152 12434 56180 16546
rect 56428 15366 56456 31078
rect 56612 30818 56640 39238
rect 56704 34746 56732 55354
rect 56888 52494 56916 56646
rect 57072 56506 57100 56782
rect 57060 56500 57112 56506
rect 57060 56442 57112 56448
rect 57532 56438 57560 56782
rect 57704 56704 57756 56710
rect 57704 56646 57756 56652
rect 57520 56432 57572 56438
rect 57520 56374 57572 56380
rect 56876 52488 56928 52494
rect 56876 52430 56928 52436
rect 57336 48544 57388 48550
rect 57336 48486 57388 48492
rect 56784 43648 56836 43654
rect 56784 43590 56836 43596
rect 56692 34740 56744 34746
rect 56692 34682 56744 34688
rect 56796 32842 56824 43590
rect 57060 40384 57112 40390
rect 57060 40326 57112 40332
rect 56876 39296 56928 39302
rect 56876 39238 56928 39244
rect 56888 34218 56916 39238
rect 57072 38706 57100 40326
rect 57244 40180 57296 40186
rect 57244 40122 57296 40128
rect 57256 39438 57284 40122
rect 57244 39432 57296 39438
rect 57244 39374 57296 39380
rect 57348 39098 57376 48486
rect 57612 40928 57664 40934
rect 57612 40870 57664 40876
rect 57152 39092 57204 39098
rect 57152 39034 57204 39040
rect 57336 39092 57388 39098
rect 57336 39034 57388 39040
rect 56980 38678 57100 38706
rect 56980 35894 57008 38678
rect 57058 38584 57114 38593
rect 57058 38519 57060 38528
rect 57112 38519 57114 38528
rect 57060 38490 57112 38496
rect 57164 37482 57192 39034
rect 57164 37454 57376 37482
rect 56980 35866 57284 35894
rect 57152 35284 57204 35290
rect 57152 35226 57204 35232
rect 57164 35154 57192 35226
rect 57152 35148 57204 35154
rect 57152 35090 57204 35096
rect 56888 34190 57192 34218
rect 56968 34128 57020 34134
rect 56968 34070 57020 34076
rect 56876 33312 56928 33318
rect 56876 33254 56928 33260
rect 56784 32836 56836 32842
rect 56784 32778 56836 32784
rect 56612 30790 56732 30818
rect 56508 27328 56560 27334
rect 56508 27270 56560 27276
rect 56520 26382 56548 27270
rect 56508 26376 56560 26382
rect 56508 26318 56560 26324
rect 56704 26234 56732 30790
rect 56888 29050 56916 33254
rect 56980 32910 57008 34070
rect 56968 32904 57020 32910
rect 56968 32846 57020 32852
rect 57060 32768 57112 32774
rect 57060 32710 57112 32716
rect 56968 32020 57020 32026
rect 56968 31962 57020 31968
rect 56980 31890 57008 31962
rect 56968 31884 57020 31890
rect 56968 31826 57020 31832
rect 56968 31408 57020 31414
rect 56968 31350 57020 31356
rect 56980 30326 57008 31350
rect 56968 30320 57020 30326
rect 56968 30262 57020 30268
rect 56980 29510 57008 30262
rect 56968 29504 57020 29510
rect 56968 29446 57020 29452
rect 56888 29022 57008 29050
rect 56980 28966 57008 29022
rect 56968 28960 57020 28966
rect 56968 28902 57020 28908
rect 56784 28416 56836 28422
rect 56784 28358 56836 28364
rect 56796 28150 56824 28358
rect 56784 28144 56836 28150
rect 56784 28086 56836 28092
rect 56612 26206 56732 26234
rect 56508 25152 56560 25158
rect 56508 25094 56560 25100
rect 56520 22098 56548 25094
rect 56508 22092 56560 22098
rect 56508 22034 56560 22040
rect 56416 15360 56468 15366
rect 56416 15302 56468 15308
rect 56428 12434 56456 15302
rect 56060 12406 56180 12434
rect 56244 12406 56456 12434
rect 56060 6798 56088 12406
rect 56140 8560 56192 8566
rect 56140 8502 56192 8508
rect 56048 6792 56100 6798
rect 56048 6734 56100 6740
rect 55956 4140 56008 4146
rect 55956 4082 56008 4088
rect 55968 3534 55996 4082
rect 55956 3528 56008 3534
rect 55956 3470 56008 3476
rect 55864 3188 55916 3194
rect 55864 3130 55916 3136
rect 56048 3052 56100 3058
rect 56048 2994 56100 3000
rect 55956 2848 56008 2854
rect 55956 2790 56008 2796
rect 55968 2446 55996 2790
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 29828 2440 29880 2446
rect 29828 2382 29880 2388
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38936 2440 38988 2446
rect 38936 2382 38988 2388
rect 40316 2440 40368 2446
rect 40316 2382 40368 2388
rect 42984 2440 43036 2446
rect 42984 2382 43036 2388
rect 43720 2440 43772 2446
rect 43720 2382 43772 2388
rect 44824 2440 44876 2446
rect 44824 2382 44876 2388
rect 45744 2440 45796 2446
rect 45744 2382 45796 2388
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 50620 2440 50672 2446
rect 50620 2382 50672 2388
rect 51448 2440 51500 2446
rect 51448 2382 51500 2388
rect 52920 2440 52972 2446
rect 52920 2382 52972 2388
rect 54392 2440 54444 2446
rect 54392 2382 54444 2388
rect 55496 2440 55548 2446
rect 55496 2382 55548 2388
rect 55772 2440 55824 2446
rect 55772 2382 55824 2388
rect 55956 2440 56008 2446
rect 55956 2382 56008 2388
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 29920 2304 29972 2310
rect 29920 2246 29972 2252
rect 31024 2304 31076 2310
rect 31024 2246 31076 2252
rect 32128 2304 32180 2310
rect 32128 2246 32180 2252
rect 33232 2304 33284 2310
rect 33232 2246 33284 2252
rect 34336 2304 34388 2310
rect 34336 2246 34388 2252
rect 28828 800 28856 2246
rect 29932 800 29960 2246
rect 31036 800 31064 2246
rect 32140 800 32168 2246
rect 33244 800 33272 2246
rect 34348 800 34376 2246
rect 36004 1714 36032 2382
rect 36544 2304 36596 2310
rect 36544 2246 36596 2252
rect 37648 2304 37700 2310
rect 37648 2246 37700 2252
rect 38752 2304 38804 2310
rect 38752 2246 38804 2252
rect 39856 2304 39908 2310
rect 39856 2246 39908 2252
rect 40960 2304 41012 2310
rect 40960 2246 41012 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 42064 2304 42116 2310
rect 42064 2246 42116 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 44272 2304 44324 2310
rect 44272 2246 44324 2252
rect 45376 2304 45428 2310
rect 45376 2246 45428 2252
rect 46480 2304 46532 2310
rect 46480 2246 46532 2252
rect 47584 2304 47636 2310
rect 47584 2246 47636 2252
rect 48688 2304 48740 2310
rect 48688 2246 48740 2252
rect 49792 2304 49844 2310
rect 49792 2246 49844 2252
rect 50896 2304 50948 2310
rect 50896 2246 50948 2252
rect 52000 2304 52052 2310
rect 52000 2246 52052 2252
rect 53104 2304 53156 2310
rect 53104 2246 53156 2252
rect 54208 2304 54260 2310
rect 54208 2246 54260 2252
rect 55312 2304 55364 2310
rect 55312 2246 55364 2252
rect 35820 1686 36032 1714
rect 35452 870 35572 898
rect 35452 800 35480 870
rect 2318 0 2374 800
rect 3422 0 3478 800
rect 4526 0 4582 800
rect 5630 0 5686 800
rect 6734 0 6790 800
rect 7838 0 7894 800
rect 8942 0 8998 800
rect 10046 0 10102 800
rect 11150 0 11206 800
rect 12254 0 12310 800
rect 13358 0 13414 800
rect 14462 0 14518 800
rect 15566 0 15622 800
rect 16670 0 16726 800
rect 17774 0 17830 800
rect 18878 0 18934 800
rect 19982 0 20038 800
rect 21086 0 21142 800
rect 22190 0 22246 800
rect 23294 0 23350 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26606 0 26662 800
rect 27710 0 27766 800
rect 28814 0 28870 800
rect 29918 0 29974 800
rect 31022 0 31078 800
rect 32126 0 32182 800
rect 33230 0 33286 800
rect 34334 0 34390 800
rect 35438 0 35494 800
rect 35544 762 35572 870
rect 35820 762 35848 1686
rect 36556 800 36584 2246
rect 37660 800 37688 2246
rect 38764 800 38792 2246
rect 39868 800 39896 2246
rect 40972 800 41000 2246
rect 41892 2106 41920 2246
rect 41880 2100 41932 2106
rect 41880 2042 41932 2048
rect 42076 800 42104 2246
rect 43180 800 43208 2246
rect 44284 800 44312 2246
rect 45388 800 45416 2246
rect 46492 800 46520 2246
rect 47596 800 47624 2246
rect 48700 800 48728 2246
rect 49804 800 49832 2246
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50908 800 50936 2246
rect 52012 800 52040 2246
rect 53116 800 53144 2246
rect 54220 800 54248 2246
rect 55324 800 55352 2246
rect 56060 1873 56088 2994
rect 56152 2582 56180 8502
rect 56140 2576 56192 2582
rect 56140 2518 56192 2524
rect 56244 2378 56272 12406
rect 56508 8832 56560 8838
rect 56508 8774 56560 8780
rect 56324 4480 56376 4486
rect 56324 4422 56376 4428
rect 56336 2689 56364 4422
rect 56520 4078 56548 8774
rect 56612 4146 56640 26206
rect 57072 24342 57100 32710
rect 57164 30190 57192 34190
rect 57152 30184 57204 30190
rect 57152 30126 57204 30132
rect 57152 30048 57204 30054
rect 57152 29990 57204 29996
rect 57164 29578 57192 29990
rect 57152 29572 57204 29578
rect 57152 29514 57204 29520
rect 57152 29028 57204 29034
rect 57152 28970 57204 28976
rect 57164 28801 57192 28970
rect 57150 28792 57206 28801
rect 57150 28727 57206 28736
rect 57152 28212 57204 28218
rect 57152 28154 57204 28160
rect 57164 27538 57192 28154
rect 57256 27538 57284 35866
rect 57348 29306 57376 37454
rect 57428 37120 57480 37126
rect 57428 37062 57480 37068
rect 57440 36174 57468 37062
rect 57428 36168 57480 36174
rect 57428 36110 57480 36116
rect 57520 35488 57572 35494
rect 57520 35430 57572 35436
rect 57532 35154 57560 35430
rect 57520 35148 57572 35154
rect 57520 35090 57572 35096
rect 57520 32836 57572 32842
rect 57520 32778 57572 32784
rect 57532 32570 57560 32778
rect 57520 32564 57572 32570
rect 57520 32506 57572 32512
rect 57428 32224 57480 32230
rect 57428 32166 57480 32172
rect 57440 31890 57468 32166
rect 57520 31952 57572 31958
rect 57520 31894 57572 31900
rect 57428 31884 57480 31890
rect 57428 31826 57480 31832
rect 57532 31482 57560 31894
rect 57520 31476 57572 31482
rect 57520 31418 57572 31424
rect 57624 31090 57652 40870
rect 57716 39438 57744 56646
rect 58084 56370 58112 57394
rect 58164 57248 58216 57254
rect 58164 57190 58216 57196
rect 58072 56364 58124 56370
rect 58072 56306 58124 56312
rect 58176 56302 58204 57190
rect 58348 56840 58400 56846
rect 58348 56782 58400 56788
rect 58360 56545 58388 56782
rect 58346 56536 58402 56545
rect 58346 56471 58402 56480
rect 58452 56370 58480 58103
rect 59176 56704 59228 56710
rect 59176 56646 59228 56652
rect 58440 56364 58492 56370
rect 58440 56306 58492 56312
rect 58164 56296 58216 56302
rect 58164 56238 58216 56244
rect 58164 56160 58216 56166
rect 58164 56102 58216 56108
rect 57980 55276 58032 55282
rect 57980 55218 58032 55224
rect 57992 55162 58020 55218
rect 57900 55134 58020 55162
rect 57900 54913 57928 55134
rect 57886 54904 57942 54913
rect 57886 54839 57942 54848
rect 57980 49088 58032 49094
rect 57980 49030 58032 49036
rect 57796 42560 57848 42566
rect 57796 42502 57848 42508
rect 57704 39432 57756 39438
rect 57704 39374 57756 39380
rect 57808 35986 57836 42502
rect 57888 40112 57940 40118
rect 57888 40054 57940 40060
rect 57900 39409 57928 40054
rect 57886 39400 57942 39409
rect 57992 39370 58020 49030
rect 57886 39335 57942 39344
rect 57980 39364 58032 39370
rect 57980 39306 58032 39312
rect 58176 38962 58204 56102
rect 58452 55962 58480 56306
rect 58440 55956 58492 55962
rect 58440 55898 58492 55904
rect 58348 55752 58400 55758
rect 58346 55720 58348 55729
rect 58400 55720 58402 55729
rect 58346 55655 58402 55664
rect 58348 54528 58400 54534
rect 58348 54470 58400 54476
rect 58360 54194 58388 54470
rect 58348 54188 58400 54194
rect 58348 54130 58400 54136
rect 58360 54097 58388 54130
rect 58346 54088 58402 54097
rect 58346 54023 58402 54032
rect 58900 53984 58952 53990
rect 58900 53926 58952 53932
rect 58348 53576 58400 53582
rect 58348 53518 58400 53524
rect 58360 53281 58388 53518
rect 58532 53440 58584 53446
rect 58532 53382 58584 53388
rect 58346 53272 58402 53281
rect 58346 53207 58402 53216
rect 58348 52488 58400 52494
rect 58346 52456 58348 52465
rect 58400 52456 58402 52465
rect 58346 52391 58402 52400
rect 58348 52012 58400 52018
rect 58348 51954 58400 51960
rect 58360 51649 58388 51954
rect 58346 51640 58402 51649
rect 58346 51575 58402 51584
rect 58348 51264 58400 51270
rect 58348 51206 58400 51212
rect 58360 50930 58388 51206
rect 58348 50924 58400 50930
rect 58348 50866 58400 50872
rect 58360 50833 58388 50866
rect 58346 50824 58402 50833
rect 58346 50759 58402 50768
rect 58348 50312 58400 50318
rect 58348 50254 58400 50260
rect 58360 50017 58388 50254
rect 58440 50176 58492 50182
rect 58440 50118 58492 50124
rect 58346 50008 58402 50017
rect 58346 49943 58402 49952
rect 58348 49224 58400 49230
rect 58346 49192 58348 49201
rect 58400 49192 58402 49201
rect 58346 49127 58402 49136
rect 58348 48748 58400 48754
rect 58348 48690 58400 48696
rect 58360 48385 58388 48690
rect 58346 48376 58402 48385
rect 58346 48311 58402 48320
rect 58348 48000 58400 48006
rect 58348 47942 58400 47948
rect 58360 47666 58388 47942
rect 58348 47660 58400 47666
rect 58348 47602 58400 47608
rect 58360 47569 58388 47602
rect 58346 47560 58402 47569
rect 58346 47495 58402 47504
rect 58256 47456 58308 47462
rect 58256 47398 58308 47404
rect 58164 38956 58216 38962
rect 58164 38898 58216 38904
rect 58176 38554 58204 38898
rect 58164 38548 58216 38554
rect 58164 38490 58216 38496
rect 58268 37942 58296 47398
rect 58348 47048 58400 47054
rect 58348 46990 58400 46996
rect 58360 46753 58388 46990
rect 58346 46744 58402 46753
rect 58346 46679 58402 46688
rect 58348 45960 58400 45966
rect 58346 45928 58348 45937
rect 58400 45928 58402 45937
rect 58346 45863 58402 45872
rect 58348 45484 58400 45490
rect 58348 45426 58400 45432
rect 58360 45121 58388 45426
rect 58346 45112 58402 45121
rect 58346 45047 58402 45056
rect 58348 44736 58400 44742
rect 58348 44678 58400 44684
rect 58360 44402 58388 44678
rect 58348 44396 58400 44402
rect 58348 44338 58400 44344
rect 58360 44305 58388 44338
rect 58346 44296 58402 44305
rect 58346 44231 58402 44240
rect 58348 43784 58400 43790
rect 58348 43726 58400 43732
rect 58360 43489 58388 43726
rect 58346 43480 58402 43489
rect 58346 43415 58402 43424
rect 58348 42696 58400 42702
rect 58346 42664 58348 42673
rect 58400 42664 58402 42673
rect 58346 42599 58402 42608
rect 58348 42220 58400 42226
rect 58348 42162 58400 42168
rect 58360 41857 58388 42162
rect 58346 41848 58402 41857
rect 58346 41783 58402 41792
rect 58348 41472 58400 41478
rect 58348 41414 58400 41420
rect 58360 41138 58388 41414
rect 58348 41132 58400 41138
rect 58348 41074 58400 41080
rect 58360 41041 58388 41074
rect 58346 41032 58402 41041
rect 58346 40967 58402 40976
rect 58348 40520 58400 40526
rect 58348 40462 58400 40468
rect 58360 40225 58388 40462
rect 58346 40216 58402 40225
rect 58346 40151 58402 40160
rect 58348 38956 58400 38962
rect 58348 38898 58400 38904
rect 58360 38593 58388 38898
rect 58346 38584 58402 38593
rect 58346 38519 58402 38528
rect 58348 38208 58400 38214
rect 58348 38150 58400 38156
rect 58256 37936 58308 37942
rect 58256 37878 58308 37884
rect 58360 37874 58388 38150
rect 58348 37868 58400 37874
rect 58348 37810 58400 37816
rect 58360 37777 58388 37810
rect 58346 37768 58402 37777
rect 58346 37703 58402 37712
rect 57888 37324 57940 37330
rect 57888 37266 57940 37272
rect 57900 36786 57928 37266
rect 58348 37256 58400 37262
rect 58348 37198 58400 37204
rect 58360 36961 58388 37198
rect 58346 36952 58402 36961
rect 57980 36916 58032 36922
rect 58346 36887 58402 36896
rect 57980 36858 58032 36864
rect 57888 36780 57940 36786
rect 57888 36722 57940 36728
rect 57900 36145 57928 36722
rect 57992 36174 58020 36858
rect 58072 36576 58124 36582
rect 58072 36518 58124 36524
rect 57980 36168 58032 36174
rect 57886 36136 57942 36145
rect 57980 36110 58032 36116
rect 57886 36071 57942 36080
rect 57808 35958 57928 35986
rect 57796 33856 57848 33862
rect 57796 33798 57848 33804
rect 57808 33522 57836 33798
rect 57796 33516 57848 33522
rect 57796 33458 57848 33464
rect 57808 32881 57836 33458
rect 57794 32872 57850 32881
rect 57794 32807 57850 32816
rect 57624 31062 57836 31090
rect 57520 30864 57572 30870
rect 57520 30806 57572 30812
rect 57428 30048 57480 30054
rect 57428 29990 57480 29996
rect 57336 29300 57388 29306
rect 57336 29242 57388 29248
rect 57336 28960 57388 28966
rect 57336 28902 57388 28908
rect 57348 28558 57376 28902
rect 57440 28558 57468 29990
rect 57532 29186 57560 30806
rect 57612 30184 57664 30190
rect 57612 30126 57664 30132
rect 57624 29306 57652 30126
rect 57704 29776 57756 29782
rect 57704 29718 57756 29724
rect 57612 29300 57664 29306
rect 57612 29242 57664 29248
rect 57532 29158 57652 29186
rect 57336 28552 57388 28558
rect 57336 28494 57388 28500
rect 57428 28552 57480 28558
rect 57428 28494 57480 28500
rect 57336 28416 57388 28422
rect 57336 28358 57388 28364
rect 57152 27532 57204 27538
rect 57152 27474 57204 27480
rect 57244 27532 57296 27538
rect 57244 27474 57296 27480
rect 57164 27130 57192 27474
rect 57152 27124 57204 27130
rect 57152 27066 57204 27072
rect 57164 25294 57192 27066
rect 57152 25288 57204 25294
rect 57152 25230 57204 25236
rect 57164 24614 57192 25230
rect 57152 24608 57204 24614
rect 57152 24550 57204 24556
rect 57244 24608 57296 24614
rect 57244 24550 57296 24556
rect 57060 24336 57112 24342
rect 57060 24278 57112 24284
rect 57164 13394 57192 24550
rect 57256 15570 57284 24550
rect 57348 16574 57376 28358
rect 57440 28218 57468 28494
rect 57428 28212 57480 28218
rect 57428 28154 57480 28160
rect 57624 27538 57652 29158
rect 57716 28626 57744 29718
rect 57704 28620 57756 28626
rect 57704 28562 57756 28568
rect 57716 28218 57744 28562
rect 57704 28212 57756 28218
rect 57704 28154 57756 28160
rect 57716 27606 57744 28154
rect 57704 27600 57756 27606
rect 57704 27542 57756 27548
rect 57612 27532 57664 27538
rect 57612 27474 57664 27480
rect 57624 26518 57652 27474
rect 57716 27130 57744 27542
rect 57704 27124 57756 27130
rect 57704 27066 57756 27072
rect 57612 26512 57664 26518
rect 57612 26454 57664 26460
rect 57520 26376 57572 26382
rect 57520 26318 57572 26324
rect 57532 26042 57560 26318
rect 57520 26036 57572 26042
rect 57520 25978 57572 25984
rect 57428 25492 57480 25498
rect 57428 25434 57480 25440
rect 57440 25294 57468 25434
rect 57716 25362 57744 27066
rect 57808 25430 57836 31062
rect 57900 28490 57928 35958
rect 57980 35828 58032 35834
rect 57980 35770 58032 35776
rect 57992 35222 58020 35770
rect 57980 35216 58032 35222
rect 57980 35158 58032 35164
rect 58084 35154 58112 36518
rect 58348 35692 58400 35698
rect 58348 35634 58400 35640
rect 58164 35488 58216 35494
rect 58164 35430 58216 35436
rect 58072 35148 58124 35154
rect 58072 35090 58124 35096
rect 58072 35012 58124 35018
rect 58072 34954 58124 34960
rect 57980 33652 58032 33658
rect 57980 33594 58032 33600
rect 57992 32910 58020 33594
rect 57980 32904 58032 32910
rect 57980 32846 58032 32852
rect 57980 31816 58032 31822
rect 57980 31758 58032 31764
rect 57888 28484 57940 28490
rect 57888 28426 57940 28432
rect 57992 26234 58020 31758
rect 58084 26518 58112 34954
rect 58176 34678 58204 35430
rect 58360 35329 58388 35634
rect 58346 35320 58402 35329
rect 58346 35255 58402 35264
rect 58164 34672 58216 34678
rect 58164 34614 58216 34620
rect 58348 34604 58400 34610
rect 58348 34546 58400 34552
rect 58360 34513 58388 34546
rect 58346 34504 58402 34513
rect 58346 34439 58402 34448
rect 58164 34400 58216 34406
rect 58164 34342 58216 34348
rect 58176 31890 58204 34342
rect 58348 33992 58400 33998
rect 58348 33934 58400 33940
rect 58360 33697 58388 33934
rect 58346 33688 58402 33697
rect 58346 33623 58402 33632
rect 58348 32428 58400 32434
rect 58348 32370 58400 32376
rect 58256 32224 58308 32230
rect 58256 32166 58308 32172
rect 58164 31884 58216 31890
rect 58164 31826 58216 31832
rect 58164 31340 58216 31346
rect 58164 31282 58216 31288
rect 58176 31249 58204 31282
rect 58162 31240 58218 31249
rect 58162 31175 58218 31184
rect 58176 30938 58204 31175
rect 58164 30932 58216 30938
rect 58164 30874 58216 30880
rect 58268 29646 58296 32166
rect 58360 32065 58388 32370
rect 58346 32056 58402 32065
rect 58346 31991 58402 32000
rect 58452 30870 58480 50118
rect 58544 33658 58572 53382
rect 58716 52624 58768 52630
rect 58716 52566 58768 52572
rect 58624 47184 58676 47190
rect 58624 47126 58676 47132
rect 58636 36038 58664 47126
rect 58624 36032 58676 36038
rect 58624 35974 58676 35980
rect 58532 33652 58584 33658
rect 58532 33594 58584 33600
rect 58532 31136 58584 31142
rect 58532 31078 58584 31084
rect 58440 30864 58492 30870
rect 58440 30806 58492 30812
rect 58440 30728 58492 30734
rect 58440 30670 58492 30676
rect 58348 30592 58400 30598
rect 58348 30534 58400 30540
rect 58256 29640 58308 29646
rect 58256 29582 58308 29588
rect 58360 27538 58388 30534
rect 58452 30433 58480 30670
rect 58438 30424 58494 30433
rect 58438 30359 58440 30368
rect 58492 30359 58494 30368
rect 58440 30330 58492 30336
rect 58438 29608 58494 29617
rect 58438 29543 58494 29552
rect 58452 29170 58480 29543
rect 58440 29164 58492 29170
rect 58440 29106 58492 29112
rect 58440 28076 58492 28082
rect 58440 28018 58492 28024
rect 58452 27985 58480 28018
rect 58438 27976 58494 27985
rect 58438 27911 58494 27920
rect 58348 27532 58400 27538
rect 58348 27474 58400 27480
rect 58164 27464 58216 27470
rect 58164 27406 58216 27412
rect 58072 26512 58124 26518
rect 58072 26454 58124 26460
rect 57992 26206 58112 26234
rect 57796 25424 57848 25430
rect 57796 25366 57848 25372
rect 57704 25356 57756 25362
rect 57704 25298 57756 25304
rect 57428 25288 57480 25294
rect 57428 25230 57480 25236
rect 57716 24614 57744 25298
rect 58084 24682 58112 26206
rect 58176 25378 58204 27406
rect 58346 27160 58402 27169
rect 58346 27095 58402 27104
rect 58360 26994 58388 27095
rect 58348 26988 58400 26994
rect 58348 26930 58400 26936
rect 58360 26586 58388 26930
rect 58348 26580 58400 26586
rect 58348 26522 58400 26528
rect 58348 26376 58400 26382
rect 58346 26344 58348 26353
rect 58400 26344 58402 26353
rect 58346 26279 58402 26288
rect 58348 25900 58400 25906
rect 58348 25842 58400 25848
rect 58360 25537 58388 25842
rect 58346 25528 58402 25537
rect 58346 25463 58402 25472
rect 58176 25350 58296 25378
rect 58544 25362 58572 31078
rect 58728 28558 58756 52566
rect 58808 50720 58860 50726
rect 58808 50662 58860 50668
rect 58716 28552 58768 28558
rect 58716 28494 58768 28500
rect 58716 28144 58768 28150
rect 58716 28086 58768 28092
rect 58164 25288 58216 25294
rect 58164 25230 58216 25236
rect 58072 24676 58124 24682
rect 58072 24618 58124 24624
rect 57704 24608 57756 24614
rect 57704 24550 57756 24556
rect 57980 22024 58032 22030
rect 57980 21966 58032 21972
rect 57992 16574 58020 21966
rect 58176 21690 58204 25230
rect 58164 21684 58216 21690
rect 58164 21626 58216 21632
rect 58268 21146 58296 25350
rect 58532 25356 58584 25362
rect 58532 25298 58584 25304
rect 58348 24812 58400 24818
rect 58348 24754 58400 24760
rect 58360 24721 58388 24754
rect 58346 24712 58402 24721
rect 58346 24647 58402 24656
rect 58360 24410 58388 24647
rect 58348 24404 58400 24410
rect 58348 24346 58400 24352
rect 58348 24200 58400 24206
rect 58348 24142 58400 24148
rect 58360 23905 58388 24142
rect 58346 23896 58402 23905
rect 58346 23831 58402 23840
rect 58728 23322 58756 28086
rect 58820 25498 58848 50662
rect 58912 31958 58940 53926
rect 59084 51808 59136 51814
rect 59084 51750 59136 51756
rect 58992 42016 59044 42022
rect 58992 41958 59044 41964
rect 58900 31952 58952 31958
rect 58900 31894 58952 31900
rect 59004 29578 59032 41958
rect 59096 31414 59124 51750
rect 59188 36922 59216 56646
rect 59544 55616 59596 55622
rect 59544 55558 59596 55564
rect 59268 45280 59320 45286
rect 59268 45222 59320 45228
rect 59176 36916 59228 36922
rect 59176 36858 59228 36864
rect 59280 34542 59308 45222
rect 59360 44192 59412 44198
rect 59360 44134 59412 44140
rect 59268 34536 59320 34542
rect 59268 34478 59320 34484
rect 59372 32026 59400 44134
rect 59452 36100 59504 36106
rect 59452 36042 59504 36048
rect 59360 32020 59412 32026
rect 59360 31962 59412 31968
rect 59084 31408 59136 31414
rect 59084 31350 59136 31356
rect 58992 29572 59044 29578
rect 58992 29514 59044 29520
rect 59464 27130 59492 36042
rect 59556 35834 59584 55558
rect 59636 45824 59688 45830
rect 59636 45766 59688 45772
rect 59544 35828 59596 35834
rect 59544 35770 59596 35776
rect 59648 35290 59676 45766
rect 59636 35284 59688 35290
rect 59636 35226 59688 35232
rect 59452 27124 59504 27130
rect 59452 27066 59504 27072
rect 58808 25492 58860 25498
rect 58808 25434 58860 25440
rect 58820 23866 58848 25434
rect 58808 23860 58860 23866
rect 58808 23802 58860 23808
rect 58716 23316 58768 23322
rect 58716 23258 58768 23264
rect 58348 23112 58400 23118
rect 58346 23080 58348 23089
rect 58400 23080 58402 23089
rect 58346 23015 58402 23024
rect 58348 22636 58400 22642
rect 58348 22578 58400 22584
rect 58360 22273 58388 22578
rect 58346 22264 58402 22273
rect 58346 22199 58402 22208
rect 58348 21548 58400 21554
rect 58348 21490 58400 21496
rect 58360 21457 58388 21490
rect 58346 21448 58402 21457
rect 58346 21383 58402 21392
rect 58256 21140 58308 21146
rect 58256 21082 58308 21088
rect 58348 20936 58400 20942
rect 58348 20878 58400 20884
rect 58360 20641 58388 20878
rect 58346 20632 58402 20641
rect 58346 20567 58402 20576
rect 58348 19848 58400 19854
rect 58346 19816 58348 19825
rect 58400 19816 58402 19825
rect 58346 19751 58402 19760
rect 58624 19712 58676 19718
rect 58624 19654 58676 19660
rect 58440 19508 58492 19514
rect 58440 19450 58492 19456
rect 58348 19372 58400 19378
rect 58348 19314 58400 19320
rect 58360 19009 58388 19314
rect 58346 19000 58402 19009
rect 58346 18935 58348 18944
rect 58400 18935 58402 18944
rect 58348 18906 58400 18912
rect 58348 18284 58400 18290
rect 58348 18226 58400 18232
rect 58360 18193 58388 18226
rect 58346 18184 58402 18193
rect 58346 18119 58402 18128
rect 58348 17672 58400 17678
rect 58348 17614 58400 17620
rect 58256 17536 58308 17542
rect 58256 17478 58308 17484
rect 57348 16546 57468 16574
rect 57992 16546 58112 16574
rect 57244 15564 57296 15570
rect 57244 15506 57296 15512
rect 57256 14074 57284 15506
rect 57336 14816 57388 14822
rect 57336 14758 57388 14764
rect 57244 14068 57296 14074
rect 57244 14010 57296 14016
rect 57348 13394 57376 14758
rect 57152 13388 57204 13394
rect 57152 13330 57204 13336
rect 57336 13388 57388 13394
rect 57336 13330 57388 13336
rect 57164 12986 57192 13330
rect 57152 12980 57204 12986
rect 57152 12922 57204 12928
rect 57164 12434 57192 12922
rect 57336 12708 57388 12714
rect 57336 12650 57388 12656
rect 56980 12406 57192 12434
rect 56692 11552 56744 11558
rect 56692 11494 56744 11500
rect 56704 6322 56732 11494
rect 56980 11218 57008 12406
rect 57244 11620 57296 11626
rect 57244 11562 57296 11568
rect 57152 11348 57204 11354
rect 57152 11290 57204 11296
rect 56968 11212 57020 11218
rect 56968 11154 57020 11160
rect 56980 10962 57008 11154
rect 56888 10934 57008 10962
rect 56888 10810 56916 10934
rect 56876 10804 56928 10810
rect 56876 10746 56928 10752
rect 56968 10804 57020 10810
rect 56968 10746 57020 10752
rect 56888 9058 56916 10746
rect 56980 9722 57008 10746
rect 56968 9716 57020 9722
rect 56968 9658 57020 9664
rect 56888 9042 57008 9058
rect 56888 9036 57020 9042
rect 56888 9030 56968 9036
rect 56968 8978 57020 8984
rect 56876 8832 56928 8838
rect 56876 8774 56928 8780
rect 56888 8566 56916 8774
rect 56876 8560 56928 8566
rect 56876 8502 56928 8508
rect 56980 8498 57008 8978
rect 56968 8492 57020 8498
rect 56968 8434 57020 8440
rect 56980 8090 57008 8434
rect 56968 8084 57020 8090
rect 56968 8026 57020 8032
rect 56980 7290 57008 8026
rect 56888 7262 57008 7290
rect 56888 6798 56916 7262
rect 56968 7200 57020 7206
rect 56968 7142 57020 7148
rect 56980 6798 57008 7142
rect 57060 6996 57112 7002
rect 57060 6938 57112 6944
rect 56876 6792 56928 6798
rect 56876 6734 56928 6740
rect 56968 6792 57020 6798
rect 56968 6734 57020 6740
rect 56888 6322 56916 6734
rect 56692 6316 56744 6322
rect 56692 6258 56744 6264
rect 56876 6316 56928 6322
rect 56876 6258 56928 6264
rect 57072 6118 57100 6938
rect 57060 6112 57112 6118
rect 57060 6054 57112 6060
rect 57072 5846 57100 6054
rect 57060 5840 57112 5846
rect 57060 5782 57112 5788
rect 56692 5704 56744 5710
rect 56692 5646 56744 5652
rect 56600 4140 56652 4146
rect 56600 4082 56652 4088
rect 56508 4072 56560 4078
rect 56508 4014 56560 4020
rect 56612 3534 56640 4082
rect 56600 3528 56652 3534
rect 56600 3470 56652 3476
rect 56704 3194 56732 5646
rect 57072 5370 57100 5782
rect 57060 5364 57112 5370
rect 57060 5306 57112 5312
rect 57164 4146 57192 11290
rect 57256 6474 57284 11562
rect 57348 9042 57376 12650
rect 57440 11626 57468 16546
rect 57796 15904 57848 15910
rect 57796 15846 57848 15852
rect 57704 14068 57756 14074
rect 57704 14010 57756 14016
rect 57716 13394 57744 14010
rect 57704 13388 57756 13394
rect 57704 13330 57756 13336
rect 57428 11620 57480 11626
rect 57428 11562 57480 11568
rect 57428 11348 57480 11354
rect 57428 11290 57480 11296
rect 57440 11150 57468 11290
rect 57716 11218 57744 13330
rect 57704 11212 57756 11218
rect 57704 11154 57756 11160
rect 57428 11144 57480 11150
rect 57428 11086 57480 11092
rect 57716 10810 57744 11154
rect 57704 10804 57756 10810
rect 57704 10746 57756 10752
rect 57808 10554 57836 15846
rect 57886 13288 57942 13297
rect 57886 13223 57942 13232
rect 57900 12850 57928 13223
rect 57888 12844 57940 12850
rect 57888 12786 57940 12792
rect 57900 12442 57928 12786
rect 57888 12436 57940 12442
rect 57888 12378 57940 12384
rect 58084 12306 58112 16546
rect 58164 14272 58216 14278
rect 58164 14214 58216 14220
rect 58072 12300 58124 12306
rect 58072 12242 58124 12248
rect 58072 12096 58124 12102
rect 58072 12038 58124 12044
rect 57980 11144 58032 11150
rect 57980 11086 58032 11092
rect 57440 10526 57836 10554
rect 57336 9036 57388 9042
rect 57336 8978 57388 8984
rect 57256 6446 57376 6474
rect 57244 6112 57296 6118
rect 57244 6054 57296 6060
rect 57152 4140 57204 4146
rect 57152 4082 57204 4088
rect 57256 3534 57284 6054
rect 57348 3890 57376 6446
rect 57440 5778 57468 10526
rect 57612 10464 57664 10470
rect 57612 10406 57664 10412
rect 57518 5944 57574 5953
rect 57518 5879 57574 5888
rect 57428 5772 57480 5778
rect 57428 5714 57480 5720
rect 57532 5370 57560 5879
rect 57624 5778 57652 10406
rect 57704 9716 57756 9722
rect 57704 9658 57756 9664
rect 57716 9042 57744 9658
rect 57796 9172 57848 9178
rect 57796 9114 57848 9120
rect 57704 9036 57756 9042
rect 57704 8978 57756 8984
rect 57716 8430 57744 8978
rect 57704 8424 57756 8430
rect 57704 8366 57756 8372
rect 57716 8090 57744 8366
rect 57704 8084 57756 8090
rect 57704 8026 57756 8032
rect 57716 7002 57744 8026
rect 57704 6996 57756 7002
rect 57704 6938 57756 6944
rect 57704 6860 57756 6866
rect 57704 6802 57756 6808
rect 57612 5772 57664 5778
rect 57612 5714 57664 5720
rect 57716 5710 57744 6802
rect 57704 5704 57756 5710
rect 57704 5646 57756 5652
rect 57716 5574 57744 5646
rect 57704 5568 57756 5574
rect 57704 5510 57756 5516
rect 57520 5364 57572 5370
rect 57520 5306 57572 5312
rect 57808 4826 57836 9114
rect 57992 4826 58020 11086
rect 58084 8634 58112 12038
rect 58176 11286 58204 14214
rect 58268 13546 58296 17478
rect 58360 17377 58388 17614
rect 58346 17368 58402 17377
rect 58346 17303 58402 17312
rect 58348 16584 58400 16590
rect 58346 16552 58348 16561
rect 58400 16552 58402 16561
rect 58346 16487 58402 16496
rect 58348 16108 58400 16114
rect 58348 16050 58400 16056
rect 58360 15745 58388 16050
rect 58346 15736 58402 15745
rect 58346 15671 58348 15680
rect 58400 15671 58402 15680
rect 58348 15642 58400 15648
rect 58348 15020 58400 15026
rect 58348 14962 58400 14968
rect 58360 14929 58388 14962
rect 58346 14920 58402 14929
rect 58346 14855 58402 14864
rect 58348 14408 58400 14414
rect 58348 14350 58400 14356
rect 58360 14113 58388 14350
rect 58346 14104 58402 14113
rect 58452 14074 58480 19450
rect 58346 14039 58402 14048
rect 58440 14068 58492 14074
rect 58440 14010 58492 14016
rect 58268 13518 58572 13546
rect 58256 13320 58308 13326
rect 58256 13262 58308 13268
rect 58164 11280 58216 11286
rect 58164 11222 58216 11228
rect 58268 10266 58296 13262
rect 58346 12472 58402 12481
rect 58346 12407 58402 12416
rect 58360 12238 58388 12407
rect 58348 12232 58400 12238
rect 58348 12174 58400 12180
rect 58348 11756 58400 11762
rect 58348 11698 58400 11704
rect 58360 11665 58388 11698
rect 58346 11656 58402 11665
rect 58346 11591 58402 11600
rect 58348 11144 58400 11150
rect 58348 11086 58400 11092
rect 58256 10260 58308 10266
rect 58256 10202 58308 10208
rect 58164 10056 58216 10062
rect 58162 10024 58164 10033
rect 58216 10024 58218 10033
rect 58162 9959 58218 9968
rect 58164 9580 58216 9586
rect 58164 9522 58216 9528
rect 58176 9217 58204 9522
rect 58360 9450 58388 11086
rect 58438 10840 58494 10849
rect 58438 10775 58494 10784
rect 58452 10674 58480 10775
rect 58440 10668 58492 10674
rect 58440 10610 58492 10616
rect 58452 10198 58480 10610
rect 58440 10192 58492 10198
rect 58440 10134 58492 10140
rect 58348 9444 58400 9450
rect 58348 9386 58400 9392
rect 58162 9208 58218 9217
rect 58162 9143 58218 9152
rect 58348 8968 58400 8974
rect 58348 8910 58400 8916
rect 58256 8832 58308 8838
rect 58256 8774 58308 8780
rect 58072 8628 58124 8634
rect 58072 8570 58124 8576
rect 58164 8492 58216 8498
rect 58164 8434 58216 8440
rect 58176 8401 58204 8434
rect 58162 8392 58218 8401
rect 58162 8327 58218 8336
rect 58176 7478 58204 8327
rect 58268 8090 58296 8774
rect 58360 8634 58388 8910
rect 58348 8628 58400 8634
rect 58348 8570 58400 8576
rect 58544 8566 58572 13518
rect 58636 13462 58664 19654
rect 58808 18080 58860 18086
rect 58808 18022 58860 18028
rect 58820 16574 58848 18022
rect 58820 16546 58940 16574
rect 58808 16448 58860 16454
rect 58808 16390 58860 16396
rect 58624 13456 58676 13462
rect 58624 13398 58676 13404
rect 58716 13388 58768 13394
rect 58716 13330 58768 13336
rect 58624 12300 58676 12306
rect 58624 12242 58676 12248
rect 58532 8560 58584 8566
rect 58532 8502 58584 8508
rect 58256 8084 58308 8090
rect 58256 8026 58308 8032
rect 58348 7880 58400 7886
rect 58348 7822 58400 7828
rect 58360 7585 58388 7822
rect 58346 7576 58402 7585
rect 58346 7511 58348 7520
rect 58400 7511 58402 7520
rect 58348 7482 58400 7488
rect 58164 7472 58216 7478
rect 58360 7451 58388 7482
rect 58164 7414 58216 7420
rect 58348 6792 58400 6798
rect 58346 6760 58348 6769
rect 58400 6760 58402 6769
rect 58346 6695 58402 6704
rect 58164 6656 58216 6662
rect 58164 6598 58216 6604
rect 58176 6458 58204 6598
rect 58164 6452 58216 6458
rect 58164 6394 58216 6400
rect 58348 6316 58400 6322
rect 58348 6258 58400 6264
rect 58164 6112 58216 6118
rect 58164 6054 58216 6060
rect 58176 5914 58204 6054
rect 58360 5953 58388 6258
rect 58346 5944 58402 5953
rect 58164 5908 58216 5914
rect 58346 5879 58402 5888
rect 58164 5850 58216 5856
rect 58256 5568 58308 5574
rect 58256 5510 58308 5516
rect 57796 4820 57848 4826
rect 57796 4762 57848 4768
rect 57980 4820 58032 4826
rect 57980 4762 58032 4768
rect 57520 4616 57572 4622
rect 57520 4558 57572 4564
rect 57428 3936 57480 3942
rect 57348 3884 57428 3890
rect 57348 3878 57480 3884
rect 57348 3862 57468 3878
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 56968 3392 57020 3398
rect 56968 3334 57020 3340
rect 56692 3188 56744 3194
rect 56692 3130 56744 3136
rect 56980 2922 57008 3334
rect 57348 3058 57376 3862
rect 57532 3505 57560 4558
rect 58072 3936 58124 3942
rect 58072 3878 58124 3884
rect 57612 3528 57664 3534
rect 57518 3496 57574 3505
rect 57612 3470 57664 3476
rect 57518 3431 57574 3440
rect 57336 3052 57388 3058
rect 57336 2994 57388 3000
rect 56968 2916 57020 2922
rect 56968 2858 57020 2864
rect 57152 2848 57204 2854
rect 57152 2790 57204 2796
rect 56322 2680 56378 2689
rect 56322 2615 56378 2624
rect 56336 2378 56364 2615
rect 57164 2514 57192 2790
rect 57624 2650 57652 3470
rect 57796 3392 57848 3398
rect 57796 3334 57848 3340
rect 57612 2644 57664 2650
rect 57612 2586 57664 2592
rect 57152 2508 57204 2514
rect 57152 2450 57204 2456
rect 57808 2446 57836 3334
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 57796 2440 57848 2446
rect 57796 2382 57848 2388
rect 56232 2372 56284 2378
rect 56232 2314 56284 2320
rect 56324 2372 56376 2378
rect 56324 2314 56376 2320
rect 56046 1864 56102 1873
rect 56046 1799 56102 1808
rect 56428 800 56456 2382
rect 57520 2304 57572 2310
rect 57520 2246 57572 2252
rect 57532 800 57560 2246
rect 58084 2106 58112 3878
rect 58268 3058 58296 5510
rect 58348 5228 58400 5234
rect 58348 5170 58400 5176
rect 58360 5137 58388 5170
rect 58346 5128 58402 5137
rect 58346 5063 58402 5072
rect 58348 4616 58400 4622
rect 58348 4558 58400 4564
rect 58360 4321 58388 4558
rect 58346 4312 58402 4321
rect 58346 4247 58402 4256
rect 58636 3602 58664 12242
rect 58728 5370 58756 13330
rect 58820 6254 58848 16390
rect 58912 8906 58940 16546
rect 58992 14068 59044 14074
rect 58992 14010 59044 14016
rect 59004 11354 59032 14010
rect 58992 11348 59044 11354
rect 58992 11290 59044 11296
rect 58900 8900 58952 8906
rect 58900 8842 58952 8848
rect 58808 6248 58860 6254
rect 58808 6190 58860 6196
rect 58716 5364 58768 5370
rect 58716 5306 58768 5312
rect 58624 3596 58676 3602
rect 58624 3538 58676 3544
rect 58348 3392 58400 3398
rect 58348 3334 58400 3340
rect 58360 3126 58388 3334
rect 58348 3120 58400 3126
rect 58348 3062 58400 3068
rect 58256 3052 58308 3058
rect 58256 2994 58308 3000
rect 58072 2100 58124 2106
rect 58072 2042 58124 2048
rect 58360 1057 58388 3062
rect 58346 1048 58402 1057
rect 58346 983 58402 992
rect 35544 734 35848 762
rect 36542 0 36598 800
rect 37646 0 37702 800
rect 38750 0 38806 800
rect 39854 0 39910 800
rect 40958 0 41014 800
rect 42062 0 42118 800
rect 43166 0 43222 800
rect 44270 0 44326 800
rect 45374 0 45430 800
rect 46478 0 46534 800
rect 47582 0 47638 800
rect 48686 0 48742 800
rect 49790 0 49846 800
rect 50894 0 50950 800
rect 51998 0 52054 800
rect 53102 0 53158 800
rect 54206 0 54262 800
rect 55310 0 55366 800
rect 56414 0 56470 800
rect 57518 0 57574 800
<< via2 >>
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 1674 55664 1730 55720
rect 3146 55664 3202 55720
rect 1674 54848 1730 54904
rect 1674 54052 1730 54088
rect 1674 54032 1676 54052
rect 1676 54032 1728 54052
rect 1728 54032 1730 54052
rect 1674 53216 1730 53272
rect 1674 52400 1730 52456
rect 1674 51584 1730 51640
rect 1674 50788 1730 50824
rect 1674 50768 1676 50788
rect 1676 50768 1728 50788
rect 1728 50768 1730 50788
rect 1674 49952 1730 50008
rect 1674 49136 1730 49192
rect 1674 48320 1730 48376
rect 1674 47524 1730 47560
rect 1674 47504 1676 47524
rect 1676 47504 1728 47524
rect 1728 47504 1730 47524
rect 1674 46688 1730 46744
rect 1674 45872 1730 45928
rect 1674 45056 1730 45112
rect 1674 44260 1730 44296
rect 1674 44240 1676 44260
rect 1676 44240 1728 44260
rect 1728 44240 1730 44260
rect 1674 43424 1730 43480
rect 1674 42608 1730 42664
rect 1674 41792 1730 41848
rect 1674 40996 1730 41032
rect 1674 40976 1676 40996
rect 1676 40976 1728 40996
rect 1728 40976 1730 40996
rect 1674 40160 1730 40216
rect 1674 39344 1730 39400
rect 1674 38528 1730 38584
rect 1674 37732 1730 37768
rect 1674 37712 1676 37732
rect 1676 37712 1728 37732
rect 1728 37712 1730 37732
rect 1674 36896 1730 36952
rect 1674 36080 1730 36136
rect 1674 35264 1730 35320
rect 1674 34468 1730 34504
rect 1674 34448 1676 34468
rect 1676 34448 1728 34468
rect 1728 34448 1730 34468
rect 1674 33632 1730 33688
rect 1674 32816 1730 32872
rect 1674 32000 1730 32056
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 1674 31204 1730 31240
rect 1674 31184 1676 31204
rect 1676 31184 1728 31204
rect 1728 31184 1730 31204
rect 1674 30368 1730 30424
rect 1674 29552 1730 29608
rect 1674 28736 1730 28792
rect 1674 27940 1730 27976
rect 1674 27920 1676 27940
rect 1676 27920 1728 27940
rect 1728 27920 1730 27940
rect 1674 27104 1730 27160
rect 1674 26288 1730 26344
rect 1674 25492 1730 25528
rect 1674 25472 1676 25492
rect 1676 25472 1728 25492
rect 1728 25472 1730 25492
rect 1674 24676 1730 24712
rect 1674 24656 1676 24676
rect 1676 24656 1728 24676
rect 1728 24656 1730 24676
rect 1674 23840 1730 23896
rect 1674 23024 1730 23080
rect 1674 22228 1730 22264
rect 1674 22208 1676 22228
rect 1676 22208 1728 22228
rect 1728 22208 1730 22228
rect 1674 21392 1730 21448
rect 1674 20596 1730 20632
rect 1674 20576 1676 20596
rect 1676 20576 1728 20596
rect 1728 20576 1730 20596
rect 1674 19760 1730 19816
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 24214 56364 24270 56400
rect 24214 56344 24216 56364
rect 24216 56344 24268 56364
rect 24268 56344 24270 56364
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 1674 18964 1730 19000
rect 1674 18944 1676 18964
rect 1676 18944 1728 18964
rect 1728 18944 1730 18964
rect 1674 18128 1730 18184
rect 1674 16496 1730 16552
rect 1674 15680 1730 15736
rect 1674 14864 1730 14920
rect 1674 13232 1730 13288
rect 2410 17312 2466 17368
rect 2410 14048 2466 14104
rect 1674 12416 1730 12472
rect 1674 11620 1730 11656
rect 1674 11600 1676 11620
rect 1676 11600 1728 11620
rect 1728 11600 1730 11620
rect 1674 10784 1730 10840
rect 1674 9968 1730 10024
rect 1674 9172 1730 9208
rect 1674 9152 1676 9172
rect 1676 9152 1728 9172
rect 1728 9152 1730 9172
rect 1674 8336 1730 8392
rect 1674 6704 1730 6760
rect 1674 5908 1730 5944
rect 1674 5888 1676 5908
rect 1676 5888 1728 5908
rect 1728 5888 1730 5908
rect 1674 5092 1730 5128
rect 1674 5072 1676 5092
rect 1676 5072 1728 5092
rect 1728 5072 1730 5092
rect 1674 4256 1730 4312
rect 2410 7520 2466 7576
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4710 16496 4766 16552
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4986 16496 5042 16552
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 25778 56364 25834 56400
rect 25778 56344 25780 56364
rect 25780 56344 25832 56364
rect 25832 56344 25834 56364
rect 26422 56364 26478 56400
rect 26422 56344 26424 56364
rect 26424 56344 26476 56364
rect 26476 56344 26478 56364
rect 27434 56344 27490 56400
rect 26882 55936 26938 55992
rect 26974 55700 26976 55720
rect 26976 55700 27028 55720
rect 27028 55700 27030 55720
rect 26974 55664 27030 55700
rect 28998 56370 29054 56400
rect 28998 56344 29006 56370
rect 29006 56344 29054 56370
rect 28354 55684 28410 55720
rect 28354 55664 28356 55684
rect 28356 55664 28408 55684
rect 28408 55664 28410 55684
rect 27526 55528 27582 55584
rect 28630 56228 28686 56264
rect 28630 56208 28632 56228
rect 28632 56208 28684 56228
rect 28684 56208 28686 56228
rect 28906 55956 28962 55992
rect 28906 55936 28908 55956
rect 28908 55936 28960 55956
rect 28960 55936 28962 55956
rect 28814 55564 28816 55584
rect 28816 55564 28868 55584
rect 28868 55564 28870 55584
rect 28814 55528 28870 55564
rect 30654 55664 30710 55720
rect 32586 56208 32642 56264
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 35162 56344 35218 56400
rect 35530 56364 35586 56400
rect 35530 56344 35532 56364
rect 35532 56344 35584 56364
rect 35584 56344 35586 56364
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 36174 56364 36230 56400
rect 36174 56344 36176 56364
rect 36176 56344 36228 56364
rect 36228 56344 36230 56364
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 38750 55800 38806 55856
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 57518 58928 57574 58984
rect 38750 55678 38752 55720
rect 38752 55678 38804 55720
rect 38804 55678 38806 55720
rect 38750 55664 38806 55678
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 57058 57296 57114 57352
rect 58438 58112 58494 58168
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 57058 38548 57114 38584
rect 57058 38528 57060 38548
rect 57060 38528 57112 38548
rect 57112 38528 57114 38548
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 57150 28736 57206 28792
rect 58346 56480 58402 56536
rect 57886 54848 57942 54904
rect 57886 39344 57942 39400
rect 58346 55700 58348 55720
rect 58348 55700 58400 55720
rect 58400 55700 58402 55720
rect 58346 55664 58402 55700
rect 58346 54032 58402 54088
rect 58346 53216 58402 53272
rect 58346 52436 58348 52456
rect 58348 52436 58400 52456
rect 58400 52436 58402 52456
rect 58346 52400 58402 52436
rect 58346 51584 58402 51640
rect 58346 50768 58402 50824
rect 58346 49952 58402 50008
rect 58346 49172 58348 49192
rect 58348 49172 58400 49192
rect 58400 49172 58402 49192
rect 58346 49136 58402 49172
rect 58346 48320 58402 48376
rect 58346 47504 58402 47560
rect 58346 46688 58402 46744
rect 58346 45908 58348 45928
rect 58348 45908 58400 45928
rect 58400 45908 58402 45928
rect 58346 45872 58402 45908
rect 58346 45056 58402 45112
rect 58346 44240 58402 44296
rect 58346 43424 58402 43480
rect 58346 42644 58348 42664
rect 58348 42644 58400 42664
rect 58400 42644 58402 42664
rect 58346 42608 58402 42644
rect 58346 41792 58402 41848
rect 58346 40976 58402 41032
rect 58346 40160 58402 40216
rect 58346 38528 58402 38584
rect 58346 37712 58402 37768
rect 58346 36896 58402 36952
rect 57886 36080 57942 36136
rect 57794 32816 57850 32872
rect 58346 35264 58402 35320
rect 58346 34448 58402 34504
rect 58346 33632 58402 33688
rect 58162 31184 58218 31240
rect 58346 32000 58402 32056
rect 58438 30388 58494 30424
rect 58438 30368 58440 30388
rect 58440 30368 58492 30388
rect 58492 30368 58494 30388
rect 58438 29552 58494 29608
rect 58438 27920 58494 27976
rect 58346 27104 58402 27160
rect 58346 26324 58348 26344
rect 58348 26324 58400 26344
rect 58400 26324 58402 26344
rect 58346 26288 58402 26324
rect 58346 25472 58402 25528
rect 58346 24656 58402 24712
rect 58346 23840 58402 23896
rect 58346 23060 58348 23080
rect 58348 23060 58400 23080
rect 58400 23060 58402 23080
rect 58346 23024 58402 23060
rect 58346 22208 58402 22264
rect 58346 21392 58402 21448
rect 58346 20576 58402 20632
rect 58346 19796 58348 19816
rect 58348 19796 58400 19816
rect 58400 19796 58402 19816
rect 58346 19760 58402 19796
rect 58346 18964 58402 19000
rect 58346 18944 58348 18964
rect 58348 18944 58400 18964
rect 58400 18944 58402 18964
rect 58346 18128 58402 18184
rect 57886 13232 57942 13288
rect 57518 5888 57574 5944
rect 58346 17312 58402 17368
rect 58346 16532 58348 16552
rect 58348 16532 58400 16552
rect 58400 16532 58402 16552
rect 58346 16496 58402 16532
rect 58346 15700 58402 15736
rect 58346 15680 58348 15700
rect 58348 15680 58400 15700
rect 58400 15680 58402 15700
rect 58346 14864 58402 14920
rect 58346 14048 58402 14104
rect 58346 12416 58402 12472
rect 58346 11600 58402 11656
rect 58162 10004 58164 10024
rect 58164 10004 58216 10024
rect 58216 10004 58218 10024
rect 58162 9968 58218 10004
rect 58438 10784 58494 10840
rect 58162 9152 58218 9208
rect 58162 8336 58218 8392
rect 58346 7540 58402 7576
rect 58346 7520 58348 7540
rect 58348 7520 58400 7540
rect 58400 7520 58402 7540
rect 58346 6740 58348 6760
rect 58348 6740 58400 6760
rect 58400 6740 58402 6760
rect 58346 6704 58402 6740
rect 58346 5888 58402 5944
rect 57518 3440 57574 3496
rect 56322 2624 56378 2680
rect 56046 1808 56102 1864
rect 58346 5072 58402 5128
rect 58346 4256 58402 4312
rect 58346 992 58402 1048
<< metal3 >>
rect 57513 58986 57579 58989
rect 59200 58986 60000 59016
rect 57513 58984 60000 58986
rect 57513 58928 57518 58984
rect 57574 58928 60000 58984
rect 57513 58926 60000 58928
rect 57513 58923 57579 58926
rect 59200 58896 60000 58926
rect 58433 58170 58499 58173
rect 59200 58170 60000 58200
rect 58433 58168 60000 58170
rect 58433 58112 58438 58168
rect 58494 58112 60000 58168
rect 58433 58110 60000 58112
rect 58433 58107 58499 58110
rect 59200 58080 60000 58110
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 57053 57354 57119 57357
rect 59200 57354 60000 57384
rect 57053 57352 60000 57354
rect 57053 57296 57058 57352
rect 57114 57296 60000 57352
rect 57053 57294 60000 57296
rect 57053 57291 57119 57294
rect 59200 57264 60000 57294
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 58341 56538 58407 56541
rect 59200 56538 60000 56568
rect 58341 56536 60000 56538
rect 58341 56480 58346 56536
rect 58402 56480 60000 56536
rect 58341 56478 60000 56480
rect 58341 56475 58407 56478
rect 59200 56448 60000 56478
rect 24209 56402 24275 56405
rect 25773 56402 25839 56405
rect 24209 56400 25839 56402
rect 24209 56344 24214 56400
rect 24270 56344 25778 56400
rect 25834 56344 25839 56400
rect 24209 56342 25839 56344
rect 24209 56339 24275 56342
rect 25773 56339 25839 56342
rect 26417 56402 26483 56405
rect 27429 56402 27495 56405
rect 26417 56400 27495 56402
rect 26417 56344 26422 56400
rect 26478 56344 27434 56400
rect 27490 56344 27495 56400
rect 26417 56342 27495 56344
rect 26417 56339 26483 56342
rect 27429 56339 27495 56342
rect 28993 56402 29059 56405
rect 35157 56402 35223 56405
rect 28993 56400 35223 56402
rect 28993 56344 28998 56400
rect 29054 56344 35162 56400
rect 35218 56344 35223 56400
rect 28993 56342 35223 56344
rect 28993 56339 29059 56342
rect 35157 56339 35223 56342
rect 35525 56402 35591 56405
rect 36169 56402 36235 56405
rect 35525 56400 36235 56402
rect 35525 56344 35530 56400
rect 35586 56344 36174 56400
rect 36230 56344 36235 56400
rect 35525 56342 36235 56344
rect 35525 56339 35591 56342
rect 36169 56339 36235 56342
rect 28625 56266 28691 56269
rect 32581 56266 32647 56269
rect 28625 56264 32647 56266
rect 28625 56208 28630 56264
rect 28686 56208 32586 56264
rect 32642 56208 32647 56264
rect 28625 56206 32647 56208
rect 28625 56203 28691 56206
rect 32581 56203 32647 56206
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 26877 55994 26943 55997
rect 28901 55994 28967 55997
rect 26877 55992 28967 55994
rect 26877 55936 26882 55992
rect 26938 55936 28906 55992
rect 28962 55936 28967 55992
rect 26877 55934 28967 55936
rect 26877 55931 26943 55934
rect 28901 55931 28967 55934
rect 38745 55858 38811 55861
rect 38702 55856 38811 55858
rect 38702 55800 38750 55856
rect 38806 55800 38811 55856
rect 38702 55795 38811 55800
rect 0 55722 800 55752
rect 38702 55725 38762 55795
rect 1669 55722 1735 55725
rect 0 55720 1735 55722
rect 0 55664 1674 55720
rect 1730 55664 1735 55720
rect 0 55662 1735 55664
rect 0 55632 800 55662
rect 1669 55659 1735 55662
rect 3141 55722 3207 55725
rect 26969 55722 27035 55725
rect 3141 55720 27035 55722
rect 3141 55664 3146 55720
rect 3202 55664 26974 55720
rect 27030 55664 27035 55720
rect 3141 55662 27035 55664
rect 3141 55659 3207 55662
rect 26969 55659 27035 55662
rect 28349 55722 28415 55725
rect 30649 55722 30715 55725
rect 28349 55720 30715 55722
rect 28349 55664 28354 55720
rect 28410 55664 30654 55720
rect 30710 55664 30715 55720
rect 28349 55662 30715 55664
rect 38702 55720 38811 55725
rect 38702 55664 38750 55720
rect 38806 55664 38811 55720
rect 38702 55662 38811 55664
rect 28349 55659 28415 55662
rect 30649 55659 30715 55662
rect 38745 55659 38811 55662
rect 58341 55722 58407 55725
rect 59200 55722 60000 55752
rect 58341 55720 60000 55722
rect 58341 55664 58346 55720
rect 58402 55664 60000 55720
rect 58341 55662 60000 55664
rect 58341 55659 58407 55662
rect 59200 55632 60000 55662
rect 27521 55586 27587 55589
rect 28809 55586 28875 55589
rect 27521 55584 28875 55586
rect 27521 55528 27526 55584
rect 27582 55528 28814 55584
rect 28870 55528 28875 55584
rect 27521 55526 28875 55528
rect 27521 55523 27587 55526
rect 28809 55523 28875 55526
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 0 54906 800 54936
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 1669 54906 1735 54909
rect 0 54904 1735 54906
rect 0 54848 1674 54904
rect 1730 54848 1735 54904
rect 0 54846 1735 54848
rect 0 54816 800 54846
rect 1669 54843 1735 54846
rect 57881 54906 57947 54909
rect 59200 54906 60000 54936
rect 57881 54904 60000 54906
rect 57881 54848 57886 54904
rect 57942 54848 60000 54904
rect 57881 54846 60000 54848
rect 57881 54843 57947 54846
rect 59200 54816 60000 54846
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 0 54090 800 54120
rect 1669 54090 1735 54093
rect 0 54088 1735 54090
rect 0 54032 1674 54088
rect 1730 54032 1735 54088
rect 0 54030 1735 54032
rect 0 54000 800 54030
rect 1669 54027 1735 54030
rect 58341 54090 58407 54093
rect 59200 54090 60000 54120
rect 58341 54088 60000 54090
rect 58341 54032 58346 54088
rect 58402 54032 60000 54088
rect 58341 54030 60000 54032
rect 58341 54027 58407 54030
rect 59200 54000 60000 54030
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 0 53274 800 53304
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 1669 53274 1735 53277
rect 0 53272 1735 53274
rect 0 53216 1674 53272
rect 1730 53216 1735 53272
rect 0 53214 1735 53216
rect 0 53184 800 53214
rect 1669 53211 1735 53214
rect 58341 53274 58407 53277
rect 59200 53274 60000 53304
rect 58341 53272 60000 53274
rect 58341 53216 58346 53272
rect 58402 53216 60000 53272
rect 58341 53214 60000 53216
rect 58341 53211 58407 53214
rect 59200 53184 60000 53214
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 0 52458 800 52488
rect 1669 52458 1735 52461
rect 0 52456 1735 52458
rect 0 52400 1674 52456
rect 1730 52400 1735 52456
rect 0 52398 1735 52400
rect 0 52368 800 52398
rect 1669 52395 1735 52398
rect 58341 52458 58407 52461
rect 59200 52458 60000 52488
rect 58341 52456 60000 52458
rect 58341 52400 58346 52456
rect 58402 52400 60000 52456
rect 58341 52398 60000 52400
rect 58341 52395 58407 52398
rect 59200 52368 60000 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51642 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 1669 51642 1735 51645
rect 0 51640 1735 51642
rect 0 51584 1674 51640
rect 1730 51584 1735 51640
rect 0 51582 1735 51584
rect 0 51552 800 51582
rect 1669 51579 1735 51582
rect 58341 51642 58407 51645
rect 59200 51642 60000 51672
rect 58341 51640 60000 51642
rect 58341 51584 58346 51640
rect 58402 51584 60000 51640
rect 58341 51582 60000 51584
rect 58341 51579 58407 51582
rect 59200 51552 60000 51582
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 0 50826 800 50856
rect 1669 50826 1735 50829
rect 0 50824 1735 50826
rect 0 50768 1674 50824
rect 1730 50768 1735 50824
rect 0 50766 1735 50768
rect 0 50736 800 50766
rect 1669 50763 1735 50766
rect 58341 50826 58407 50829
rect 59200 50826 60000 50856
rect 58341 50824 60000 50826
rect 58341 50768 58346 50824
rect 58402 50768 60000 50824
rect 58341 50766 60000 50768
rect 58341 50763 58407 50766
rect 59200 50736 60000 50766
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 0 50010 800 50040
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 1669 50010 1735 50013
rect 0 50008 1735 50010
rect 0 49952 1674 50008
rect 1730 49952 1735 50008
rect 0 49950 1735 49952
rect 0 49920 800 49950
rect 1669 49947 1735 49950
rect 58341 50010 58407 50013
rect 59200 50010 60000 50040
rect 58341 50008 60000 50010
rect 58341 49952 58346 50008
rect 58402 49952 60000 50008
rect 58341 49950 60000 49952
rect 58341 49947 58407 49950
rect 59200 49920 60000 49950
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 0 49194 800 49224
rect 1669 49194 1735 49197
rect 0 49192 1735 49194
rect 0 49136 1674 49192
rect 1730 49136 1735 49192
rect 0 49134 1735 49136
rect 0 49104 800 49134
rect 1669 49131 1735 49134
rect 58341 49194 58407 49197
rect 59200 49194 60000 49224
rect 58341 49192 60000 49194
rect 58341 49136 58346 49192
rect 58402 49136 60000 49192
rect 58341 49134 60000 49136
rect 58341 49131 58407 49134
rect 59200 49104 60000 49134
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 0 48378 800 48408
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 1669 48378 1735 48381
rect 0 48376 1735 48378
rect 0 48320 1674 48376
rect 1730 48320 1735 48376
rect 0 48318 1735 48320
rect 0 48288 800 48318
rect 1669 48315 1735 48318
rect 58341 48378 58407 48381
rect 59200 48378 60000 48408
rect 58341 48376 60000 48378
rect 58341 48320 58346 48376
rect 58402 48320 60000 48376
rect 58341 48318 60000 48320
rect 58341 48315 58407 48318
rect 59200 48288 60000 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 0 47562 800 47592
rect 1669 47562 1735 47565
rect 0 47560 1735 47562
rect 0 47504 1674 47560
rect 1730 47504 1735 47560
rect 0 47502 1735 47504
rect 0 47472 800 47502
rect 1669 47499 1735 47502
rect 58341 47562 58407 47565
rect 59200 47562 60000 47592
rect 58341 47560 60000 47562
rect 58341 47504 58346 47560
rect 58402 47504 60000 47560
rect 58341 47502 60000 47504
rect 58341 47499 58407 47502
rect 59200 47472 60000 47502
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 0 46746 800 46776
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 1669 46746 1735 46749
rect 0 46744 1735 46746
rect 0 46688 1674 46744
rect 1730 46688 1735 46744
rect 0 46686 1735 46688
rect 0 46656 800 46686
rect 1669 46683 1735 46686
rect 58341 46746 58407 46749
rect 59200 46746 60000 46776
rect 58341 46744 60000 46746
rect 58341 46688 58346 46744
rect 58402 46688 60000 46744
rect 58341 46686 60000 46688
rect 58341 46683 58407 46686
rect 59200 46656 60000 46686
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 0 45930 800 45960
rect 1669 45930 1735 45933
rect 0 45928 1735 45930
rect 0 45872 1674 45928
rect 1730 45872 1735 45928
rect 0 45870 1735 45872
rect 0 45840 800 45870
rect 1669 45867 1735 45870
rect 58341 45930 58407 45933
rect 59200 45930 60000 45960
rect 58341 45928 60000 45930
rect 58341 45872 58346 45928
rect 58402 45872 60000 45928
rect 58341 45870 60000 45872
rect 58341 45867 58407 45870
rect 59200 45840 60000 45870
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 0 45114 800 45144
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 1669 45114 1735 45117
rect 0 45112 1735 45114
rect 0 45056 1674 45112
rect 1730 45056 1735 45112
rect 0 45054 1735 45056
rect 0 45024 800 45054
rect 1669 45051 1735 45054
rect 58341 45114 58407 45117
rect 59200 45114 60000 45144
rect 58341 45112 60000 45114
rect 58341 45056 58346 45112
rect 58402 45056 60000 45112
rect 58341 45054 60000 45056
rect 58341 45051 58407 45054
rect 59200 45024 60000 45054
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 0 44298 800 44328
rect 1669 44298 1735 44301
rect 0 44296 1735 44298
rect 0 44240 1674 44296
rect 1730 44240 1735 44296
rect 0 44238 1735 44240
rect 0 44208 800 44238
rect 1669 44235 1735 44238
rect 58341 44298 58407 44301
rect 59200 44298 60000 44328
rect 58341 44296 60000 44298
rect 58341 44240 58346 44296
rect 58402 44240 60000 44296
rect 58341 44238 60000 44240
rect 58341 44235 58407 44238
rect 59200 44208 60000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 0 43482 800 43512
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 1669 43482 1735 43485
rect 0 43480 1735 43482
rect 0 43424 1674 43480
rect 1730 43424 1735 43480
rect 0 43422 1735 43424
rect 0 43392 800 43422
rect 1669 43419 1735 43422
rect 58341 43482 58407 43485
rect 59200 43482 60000 43512
rect 58341 43480 60000 43482
rect 58341 43424 58346 43480
rect 58402 43424 60000 43480
rect 58341 43422 60000 43424
rect 58341 43419 58407 43422
rect 59200 43392 60000 43422
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 0 42666 800 42696
rect 1669 42666 1735 42669
rect 0 42664 1735 42666
rect 0 42608 1674 42664
rect 1730 42608 1735 42664
rect 0 42606 1735 42608
rect 0 42576 800 42606
rect 1669 42603 1735 42606
rect 58341 42666 58407 42669
rect 59200 42666 60000 42696
rect 58341 42664 60000 42666
rect 58341 42608 58346 42664
rect 58402 42608 60000 42664
rect 58341 42606 60000 42608
rect 58341 42603 58407 42606
rect 59200 42576 60000 42606
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 0 41850 800 41880
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 1669 41850 1735 41853
rect 0 41848 1735 41850
rect 0 41792 1674 41848
rect 1730 41792 1735 41848
rect 0 41790 1735 41792
rect 0 41760 800 41790
rect 1669 41787 1735 41790
rect 58341 41850 58407 41853
rect 59200 41850 60000 41880
rect 58341 41848 60000 41850
rect 58341 41792 58346 41848
rect 58402 41792 60000 41848
rect 58341 41790 60000 41792
rect 58341 41787 58407 41790
rect 59200 41760 60000 41790
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41034 800 41064
rect 1669 41034 1735 41037
rect 0 41032 1735 41034
rect 0 40976 1674 41032
rect 1730 40976 1735 41032
rect 0 40974 1735 40976
rect 0 40944 800 40974
rect 1669 40971 1735 40974
rect 58341 41034 58407 41037
rect 59200 41034 60000 41064
rect 58341 41032 60000 41034
rect 58341 40976 58346 41032
rect 58402 40976 60000 41032
rect 58341 40974 60000 40976
rect 58341 40971 58407 40974
rect 59200 40944 60000 40974
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 0 40218 800 40248
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 1669 40218 1735 40221
rect 0 40216 1735 40218
rect 0 40160 1674 40216
rect 1730 40160 1735 40216
rect 0 40158 1735 40160
rect 0 40128 800 40158
rect 1669 40155 1735 40158
rect 58341 40218 58407 40221
rect 59200 40218 60000 40248
rect 58341 40216 60000 40218
rect 58341 40160 58346 40216
rect 58402 40160 60000 40216
rect 58341 40158 60000 40160
rect 58341 40155 58407 40158
rect 59200 40128 60000 40158
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39402 800 39432
rect 1669 39402 1735 39405
rect 0 39400 1735 39402
rect 0 39344 1674 39400
rect 1730 39344 1735 39400
rect 0 39342 1735 39344
rect 0 39312 800 39342
rect 1669 39339 1735 39342
rect 57881 39402 57947 39405
rect 59200 39402 60000 39432
rect 57881 39400 60000 39402
rect 57881 39344 57886 39400
rect 57942 39344 60000 39400
rect 57881 39342 60000 39344
rect 57881 39339 57947 39342
rect 59200 39312 60000 39342
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 0 38586 800 38616
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 1669 38586 1735 38589
rect 0 38584 1735 38586
rect 0 38528 1674 38584
rect 1730 38528 1735 38584
rect 0 38526 1735 38528
rect 0 38496 800 38526
rect 1669 38523 1735 38526
rect 57053 38586 57119 38589
rect 58341 38586 58407 38589
rect 59200 38586 60000 38616
rect 57053 38584 60000 38586
rect 57053 38528 57058 38584
rect 57114 38528 58346 38584
rect 58402 38528 60000 38584
rect 57053 38526 60000 38528
rect 57053 38523 57119 38526
rect 58341 38523 58407 38526
rect 59200 38496 60000 38526
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 0 37770 800 37800
rect 1669 37770 1735 37773
rect 0 37768 1735 37770
rect 0 37712 1674 37768
rect 1730 37712 1735 37768
rect 0 37710 1735 37712
rect 0 37680 800 37710
rect 1669 37707 1735 37710
rect 58341 37770 58407 37773
rect 59200 37770 60000 37800
rect 58341 37768 60000 37770
rect 58341 37712 58346 37768
rect 58402 37712 60000 37768
rect 58341 37710 60000 37712
rect 58341 37707 58407 37710
rect 59200 37680 60000 37710
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 0 36954 800 36984
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 1669 36954 1735 36957
rect 0 36952 1735 36954
rect 0 36896 1674 36952
rect 1730 36896 1735 36952
rect 0 36894 1735 36896
rect 0 36864 800 36894
rect 1669 36891 1735 36894
rect 58341 36954 58407 36957
rect 59200 36954 60000 36984
rect 58341 36952 60000 36954
rect 58341 36896 58346 36952
rect 58402 36896 60000 36952
rect 58341 36894 60000 36896
rect 58341 36891 58407 36894
rect 59200 36864 60000 36894
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 36138 800 36168
rect 1669 36138 1735 36141
rect 0 36136 1735 36138
rect 0 36080 1674 36136
rect 1730 36080 1735 36136
rect 0 36078 1735 36080
rect 0 36048 800 36078
rect 1669 36075 1735 36078
rect 57881 36138 57947 36141
rect 59200 36138 60000 36168
rect 57881 36136 60000 36138
rect 57881 36080 57886 36136
rect 57942 36080 60000 36136
rect 57881 36078 60000 36080
rect 57881 36075 57947 36078
rect 59200 36048 60000 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 0 35322 800 35352
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 1669 35322 1735 35325
rect 0 35320 1735 35322
rect 0 35264 1674 35320
rect 1730 35264 1735 35320
rect 0 35262 1735 35264
rect 0 35232 800 35262
rect 1669 35259 1735 35262
rect 58341 35322 58407 35325
rect 59200 35322 60000 35352
rect 58341 35320 60000 35322
rect 58341 35264 58346 35320
rect 58402 35264 60000 35320
rect 58341 35262 60000 35264
rect 58341 35259 58407 35262
rect 59200 35232 60000 35262
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 0 34506 800 34536
rect 1669 34506 1735 34509
rect 0 34504 1735 34506
rect 0 34448 1674 34504
rect 1730 34448 1735 34504
rect 0 34446 1735 34448
rect 0 34416 800 34446
rect 1669 34443 1735 34446
rect 58341 34506 58407 34509
rect 59200 34506 60000 34536
rect 58341 34504 60000 34506
rect 58341 34448 58346 34504
rect 58402 34448 60000 34504
rect 58341 34446 60000 34448
rect 58341 34443 58407 34446
rect 59200 34416 60000 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 0 33690 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 1669 33690 1735 33693
rect 0 33688 1735 33690
rect 0 33632 1674 33688
rect 1730 33632 1735 33688
rect 0 33630 1735 33632
rect 0 33600 800 33630
rect 1669 33627 1735 33630
rect 58341 33690 58407 33693
rect 59200 33690 60000 33720
rect 58341 33688 60000 33690
rect 58341 33632 58346 33688
rect 58402 33632 60000 33688
rect 58341 33630 60000 33632
rect 58341 33627 58407 33630
rect 59200 33600 60000 33630
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 0 32874 800 32904
rect 1669 32874 1735 32877
rect 0 32872 1735 32874
rect 0 32816 1674 32872
rect 1730 32816 1735 32872
rect 0 32814 1735 32816
rect 0 32784 800 32814
rect 1669 32811 1735 32814
rect 57789 32874 57855 32877
rect 59200 32874 60000 32904
rect 57789 32872 60000 32874
rect 57789 32816 57794 32872
rect 57850 32816 60000 32872
rect 57789 32814 60000 32816
rect 57789 32811 57855 32814
rect 59200 32784 60000 32814
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1669 32058 1735 32061
rect 0 32056 1735 32058
rect 0 32000 1674 32056
rect 1730 32000 1735 32056
rect 0 31998 1735 32000
rect 0 31968 800 31998
rect 1669 31995 1735 31998
rect 58341 32058 58407 32061
rect 59200 32058 60000 32088
rect 58341 32056 60000 32058
rect 58341 32000 58346 32056
rect 58402 32000 60000 32056
rect 58341 31998 60000 32000
rect 58341 31995 58407 31998
rect 59200 31968 60000 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 0 31242 800 31272
rect 1669 31242 1735 31245
rect 0 31240 1735 31242
rect 0 31184 1674 31240
rect 1730 31184 1735 31240
rect 0 31182 1735 31184
rect 0 31152 800 31182
rect 1669 31179 1735 31182
rect 58157 31242 58223 31245
rect 59200 31242 60000 31272
rect 58157 31240 60000 31242
rect 58157 31184 58162 31240
rect 58218 31184 60000 31240
rect 58157 31182 60000 31184
rect 58157 31179 58223 31182
rect 59200 31152 60000 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 0 30426 800 30456
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 1669 30426 1735 30429
rect 0 30424 1735 30426
rect 0 30368 1674 30424
rect 1730 30368 1735 30424
rect 0 30366 1735 30368
rect 0 30336 800 30366
rect 1669 30363 1735 30366
rect 58433 30426 58499 30429
rect 59200 30426 60000 30456
rect 58433 30424 60000 30426
rect 58433 30368 58438 30424
rect 58494 30368 60000 30424
rect 58433 30366 60000 30368
rect 58433 30363 58499 30366
rect 59200 30336 60000 30366
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 0 29610 800 29640
rect 1669 29610 1735 29613
rect 0 29608 1735 29610
rect 0 29552 1674 29608
rect 1730 29552 1735 29608
rect 0 29550 1735 29552
rect 0 29520 800 29550
rect 1669 29547 1735 29550
rect 58433 29610 58499 29613
rect 59200 29610 60000 29640
rect 58433 29608 60000 29610
rect 58433 29552 58438 29608
rect 58494 29552 60000 29608
rect 58433 29550 60000 29552
rect 58433 29547 58499 29550
rect 59200 29520 60000 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 0 28794 800 28824
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 1669 28794 1735 28797
rect 0 28792 1735 28794
rect 0 28736 1674 28792
rect 1730 28736 1735 28792
rect 0 28734 1735 28736
rect 0 28704 800 28734
rect 1669 28731 1735 28734
rect 57145 28794 57211 28797
rect 59200 28794 60000 28824
rect 57145 28792 60000 28794
rect 57145 28736 57150 28792
rect 57206 28736 60000 28792
rect 57145 28734 60000 28736
rect 57145 28731 57211 28734
rect 59200 28704 60000 28734
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 0 27978 800 28008
rect 1669 27978 1735 27981
rect 0 27976 1735 27978
rect 0 27920 1674 27976
rect 1730 27920 1735 27976
rect 0 27918 1735 27920
rect 0 27888 800 27918
rect 1669 27915 1735 27918
rect 58433 27978 58499 27981
rect 59200 27978 60000 28008
rect 58433 27976 60000 27978
rect 58433 27920 58438 27976
rect 58494 27920 60000 27976
rect 58433 27918 60000 27920
rect 58433 27915 58499 27918
rect 59200 27888 60000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 0 27162 800 27192
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 1669 27162 1735 27165
rect 0 27160 1735 27162
rect 0 27104 1674 27160
rect 1730 27104 1735 27160
rect 0 27102 1735 27104
rect 0 27072 800 27102
rect 1669 27099 1735 27102
rect 58341 27162 58407 27165
rect 59200 27162 60000 27192
rect 58341 27160 60000 27162
rect 58341 27104 58346 27160
rect 58402 27104 60000 27160
rect 58341 27102 60000 27104
rect 58341 27099 58407 27102
rect 59200 27072 60000 27102
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 0 26346 800 26376
rect 1669 26346 1735 26349
rect 0 26344 1735 26346
rect 0 26288 1674 26344
rect 1730 26288 1735 26344
rect 0 26286 1735 26288
rect 0 26256 800 26286
rect 1669 26283 1735 26286
rect 58341 26346 58407 26349
rect 59200 26346 60000 26376
rect 58341 26344 60000 26346
rect 58341 26288 58346 26344
rect 58402 26288 60000 26344
rect 58341 26286 60000 26288
rect 58341 26283 58407 26286
rect 59200 26256 60000 26286
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 0 25530 800 25560
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 1669 25530 1735 25533
rect 0 25528 1735 25530
rect 0 25472 1674 25528
rect 1730 25472 1735 25528
rect 0 25470 1735 25472
rect 0 25440 800 25470
rect 1669 25467 1735 25470
rect 58341 25530 58407 25533
rect 59200 25530 60000 25560
rect 58341 25528 60000 25530
rect 58341 25472 58346 25528
rect 58402 25472 60000 25528
rect 58341 25470 60000 25472
rect 58341 25467 58407 25470
rect 59200 25440 60000 25470
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 0 24714 800 24744
rect 1669 24714 1735 24717
rect 0 24712 1735 24714
rect 0 24656 1674 24712
rect 1730 24656 1735 24712
rect 0 24654 1735 24656
rect 0 24624 800 24654
rect 1669 24651 1735 24654
rect 58341 24714 58407 24717
rect 59200 24714 60000 24744
rect 58341 24712 60000 24714
rect 58341 24656 58346 24712
rect 58402 24656 60000 24712
rect 58341 24654 60000 24656
rect 58341 24651 58407 24654
rect 59200 24624 60000 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 0 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 1669 23898 1735 23901
rect 0 23896 1735 23898
rect 0 23840 1674 23896
rect 1730 23840 1735 23896
rect 0 23838 1735 23840
rect 0 23808 800 23838
rect 1669 23835 1735 23838
rect 58341 23898 58407 23901
rect 59200 23898 60000 23928
rect 58341 23896 60000 23898
rect 58341 23840 58346 23896
rect 58402 23840 60000 23896
rect 58341 23838 60000 23840
rect 58341 23835 58407 23838
rect 59200 23808 60000 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23082 800 23112
rect 1669 23082 1735 23085
rect 0 23080 1735 23082
rect 0 23024 1674 23080
rect 1730 23024 1735 23080
rect 0 23022 1735 23024
rect 0 22992 800 23022
rect 1669 23019 1735 23022
rect 58341 23082 58407 23085
rect 59200 23082 60000 23112
rect 58341 23080 60000 23082
rect 58341 23024 58346 23080
rect 58402 23024 60000 23080
rect 58341 23022 60000 23024
rect 58341 23019 58407 23022
rect 59200 22992 60000 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4210 22336 4526 22337
rect 0 22266 800 22296
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 1669 22266 1735 22269
rect 0 22264 1735 22266
rect 0 22208 1674 22264
rect 1730 22208 1735 22264
rect 0 22206 1735 22208
rect 0 22176 800 22206
rect 1669 22203 1735 22206
rect 58341 22266 58407 22269
rect 59200 22266 60000 22296
rect 58341 22264 60000 22266
rect 58341 22208 58346 22264
rect 58402 22208 60000 22264
rect 58341 22206 60000 22208
rect 58341 22203 58407 22206
rect 59200 22176 60000 22206
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 0 21450 800 21480
rect 1669 21450 1735 21453
rect 0 21448 1735 21450
rect 0 21392 1674 21448
rect 1730 21392 1735 21448
rect 0 21390 1735 21392
rect 0 21360 800 21390
rect 1669 21387 1735 21390
rect 58341 21450 58407 21453
rect 59200 21450 60000 21480
rect 58341 21448 60000 21450
rect 58341 21392 58346 21448
rect 58402 21392 60000 21448
rect 58341 21390 60000 21392
rect 58341 21387 58407 21390
rect 59200 21360 60000 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 0 20634 800 20664
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 1669 20634 1735 20637
rect 0 20632 1735 20634
rect 0 20576 1674 20632
rect 1730 20576 1735 20632
rect 0 20574 1735 20576
rect 0 20544 800 20574
rect 1669 20571 1735 20574
rect 58341 20634 58407 20637
rect 59200 20634 60000 20664
rect 58341 20632 60000 20634
rect 58341 20576 58346 20632
rect 58402 20576 60000 20632
rect 58341 20574 60000 20576
rect 58341 20571 58407 20574
rect 59200 20544 60000 20574
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 0 19818 800 19848
rect 1669 19818 1735 19821
rect 0 19816 1735 19818
rect 0 19760 1674 19816
rect 1730 19760 1735 19816
rect 0 19758 1735 19760
rect 0 19728 800 19758
rect 1669 19755 1735 19758
rect 58341 19818 58407 19821
rect 59200 19818 60000 19848
rect 58341 19816 60000 19818
rect 58341 19760 58346 19816
rect 58402 19760 60000 19816
rect 58341 19758 60000 19760
rect 58341 19755 58407 19758
rect 59200 19728 60000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 0 19002 800 19032
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 1669 19002 1735 19005
rect 0 19000 1735 19002
rect 0 18944 1674 19000
rect 1730 18944 1735 19000
rect 0 18942 1735 18944
rect 0 18912 800 18942
rect 1669 18939 1735 18942
rect 58341 19002 58407 19005
rect 59200 19002 60000 19032
rect 58341 19000 60000 19002
rect 58341 18944 58346 19000
rect 58402 18944 60000 19000
rect 58341 18942 60000 18944
rect 58341 18939 58407 18942
rect 59200 18912 60000 18942
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 0 18186 800 18216
rect 1669 18186 1735 18189
rect 0 18184 1735 18186
rect 0 18128 1674 18184
rect 1730 18128 1735 18184
rect 0 18126 1735 18128
rect 0 18096 800 18126
rect 1669 18123 1735 18126
rect 58341 18186 58407 18189
rect 59200 18186 60000 18216
rect 58341 18184 60000 18186
rect 58341 18128 58346 18184
rect 58402 18128 60000 18184
rect 58341 18126 60000 18128
rect 58341 18123 58407 18126
rect 59200 18096 60000 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 0 17370 800 17400
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 2405 17370 2471 17373
rect 0 17368 2471 17370
rect 0 17312 2410 17368
rect 2466 17312 2471 17368
rect 0 17310 2471 17312
rect 0 17280 800 17310
rect 2405 17307 2471 17310
rect 58341 17370 58407 17373
rect 59200 17370 60000 17400
rect 58341 17368 60000 17370
rect 58341 17312 58346 17368
rect 58402 17312 60000 17368
rect 58341 17310 60000 17312
rect 58341 17307 58407 17310
rect 59200 17280 60000 17310
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 0 16554 800 16584
rect 1669 16554 1735 16557
rect 0 16552 1735 16554
rect 0 16496 1674 16552
rect 1730 16496 1735 16552
rect 0 16494 1735 16496
rect 0 16464 800 16494
rect 1669 16491 1735 16494
rect 4705 16554 4771 16557
rect 4981 16554 5047 16557
rect 4705 16552 5047 16554
rect 4705 16496 4710 16552
rect 4766 16496 4986 16552
rect 5042 16496 5047 16552
rect 4705 16494 5047 16496
rect 4705 16491 4771 16494
rect 4981 16491 5047 16494
rect 58341 16554 58407 16557
rect 59200 16554 60000 16584
rect 58341 16552 60000 16554
rect 58341 16496 58346 16552
rect 58402 16496 60000 16552
rect 58341 16494 60000 16496
rect 58341 16491 58407 16494
rect 59200 16464 60000 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 0 15736 1735 15738
rect 0 15680 1674 15736
rect 1730 15680 1735 15736
rect 0 15678 1735 15680
rect 0 15648 800 15678
rect 1669 15675 1735 15678
rect 58341 15738 58407 15741
rect 59200 15738 60000 15768
rect 58341 15736 60000 15738
rect 58341 15680 58346 15736
rect 58402 15680 60000 15736
rect 58341 15678 60000 15680
rect 58341 15675 58407 15678
rect 59200 15648 60000 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 0 14922 800 14952
rect 1669 14922 1735 14925
rect 0 14920 1735 14922
rect 0 14864 1674 14920
rect 1730 14864 1735 14920
rect 0 14862 1735 14864
rect 0 14832 800 14862
rect 1669 14859 1735 14862
rect 58341 14922 58407 14925
rect 59200 14922 60000 14952
rect 58341 14920 60000 14922
rect 58341 14864 58346 14920
rect 58402 14864 60000 14920
rect 58341 14862 60000 14864
rect 58341 14859 58407 14862
rect 59200 14832 60000 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 0 14106 800 14136
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 2405 14106 2471 14109
rect 0 14104 2471 14106
rect 0 14048 2410 14104
rect 2466 14048 2471 14104
rect 0 14046 2471 14048
rect 0 14016 800 14046
rect 2405 14043 2471 14046
rect 58341 14106 58407 14109
rect 59200 14106 60000 14136
rect 58341 14104 60000 14106
rect 58341 14048 58346 14104
rect 58402 14048 60000 14104
rect 58341 14046 60000 14048
rect 58341 14043 58407 14046
rect 59200 14016 60000 14046
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 0 13290 800 13320
rect 1669 13290 1735 13293
rect 0 13288 1735 13290
rect 0 13232 1674 13288
rect 1730 13232 1735 13288
rect 0 13230 1735 13232
rect 0 13200 800 13230
rect 1669 13227 1735 13230
rect 57881 13290 57947 13293
rect 59200 13290 60000 13320
rect 57881 13288 60000 13290
rect 57881 13232 57886 13288
rect 57942 13232 60000 13288
rect 57881 13230 60000 13232
rect 57881 13227 57947 13230
rect 59200 13200 60000 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 0 12474 800 12504
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 1669 12474 1735 12477
rect 0 12472 1735 12474
rect 0 12416 1674 12472
rect 1730 12416 1735 12472
rect 0 12414 1735 12416
rect 0 12384 800 12414
rect 1669 12411 1735 12414
rect 58341 12474 58407 12477
rect 59200 12474 60000 12504
rect 58341 12472 60000 12474
rect 58341 12416 58346 12472
rect 58402 12416 60000 12472
rect 58341 12414 60000 12416
rect 58341 12411 58407 12414
rect 59200 12384 60000 12414
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 0 11658 800 11688
rect 1669 11658 1735 11661
rect 0 11656 1735 11658
rect 0 11600 1674 11656
rect 1730 11600 1735 11656
rect 0 11598 1735 11600
rect 0 11568 800 11598
rect 1669 11595 1735 11598
rect 58341 11658 58407 11661
rect 59200 11658 60000 11688
rect 58341 11656 60000 11658
rect 58341 11600 58346 11656
rect 58402 11600 60000 11656
rect 58341 11598 60000 11600
rect 58341 11595 58407 11598
rect 59200 11568 60000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 0 10842 800 10872
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 1669 10842 1735 10845
rect 0 10840 1735 10842
rect 0 10784 1674 10840
rect 1730 10784 1735 10840
rect 0 10782 1735 10784
rect 0 10752 800 10782
rect 1669 10779 1735 10782
rect 58433 10842 58499 10845
rect 59200 10842 60000 10872
rect 58433 10840 60000 10842
rect 58433 10784 58438 10840
rect 58494 10784 60000 10840
rect 58433 10782 60000 10784
rect 58433 10779 58499 10782
rect 59200 10752 60000 10782
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 0 10026 800 10056
rect 1669 10026 1735 10029
rect 0 10024 1735 10026
rect 0 9968 1674 10024
rect 1730 9968 1735 10024
rect 0 9966 1735 9968
rect 0 9936 800 9966
rect 1669 9963 1735 9966
rect 58157 10026 58223 10029
rect 59200 10026 60000 10056
rect 58157 10024 60000 10026
rect 58157 9968 58162 10024
rect 58218 9968 60000 10024
rect 58157 9966 60000 9968
rect 58157 9963 58223 9966
rect 59200 9936 60000 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 0 9210 800 9240
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 1669 9210 1735 9213
rect 0 9208 1735 9210
rect 0 9152 1674 9208
rect 1730 9152 1735 9208
rect 0 9150 1735 9152
rect 0 9120 800 9150
rect 1669 9147 1735 9150
rect 58157 9210 58223 9213
rect 59200 9210 60000 9240
rect 58157 9208 60000 9210
rect 58157 9152 58162 9208
rect 58218 9152 60000 9208
rect 58157 9150 60000 9152
rect 58157 9147 58223 9150
rect 59200 9120 60000 9150
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 0 8394 800 8424
rect 1669 8394 1735 8397
rect 0 8392 1735 8394
rect 0 8336 1674 8392
rect 1730 8336 1735 8392
rect 0 8334 1735 8336
rect 0 8304 800 8334
rect 1669 8331 1735 8334
rect 58157 8394 58223 8397
rect 59200 8394 60000 8424
rect 58157 8392 60000 8394
rect 58157 8336 58162 8392
rect 58218 8336 60000 8392
rect 58157 8334 60000 8336
rect 58157 8331 58223 8334
rect 59200 8304 60000 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 2405 7578 2471 7581
rect 0 7576 2471 7578
rect 0 7520 2410 7576
rect 2466 7520 2471 7576
rect 0 7518 2471 7520
rect 0 7488 800 7518
rect 2405 7515 2471 7518
rect 58341 7578 58407 7581
rect 59200 7578 60000 7608
rect 58341 7576 60000 7578
rect 58341 7520 58346 7576
rect 58402 7520 60000 7576
rect 58341 7518 60000 7520
rect 58341 7515 58407 7518
rect 59200 7488 60000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6762 800 6792
rect 1669 6762 1735 6765
rect 0 6760 1735 6762
rect 0 6704 1674 6760
rect 1730 6704 1735 6760
rect 0 6702 1735 6704
rect 0 6672 800 6702
rect 1669 6699 1735 6702
rect 58341 6762 58407 6765
rect 59200 6762 60000 6792
rect 58341 6760 60000 6762
rect 58341 6704 58346 6760
rect 58402 6704 60000 6760
rect 58341 6702 60000 6704
rect 58341 6699 58407 6702
rect 59200 6672 60000 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 0 5946 800 5976
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 1669 5946 1735 5949
rect 0 5944 1735 5946
rect 0 5888 1674 5944
rect 1730 5888 1735 5944
rect 0 5886 1735 5888
rect 0 5856 800 5886
rect 1669 5883 1735 5886
rect 57513 5946 57579 5949
rect 58341 5946 58407 5949
rect 59200 5946 60000 5976
rect 57513 5944 60000 5946
rect 57513 5888 57518 5944
rect 57574 5888 58346 5944
rect 58402 5888 60000 5944
rect 57513 5886 60000 5888
rect 57513 5883 57579 5886
rect 58341 5883 58407 5886
rect 59200 5856 60000 5886
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 0 5130 800 5160
rect 1669 5130 1735 5133
rect 0 5128 1735 5130
rect 0 5072 1674 5128
rect 1730 5072 1735 5128
rect 0 5070 1735 5072
rect 0 5040 800 5070
rect 1669 5067 1735 5070
rect 58341 5130 58407 5133
rect 59200 5130 60000 5160
rect 58341 5128 60000 5130
rect 58341 5072 58346 5128
rect 58402 5072 60000 5128
rect 58341 5070 60000 5072
rect 58341 5067 58407 5070
rect 59200 5040 60000 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 0 4314 800 4344
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 800 4254
rect 1669 4251 1735 4254
rect 58341 4314 58407 4317
rect 59200 4314 60000 4344
rect 58341 4312 60000 4314
rect 58341 4256 58346 4312
rect 58402 4256 60000 4312
rect 58341 4254 60000 4256
rect 58341 4251 58407 4254
rect 59200 4224 60000 4254
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 57513 3498 57579 3501
rect 59200 3498 60000 3528
rect 57513 3496 60000 3498
rect 57513 3440 57518 3496
rect 57574 3440 60000 3496
rect 57513 3438 60000 3440
rect 57513 3435 57579 3438
rect 59200 3408 60000 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 56317 2682 56383 2685
rect 59200 2682 60000 2712
rect 56317 2680 60000 2682
rect 56317 2624 56322 2680
rect 56378 2624 60000 2680
rect 56317 2622 60000 2624
rect 56317 2619 56383 2622
rect 59200 2592 60000 2622
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 56041 1866 56107 1869
rect 59200 1866 60000 1896
rect 56041 1864 60000 1866
rect 56041 1808 56046 1864
rect 56102 1808 60000 1864
rect 56041 1806 60000 1808
rect 56041 1803 56107 1806
rect 59200 1776 60000 1806
rect 58341 1050 58407 1053
rect 59200 1050 60000 1080
rect 58341 1048 60000 1050
rect 58341 992 58346 1048
rect 58402 992 60000 1048
rect 58341 990 60000 992
rect 58341 987 58407 990
rect 59200 960 60000 990
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4048 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A1
timestamp 1666464484
transform 1 0 4508 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__S
timestamp 1666464484
transform 1 0 2300 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A0
timestamp 1666464484
transform -1 0 6992 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A1
timestamp 1666464484
transform 1 0 6992 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__S
timestamp 1666464484
transform 1 0 7360 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A0
timestamp 1666464484
transform -1 0 13156 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A1
timestamp 1666464484
transform 1 0 11684 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__S
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A0
timestamp 1666464484
transform -1 0 9292 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A1
timestamp 1666464484
transform 1 0 9200 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__S
timestamp 1666464484
transform 1 0 9660 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A0
timestamp 1666464484
transform 1 0 16652 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A1
timestamp 1666464484
transform 1 0 16468 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__S
timestamp 1666464484
transform 1 0 18032 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A0
timestamp 1666464484
transform 1 0 18400 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A1
timestamp 1666464484
transform 1 0 18584 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__S
timestamp 1666464484
transform 1 0 20148 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A0
timestamp 1666464484
transform 1 0 18768 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1666464484
transform 1 0 18216 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__S
timestamp 1666464484
transform 1 0 20792 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A0
timestamp 1666464484
transform 1 0 18584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1
timestamp 1666464484
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__S
timestamp 1666464484
transform 1 0 19596 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A0
timestamp 1666464484
transform -1 0 20792 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A1
timestamp 1666464484
transform 1 0 18768 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__S
timestamp 1666464484
transform -1 0 20424 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A1
timestamp 1666464484
transform -1 0 20240 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__S
timestamp 1666464484
transform 1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A1
timestamp 1666464484
transform 1 0 20976 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__S
timestamp 1666464484
transform -1 0 22908 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A1
timestamp 1666464484
transform -1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__S
timestamp 1666464484
transform 1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1666464484
transform 1 0 38180 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1666464484
transform 1 0 37536 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A
timestamp 1666464484
transform 1 0 33856 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666464484
transform 1 0 29072 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1666464484
transform 1 0 28980 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__C_N
timestamp 1666464484
transform 1 0 28796 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A
timestamp 1666464484
transform 1 0 29164 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A_N
timestamp 1666464484
transform -1 0 32476 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__B
timestamp 1666464484
transform 1 0 31832 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1666464484
transform -1 0 38548 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1666464484
transform 1 0 40572 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__B
timestamp 1666464484
transform -1 0 41216 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__C
timestamp 1666464484
transform -1 0 41768 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A_N
timestamp 1666464484
transform 1 0 40204 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__B
timestamp 1666464484
transform 1 0 39652 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__C
timestamp 1666464484
transform 1 0 39376 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A_N
timestamp 1666464484
transform -1 0 40204 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__B
timestamp 1666464484
transform -1 0 39744 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__C
timestamp 1666464484
transform 1 0 39284 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__C
timestamp 1666464484
transform 1 0 33948 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1666464484
transform 1 0 31648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1666464484
transform 1 0 22816 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A1
timestamp 1666464484
transform -1 0 27140 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A1
timestamp 1666464484
transform 1 0 23920 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A1
timestamp 1666464484
transform -1 0 26680 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A1
timestamp 1666464484
transform -1 0 29716 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A1
timestamp 1666464484
transform 1 0 36892 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A1
timestamp 1666464484
transform -1 0 31096 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1666464484
transform 1 0 56396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1666464484
transform 1 0 55568 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__S0
timestamp 1666464484
transform -1 0 57040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__S1
timestamp 1666464484
transform -1 0 56120 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__S0
timestamp 1666464484
transform 1 0 57592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__S1
timestamp 1666464484
transform 1 0 57040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__S0
timestamp 1666464484
transform 1 0 57592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__S1
timestamp 1666464484
transform 1 0 57040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A
timestamp 1666464484
transform 1 0 40020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__S0
timestamp 1666464484
transform 1 0 56856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__S1
timestamp 1666464484
transform -1 0 56120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__S0
timestamp 1666464484
transform 1 0 57408 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__S1
timestamp 1666464484
transform 1 0 56856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__S0
timestamp 1666464484
transform -1 0 58420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__S1
timestamp 1666464484
transform 1 0 57408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A3
timestamp 1666464484
transform -1 0 57776 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__S0
timestamp 1666464484
transform 1 0 57408 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__S1
timestamp 1666464484
transform 1 0 56856 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A3
timestamp 1666464484
transform -1 0 58420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__S0
timestamp 1666464484
transform 1 0 57408 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__S1
timestamp 1666464484
transform 1 0 56856 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A3
timestamp 1666464484
transform 1 0 56856 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__S0
timestamp 1666464484
transform -1 0 58420 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__S1
timestamp 1666464484
transform -1 0 57592 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1666464484
transform 1 0 46920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A3
timestamp 1666464484
transform -1 0 56120 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__S0
timestamp 1666464484
transform 1 0 57408 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__S1
timestamp 1666464484
transform 1 0 56856 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A
timestamp 1666464484
transform -1 0 55384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A3
timestamp 1666464484
transform 1 0 57408 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__S0
timestamp 1666464484
transform 1 0 56120 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__S1
timestamp 1666464484
transform 1 0 55752 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1666464484
transform 1 0 48944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A3
timestamp 1666464484
transform -1 0 57592 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__S0
timestamp 1666464484
transform 1 0 56028 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__S1
timestamp 1666464484
transform 1 0 55660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A3
timestamp 1666464484
transform 1 0 56672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__S0
timestamp 1666464484
transform 1 0 54188 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__S1
timestamp 1666464484
transform 1 0 53820 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A3
timestamp 1666464484
transform 1 0 57408 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__S0
timestamp 1666464484
transform 1 0 56120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__S1
timestamp 1666464484
transform 1 0 55752 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A3
timestamp 1666464484
transform 1 0 57408 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__S0
timestamp 1666464484
transform 1 0 56580 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__S1
timestamp 1666464484
transform 1 0 56212 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1666464484
transform 1 0 53544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A3
timestamp 1666464484
transform -1 0 56580 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__S0
timestamp 1666464484
transform 1 0 54188 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__S1
timestamp 1666464484
transform 1 0 53820 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1666464484
transform -1 0 54832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A3
timestamp 1666464484
transform -1 0 57684 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__S0
timestamp 1666464484
transform 1 0 55660 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__S1
timestamp 1666464484
transform 1 0 55292 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1666464484
transform 1 0 55752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__S0
timestamp 1666464484
transform -1 0 56580 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__S1
timestamp 1666464484
transform -1 0 56212 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1666464484
transform 1 0 56580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1666464484
transform -1 0 21804 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__B
timestamp 1666464484
transform -1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1666464484
transform -1 0 18584 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A0
timestamp 1666464484
transform -1 0 4692 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A1
timestamp 1666464484
transform 1 0 3956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__S
timestamp 1666464484
transform -1 0 3680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A0
timestamp 1666464484
transform -1 0 9292 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A1
timestamp 1666464484
transform 1 0 9568 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__S
timestamp 1666464484
transform 1 0 8464 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A0
timestamp 1666464484
transform 1 0 10120 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A1
timestamp 1666464484
transform 1 0 10304 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__S
timestamp 1666464484
transform 1 0 10672 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A0
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A1
timestamp 1666464484
transform 1 0 3956 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__S
timestamp 1666464484
transform 1 0 3404 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A0
timestamp 1666464484
transform 1 0 7084 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A1
timestamp 1666464484
transform 1 0 6532 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__S
timestamp 1666464484
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A0
timestamp 1666464484
transform 1 0 5796 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A1
timestamp 1666464484
transform 1 0 5612 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__S
timestamp 1666464484
transform 1 0 5244 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A0
timestamp 1666464484
transform 1 0 7176 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A1
timestamp 1666464484
transform 1 0 7636 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__S
timestamp 1666464484
transform 1 0 5888 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A0
timestamp 1666464484
transform 1 0 11224 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A1
timestamp 1666464484
transform 1 0 11684 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__S
timestamp 1666464484
transform -1 0 12420 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A0
timestamp 1666464484
transform 1 0 11684 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A1
timestamp 1666464484
transform 1 0 10120 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__S
timestamp 1666464484
transform 1 0 11040 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A0
timestamp 1666464484
transform 1 0 18124 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A1
timestamp 1666464484
transform 1 0 16192 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__S
timestamp 1666464484
transform 1 0 17756 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A0
timestamp 1666464484
transform 1 0 19412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A1
timestamp 1666464484
transform 1 0 19596 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__S
timestamp 1666464484
transform 1 0 20792 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A0
timestamp 1666464484
transform 1 0 18400 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A1
timestamp 1666464484
transform 1 0 18584 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__S
timestamp 1666464484
transform 1 0 20148 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A0
timestamp 1666464484
transform 1 0 19780 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A1
timestamp 1666464484
transform 1 0 18032 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__S
timestamp 1666464484
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A1
timestamp 1666464484
transform -1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__S
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A1
timestamp 1666464484
transform 1 0 20700 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__S
timestamp 1666464484
transform 1 0 22080 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A1
timestamp 1666464484
transform -1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__S
timestamp 1666464484
transform 1 0 21988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1666464484
transform -1 0 23184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__B
timestamp 1666464484
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A0
timestamp 1666464484
transform 1 0 2944 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__S
timestamp 1666464484
transform -1 0 3680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A0
timestamp 1666464484
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__S
timestamp 1666464484
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A0
timestamp 1666464484
transform 1 0 3864 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__S
timestamp 1666464484
transform 1 0 3036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A0
timestamp 1666464484
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__S
timestamp 1666464484
transform 1 0 2760 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A0
timestamp 1666464484
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__S
timestamp 1666464484
transform 1 0 3220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A0
timestamp 1666464484
transform 1 0 2944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__S
timestamp 1666464484
transform 1 0 2392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A0
timestamp 1666464484
transform 1 0 2944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__S
timestamp 1666464484
transform -1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A0
timestamp 1666464484
transform 1 0 12880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__S
timestamp 1666464484
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A0
timestamp 1666464484
transform 1 0 19136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A1
timestamp 1666464484
transform -1 0 18768 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__S
timestamp 1666464484
transform -1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A0
timestamp 1666464484
transform 1 0 18308 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A1
timestamp 1666464484
transform -1 0 18676 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__S
timestamp 1666464484
transform 1 0 19688 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A0
timestamp 1666464484
transform 1 0 19412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A1
timestamp 1666464484
transform 1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A0
timestamp 1666464484
transform 1 0 19504 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A1
timestamp 1666464484
transform 1 0 18768 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A0
timestamp 1666464484
transform -1 0 17756 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A1
timestamp 1666464484
transform 1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A1
timestamp 1666464484
transform 1 0 20424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A1
timestamp 1666464484
transform -1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A1
timestamp 1666464484
transform 1 0 21620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A_N
timestamp 1666464484
transform 1 0 21988 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__B
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A0
timestamp 1666464484
transform 1 0 3772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__S
timestamp 1666464484
transform 1 0 3036 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A0
timestamp 1666464484
transform 1 0 3128 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__S
timestamp 1666464484
transform 1 0 2760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A0
timestamp 1666464484
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__S
timestamp 1666464484
transform -1 0 3128 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A0
timestamp 1666464484
transform 1 0 2944 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__S
timestamp 1666464484
transform 1 0 3036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A0
timestamp 1666464484
transform 1 0 3128 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__S
timestamp 1666464484
transform 1 0 2944 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A0
timestamp 1666464484
transform 1 0 2944 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__S
timestamp 1666464484
transform 1 0 4048 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A0
timestamp 1666464484
transform -1 0 13892 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A1
timestamp 1666464484
transform -1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__S
timestamp 1666464484
transform -1 0 13708 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A0
timestamp 1666464484
transform 1 0 11500 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__S
timestamp 1666464484
transform 1 0 10488 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A0
timestamp 1666464484
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A1
timestamp 1666464484
transform -1 0 15640 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__S
timestamp 1666464484
transform 1 0 15088 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A0
timestamp 1666464484
transform 1 0 18768 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A1
timestamp 1666464484
transform -1 0 18400 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__S
timestamp 1666464484
transform 1 0 17848 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A0
timestamp 1666464484
transform 1 0 18952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A1
timestamp 1666464484
transform -1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A0
timestamp 1666464484
transform 1 0 19504 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A1
timestamp 1666464484
transform -1 0 20792 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A0
timestamp 1666464484
transform 1 0 19412 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A1
timestamp 1666464484
transform -1 0 20240 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A1
timestamp 1666464484
transform 1 0 19688 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A1
timestamp 1666464484
transform -1 0 20424 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A1
timestamp 1666464484
transform 1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A_N
timestamp 1666464484
transform 1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__B
timestamp 1666464484
transform -1 0 23736 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A0
timestamp 1666464484
transform 1 0 3680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A1
timestamp 1666464484
transform 1 0 3128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__S
timestamp 1666464484
transform 1 0 2760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A0
timestamp 1666464484
transform 1 0 2944 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A1
timestamp 1666464484
transform 1 0 3128 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__S
timestamp 1666464484
transform 1 0 2760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A0
timestamp 1666464484
transform 1 0 11040 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A1
timestamp 1666464484
transform -1 0 13064 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__S
timestamp 1666464484
transform 1 0 12512 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A0
timestamp 1666464484
transform 1 0 3496 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A1
timestamp 1666464484
transform 1 0 3956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__S
timestamp 1666464484
transform -1 0 1748 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__D
timestamp 1666464484
transform -1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__D
timestamp 1666464484
transform -1 0 6072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__D
timestamp 1666464484
transform -1 0 13524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__D
timestamp 1666464484
transform -1 0 12788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__D
timestamp 1666464484
transform -1 0 12144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__D
timestamp 1666464484
transform -1 0 6808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_reg_wr_i_A
timestamp 1666464484
transform -1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_reg_wr_i_A
timestamp 1666464484
transform 1 0 10028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_reg_wr_i_A
timestamp 1666464484
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_reg_wr_i_A
timestamp 1666464484
transform -1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_reg_wr_i_A
timestamp 1666464484
transform 1 0 12420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_reg_wr_i_A
timestamp 1666464484
transform 1 0 10028 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_reg_wr_i_A
timestamp 1666464484
transform 1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_reg_wr_i_A
timestamp 1666464484
transform 1 0 12420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_reg_wr_i_A
timestamp 1666464484
transform 1 0 12420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout235_A
timestamp 1666464484
transform -1 0 6716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout236_A
timestamp 1666464484
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout237_A
timestamp 1666464484
transform -1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout238_A
timestamp 1666464484
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout239_A
timestamp 1666464484
transform 1 0 6532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout240_A
timestamp 1666464484
transform 1 0 5704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout241_A
timestamp 1666464484
transform 1 0 14352 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout242_A
timestamp 1666464484
transform -1 0 12052 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 54280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 1932 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 4324 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 6716 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 6348 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 8648 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 9292 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 9936 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 11224 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 12696 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 13800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 15088 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 16376 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 17480 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 18308 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 19872 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 20700 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 22264 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 23092 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 24748 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1666464484
transform -1 0 25484 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1666464484
transform -1 0 26680 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1666464484
transform -1 0 28244 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1666464484
transform -1 0 29256 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1666464484
transform -1 0 31464 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1666464484
transform -1 0 32292 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1666464484
transform -1 0 33856 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1666464484
transform -1 0 34408 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1666464484
transform -1 0 35512 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1666464484
transform -1 0 36616 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1666464484
transform -1 0 38640 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1666464484
transform -1 0 38180 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1666464484
transform -1 0 41032 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1666464484
transform -1 0 41400 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1666464484
transform -1 0 43424 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1666464484
transform -1 0 44620 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1666464484
transform -1 0 45356 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1666464484
transform -1 0 47012 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1666464484
transform -1 0 47748 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1666464484
transform -1 0 49404 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1666464484
transform -1 0 50508 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1666464484
transform -1 0 51796 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1666464484
transform -1 0 52164 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1666464484
transform -1 0 54188 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1666464484
transform -1 0 54556 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1666464484
transform -1 0 56580 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1666464484
transform -1 0 56488 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1666464484
transform -1 0 56212 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1666464484
transform -1 0 24564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1666464484
transform -1 0 25576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1666464484
transform -1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1666464484
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1666464484
transform -1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1666464484
transform -1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1666464484
transform -1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1666464484
transform -1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1666464484
transform -1 0 20148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1666464484
transform -1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1666464484
transform -1 0 20240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1666464484
transform -1 0 24012 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1666464484
transform -1 0 7544 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1666464484
transform -1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1666464484
transform -1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1666464484
transform -1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1666464484
transform -1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1666464484
transform -1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1666464484
transform -1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1666464484
transform -1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1666464484
transform -1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1666464484
transform -1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1666464484
transform -1 0 58420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1666464484
transform -1 0 55476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1666464484
transform -1 0 56028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1666464484
transform -1 0 57132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1666464484
transform -1 0 56580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1666464484
transform -1 0 56488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1666464484
transform -1 0 57776 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1666464484
transform -1 0 56948 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1666464484
transform -1 0 56396 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1666464484
transform -1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1666464484
transform -1 0 57592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1666464484
transform -1 0 57776 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1666464484
transform -1 0 57224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1666464484
transform -1 0 57776 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1666464484
transform -1 0 57040 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1666464484
transform -1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1666464484
transform -1 0 57224 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1666464484
transform -1 0 56488 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1666464484
transform -1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1666464484
transform -1 0 57040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1666464484
transform -1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1666464484
transform -1 0 58420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1666464484
transform -1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1666464484
transform -1 0 57224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1666464484
transform -1 0 58420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1666464484
transform -1 0 57132 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1666464484
transform -1 0 57592 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1666464484
transform -1 0 57776 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1666464484
transform -1 0 57592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1666464484
transform -1 0 57776 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1666464484
transform -1 0 57224 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1666464484
transform -1 0 57592 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1666464484
transform -1 0 57040 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1666464484
transform -1 0 57776 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1666464484
transform -1 0 57224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1666464484
transform -1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1666464484
transform -1 0 57776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1666464484
transform -1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1666464484
transform -1 0 57224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1666464484
transform -1 0 57776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1666464484
transform -1 0 57776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1666464484
transform -1 0 57592 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1666464484
transform -1 0 57776 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1666464484
transform -1 0 57592 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1666464484
transform -1 0 57776 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1666464484
transform -1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1666464484
transform -1 0 57592 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1666464484
transform -1 0 57776 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1666464484
transform -1 0 57776 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1666464484
transform -1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1666464484
transform -1 0 57592 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1666464484
transform -1 0 57776 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1666464484
transform -1 0 57776 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1666464484
transform -1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1666464484
transform -1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1666464484
transform -1 0 57776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1666464484
transform -1 0 57776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1666464484
transform -1 0 57592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1666464484
transform -1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1666464484
transform -1 0 57776 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1666464484
transform -1 0 57776 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1666464484
transform -1 0 57224 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1666464484
transform -1 0 56764 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1666464484
transform -1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1666464484
transform -1 0 57592 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1666464484
transform -1 0 57776 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input138_A
timestamp 1666464484
transform -1 0 57776 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input139_A
timestamp 1666464484
transform -1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input140_A
timestamp 1666464484
transform -1 0 57592 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input141_A
timestamp 1666464484
transform -1 0 57776 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input142_A
timestamp 1666464484
transform -1 0 55936 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input143_A
timestamp 1666464484
transform -1 0 57316 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input144_A
timestamp 1666464484
transform -1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input145_A
timestamp 1666464484
transform -1 0 36064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output147_A
timestamp 1666464484
transform -1 0 27416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output148_A
timestamp 1666464484
transform 1 0 28704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output149_A
timestamp 1666464484
transform 1 0 29808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1666464484
transform 1 0 30912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output151_A
timestamp 1666464484
transform -1 0 32476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output152_A
timestamp 1666464484
transform 1 0 33120 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output154_A
timestamp 1666464484
transform 1 0 1932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output155_A
timestamp 1666464484
transform 1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output156_A
timestamp 1666464484
transform -1 0 4140 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output157_A
timestamp 1666464484
transform -1 0 3864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output158_A
timestamp 1666464484
transform 1 0 1932 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output159_A
timestamp 1666464484
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output167_A
timestamp 1666464484
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1666464484
transform 1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1666464484
transform 1 0 2300 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1666464484
transform 1 0 2300 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output172_A
timestamp 1666464484
transform -1 0 2116 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output173_A
timestamp 1666464484
transform 1 0 2300 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1666464484
transform 1 0 2300 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1666464484
transform -1 0 2484 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output181_A
timestamp 1666464484
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output183_A
timestamp 1666464484
transform 1 0 3404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output184_A
timestamp 1666464484
transform 1 0 2852 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output185_A
timestamp 1666464484
transform -1 0 2484 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output186_A
timestamp 1666464484
transform 1 0 2300 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output187_A
timestamp 1666464484
transform -1 0 2484 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output188_A
timestamp 1666464484
transform -1 0 2484 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output189_A
timestamp 1666464484
transform 1 0 2300 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output190_A
timestamp 1666464484
transform 1 0 2300 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output191_A
timestamp 1666464484
transform -1 0 2484 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output192_A
timestamp 1666464484
transform 1 0 2300 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output193_A
timestamp 1666464484
transform 1 0 2300 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output194_A
timestamp 1666464484
transform -1 0 2484 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output195_A
timestamp 1666464484
transform -1 0 2484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output196_A
timestamp 1666464484
transform 1 0 2300 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output197_A
timestamp 1666464484
transform 1 0 2300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output198_A
timestamp 1666464484
transform -1 0 2484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output199_A
timestamp 1666464484
transform -1 0 2484 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output200_A
timestamp 1666464484
transform 1 0 2300 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output201_A
timestamp 1666464484
transform -1 0 2484 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output202_A
timestamp 1666464484
transform 1 0 2300 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output203_A
timestamp 1666464484
transform -1 0 2484 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output204_A
timestamp 1666464484
transform -1 0 2484 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output205_A
timestamp 1666464484
transform 1 0 2300 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output206_A
timestamp 1666464484
transform 1 0 2300 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output207_A
timestamp 1666464484
transform -1 0 2484 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output208_A
timestamp 1666464484
transform 1 0 2300 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output209_A
timestamp 1666464484
transform 1 0 2300 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output210_A
timestamp 1666464484
transform -1 0 2484 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1666464484
transform -1 0 2484 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output212_A
timestamp 1666464484
transform 1 0 2300 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output213_A
timestamp 1666464484
transform 1 0 2300 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output214_A
timestamp 1666464484
transform -1 0 2484 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output215_A
timestamp 1666464484
transform -1 0 2484 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output216_A
timestamp 1666464484
transform 1 0 2300 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output217_A
timestamp 1666464484
transform 1 0 37812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output218_A
timestamp 1666464484
transform 1 0 38548 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output220_A
timestamp 1666464484
transform 1 0 40388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output221_A
timestamp 1666464484
transform 1 0 41768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output222_A
timestamp 1666464484
transform 1 0 42964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output223_A
timestamp 1666464484
transform 1 0 43700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output226_A
timestamp 1666464484
transform 1 0 44712 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1666464484
transform 1 0 49496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output231_A
timestamp 1666464484
transform 1 0 50692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output232_A
timestamp 1666464484
transform 1 0 51428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10
timestamp 1666464484
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp 1666464484
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1666464484
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1666464484
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66
timestamp 1666464484
transform 1 0 7176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1666464484
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91
timestamp 1666464484
transform 1 0 9476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1666464484
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666464484
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1666464484
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126
timestamp 1666464484
transform 1 0 12696 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666464484
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1666464484
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_150
timestamp 1666464484
transform 1 0 14904 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1666464484
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1666464484
transform 1 0 17204 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1666464484
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1666464484
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1666464484
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_229
timestamp 1666464484
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_233
timestamp 1666464484
transform 1 0 22540 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_239
timestamp 1666464484
transform 1 0 23092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1666464484
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_261
timestamp 1666464484
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_270
timestamp 1666464484
transform 1 0 25944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1666464484
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_294
timestamp 1666464484
transform 1 0 28152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1666464484
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_313
timestamp 1666464484
transform 1 0 29900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_318
timestamp 1666464484
transform 1 0 30360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1666464484
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_343
timestamp 1666464484
transform 1 0 32660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_349
timestamp 1666464484
transform 1 0 33212 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_354
timestamp 1666464484
transform 1 0 33672 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1666464484
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_376
timestamp 1666464484
transform 1 0 35696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_386
timestamp 1666464484
transform 1 0 36616 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_399
timestamp 1666464484
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_407
timestamp 1666464484
transform 1 0 38548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1666464484
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_427
timestamp 1666464484
transform 1 0 40388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1666464484
transform 1 0 40940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_438
timestamp 1666464484
transform 1 0 41400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1666464484
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_455
timestamp 1666464484
transform 1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_463
timestamp 1666464484
transform 1 0 43700 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_469
timestamp 1666464484
transform 1 0 44252 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1666464484
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1666464484
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_481
timestamp 1666464484
transform 1 0 45356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_486
timestamp 1666464484
transform 1 0 45816 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1666464484
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_511
timestamp 1666464484
transform 1 0 48116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_517
timestamp 1666464484
transform 1 0 48668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_522
timestamp 1666464484
transform 1 0 49128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_528
timestamp 1666464484
transform 1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1666464484
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1666464484
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_547
timestamp 1666464484
transform 1 0 51428 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_553
timestamp 1666464484
transform 1 0 51980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1666464484
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_565
timestamp 1666464484
transform 1 0 53084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_570
timestamp 1666464484
transform 1 0 53544 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_582
timestamp 1666464484
transform 1 0 54648 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_595
timestamp 1666464484
transform 1 0 55844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_601
timestamp 1666464484
transform 1 0 56396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_605
timestamp 1666464484
transform 1 0 56764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1666464484
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1666464484
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1666464484
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11
timestamp 1666464484
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19
timestamp 1666464484
transform 1 0 2852 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1666464484
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1666464484
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1666464484
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_61
timestamp 1666464484
transform 1 0 6716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_67
timestamp 1666464484
transform 1 0 7268 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1666464484
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1666464484
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_101
timestamp 1666464484
transform 1 0 10396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_107
timestamp 1666464484
transform 1 0 10948 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1666464484
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_127
timestamp 1666464484
transform 1 0 12788 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1666464484
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_159
timestamp 1666464484
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_163
timestamp 1666464484
transform 1 0 16100 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666464484
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175
timestamp 1666464484
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1666464484
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1666464484
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_199
timestamp 1666464484
transform 1 0 19412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_216
timestamp 1666464484
transform 1 0 20976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666464484
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1666464484
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_240
timestamp 1666464484
transform 1 0 23184 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_246
timestamp 1666464484
transform 1 0 23736 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_255
timestamp 1666464484
transform 1 0 24564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_263
timestamp 1666464484
transform 1 0 25300 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_266 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1666464484
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1666464484
transform 1 0 27416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_294
timestamp 1666464484
transform 1 0 28152 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_302
timestamp 1666464484
transform 1 0 28888 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_310
timestamp 1666464484
transform 1 0 29624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_314
timestamp 1666464484
transform 1 0 29992 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_322
timestamp 1666464484
transform 1 0 30728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_326
timestamp 1666464484
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1666464484
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_341
timestamp 1666464484
transform 1 0 32476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_347
timestamp 1666464484
transform 1 0 33028 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_350
timestamp 1666464484
transform 1 0 33304 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_362
timestamp 1666464484
transform 1 0 34408 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_374
timestamp 1666464484
transform 1 0 35512 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_380
timestamp 1666464484
transform 1 0 36064 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_401
timestamp 1666464484
transform 1 0 37996 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_409
timestamp 1666464484
transform 1 0 38732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_421
timestamp 1666464484
transform 1 0 39836 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1666464484
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1666464484
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1666464484
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_449
timestamp 1666464484
transform 1 0 42412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_457
timestamp 1666464484
transform 1 0 43148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_465
timestamp 1666464484
transform 1 0 43884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_473
timestamp 1666464484
transform 1 0 44620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_476
timestamp 1666464484
transform 1 0 44896 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_488
timestamp 1666464484
transform 1 0 46000 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1666464484
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1666464484
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1666464484
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_529
timestamp 1666464484
transform 1 0 49772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_537
timestamp 1666464484
transform 1 0 50508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_541
timestamp 1666464484
transform 1 0 50876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_549
timestamp 1666464484
transform 1 0 51612 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1666464484
transform 1 0 52348 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_573
timestamp 1666464484
transform 1 0 53820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1666464484
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_584
timestamp 1666464484
transform 1 0 54832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_588
timestamp 1666464484
transform 1 0 55200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_591
timestamp 1666464484
transform 1 0 55476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_598
timestamp 1666464484
transform 1 0 56120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_605
timestamp 1666464484
transform 1 0 56764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_612
timestamp 1666464484
transform 1 0 57408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_617
timestamp 1666464484
transform 1 0 57868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_622
timestamp 1666464484
transform 1 0 58328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_18
timestamp 1666464484
transform 1 0 2760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1666464484
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1666464484
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_69
timestamp 1666464484
transform 1 0 7452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1666464484
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_89
timestamp 1666464484
transform 1 0 9292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_101
timestamp 1666464484
transform 1 0 10396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_107
timestamp 1666464484
transform 1 0 10948 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1666464484
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1666464484
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1666464484
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1666464484
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_172
timestamp 1666464484
transform 1 0 16928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1666464484
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1666464484
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1666464484
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1666464484
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_205
timestamp 1666464484
transform 1 0 19964 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_218
timestamp 1666464484
transform 1 0 21160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_226
timestamp 1666464484
transform 1 0 21896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1666464484
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1666464484
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1666464484
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1666464484
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1666464484
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1666464484
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1666464484
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1666464484
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_401
timestamp 1666464484
transform 1 0 37996 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_409
timestamp 1666464484
transform 1 0 38732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_414
timestamp 1666464484
transform 1 0 39192 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_425
timestamp 1666464484
transform 1 0 40204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_437
timestamp 1666464484
transform 1 0 41308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_449
timestamp 1666464484
transform 1 0 42412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_461
timestamp 1666464484
transform 1 0 43516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1666464484
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1666464484
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_489
timestamp 1666464484
transform 1 0 46092 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_494
timestamp 1666464484
transform 1 0 46552 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_500
timestamp 1666464484
transform 1 0 47104 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_512
timestamp 1666464484
transform 1 0 48208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_516
timestamp 1666464484
transform 1 0 48576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_522
timestamp 1666464484
transform 1 0 49128 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_530
timestamp 1666464484
transform 1 0 49864 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1666464484
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1666464484
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_557
timestamp 1666464484
transform 1 0 52348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_566
timestamp 1666464484
transform 1 0 53176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_572
timestamp 1666464484
transform 1 0 53728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_578
timestamp 1666464484
transform 1 0 54280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_582
timestamp 1666464484
transform 1 0 54648 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_589
timestamp 1666464484
transform 1 0 55292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_594
timestamp 1666464484
transform 1 0 55752 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_603
timestamp 1666464484
transform 1 0 56580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_610
timestamp 1666464484
transform 1 0 57224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_617
timestamp 1666464484
transform 1 0 57868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_623
timestamp 1666464484
transform 1 0 58420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1666464484
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_24
timestamp 1666464484
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_36
timestamp 1666464484
transform 1 0 4416 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1666464484
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1666464484
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_122
timestamp 1666464484
transform 1 0 12328 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_134
timestamp 1666464484
transform 1 0 13432 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1666464484
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_173
timestamp 1666464484
transform 1 0 17020 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_186
timestamp 1666464484
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1666464484
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_212
timestamp 1666464484
transform 1 0 20608 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1666464484
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_239
timestamp 1666464484
transform 1 0 23092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_251
timestamp 1666464484
transform 1 0 24196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_263
timestamp 1666464484
transform 1 0 25300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1666464484
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1666464484
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1666464484
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1666464484
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1666464484
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666464484
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1666464484
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1666464484
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1666464484
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1666464484
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1666464484
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1666464484
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1666464484
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1666464484
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1666464484
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1666464484
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1666464484
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1666464484
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1666464484
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1666464484
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1666464484
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1666464484
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1666464484
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1666464484
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1666464484
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1666464484
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_585
timestamp 1666464484
transform 1 0 54924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_590
timestamp 1666464484
transform 1 0 55384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_596
timestamp 1666464484
transform 1 0 55936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_602
timestamp 1666464484
transform 1 0 56488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_605
timestamp 1666464484
transform 1 0 56764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_614
timestamp 1666464484
transform 1 0 57592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1666464484
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_622
timestamp 1666464484
transform 1 0 58328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_9
timestamp 1666464484
transform 1 0 1932 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_17
timestamp 1666464484
transform 1 0 2668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1666464484
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp 1666464484
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1666464484
transform 1 0 6072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1666464484
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_158
timestamp 1666464484
transform 1 0 15640 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_170
timestamp 1666464484
transform 1 0 16744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666464484
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1666464484
transform 1 0 19596 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_207
timestamp 1666464484
transform 1 0 20148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1666464484
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_225
timestamp 1666464484
transform 1 0 21804 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_238
timestamp 1666464484
transform 1 0 23000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1666464484
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1666464484
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1666464484
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666464484
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666464484
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666464484
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666464484
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1666464484
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1666464484
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666464484
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1666464484
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1666464484
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1666464484
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1666464484
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1666464484
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666464484
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1666464484
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1666464484
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1666464484
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1666464484
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1666464484
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1666464484
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1666464484
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1666464484
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1666464484
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1666464484
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1666464484
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_589
timestamp 1666464484
transform 1 0 55292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_597
timestamp 1666464484
transform 1 0 56028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_603
timestamp 1666464484
transform 1 0 56580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_609
timestamp 1666464484
transform 1 0 57132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_616
timestamp 1666464484
transform 1 0 57776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1666464484
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1666464484
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1666464484
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1666464484
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1666464484
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1666464484
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_77
timestamp 1666464484
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_101
timestamp 1666464484
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1666464484
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_121
timestamp 1666464484
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp 1666464484
transform 1 0 19412 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_202
timestamp 1666464484
transform 1 0 19688 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214
timestamp 1666464484
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1666464484
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1666464484
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1666464484
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1666464484
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666464484
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666464484
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666464484
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666464484
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1666464484
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1666464484
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1666464484
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1666464484
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666464484
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1666464484
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1666464484
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1666464484
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1666464484
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666464484
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1666464484
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1666464484
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1666464484
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1666464484
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1666464484
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1666464484
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1666464484
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1666464484
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_597
timestamp 1666464484
transform 1 0 56028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_602
timestamp 1666464484
transform 1 0 56488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_608
timestamp 1666464484
transform 1 0 57040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_614
timestamp 1666464484
transform 1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_617
timestamp 1666464484
transform 1 0 57868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1666464484
transform 1 0 58420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_9
timestamp 1666464484
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1666464484
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1666464484
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_120
timestamp 1666464484
transform 1 0 12144 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1666464484
transform 1 0 13248 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1666464484
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_201
timestamp 1666464484
transform 1 0 19596 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_211
timestamp 1666464484
transform 1 0 20516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_223
timestamp 1666464484
transform 1 0 21620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_235
timestamp 1666464484
transform 1 0 22724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1666464484
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1666464484
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1666464484
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666464484
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666464484
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666464484
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666464484
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666464484
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666464484
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666464484
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666464484
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666464484
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666464484
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666464484
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666464484
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666464484
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666464484
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666464484
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1666464484
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1666464484
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1666464484
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1666464484
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1666464484
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1666464484
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1666464484
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_589
timestamp 1666464484
transform 1 0 55292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_595
timestamp 1666464484
transform 1 0 55844 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_598
timestamp 1666464484
transform 1 0 56120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_623
timestamp 1666464484
transform 1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_9
timestamp 1666464484
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1666464484
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_25
timestamp 1666464484
transform 1 0 3404 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_33
timestamp 1666464484
transform 1 0 4140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1666464484
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_99
timestamp 1666464484
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1666464484
transform 1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_152
timestamp 1666464484
transform 1 0 15088 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1666464484
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1666464484
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_192
timestamp 1666464484
transform 1 0 18768 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_198
timestamp 1666464484
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1666464484
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_229
timestamp 1666464484
transform 1 0 22172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_241
timestamp 1666464484
transform 1 0 23276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_253
timestamp 1666464484
transform 1 0 24380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_265
timestamp 1666464484
transform 1 0 25484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1666464484
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1666464484
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1666464484
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1666464484
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666464484
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666464484
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666464484
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666464484
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666464484
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666464484
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666464484
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666464484
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666464484
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666464484
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666464484
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666464484
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666464484
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666464484
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1666464484
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1666464484
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1666464484
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1666464484
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1666464484
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1666464484
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_585
timestamp 1666464484
transform 1 0 54924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_614
timestamp 1666464484
transform 1 0 57592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_617
timestamp 1666464484
transform 1 0 57868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 1666464484
transform 1 0 58420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1666464484
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1666464484
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1666464484
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_61
timestamp 1666464484
transform 1 0 6716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1666464484
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_203
timestamp 1666464484
transform 1 0 19780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_216
timestamp 1666464484
transform 1 0 20976 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_220
timestamp 1666464484
transform 1 0 21344 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1666464484
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_238
timestamp 1666464484
transform 1 0 23000 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1666464484
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1666464484
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1666464484
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666464484
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1666464484
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666464484
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666464484
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666464484
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666464484
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666464484
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666464484
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666464484
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666464484
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666464484
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666464484
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666464484
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666464484
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666464484
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1666464484
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1666464484
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1666464484
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1666464484
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1666464484
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1666464484
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1666464484
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1666464484
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_589
timestamp 1666464484
transform 1 0 55292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_594
timestamp 1666464484
transform 1 0 55752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_604
timestamp 1666464484
transform 1 0 56672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_610
timestamp 1666464484
transform 1 0 57224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_616
timestamp 1666464484
transform 1 0 57776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_623
timestamp 1666464484
transform 1 0 58420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1666464484
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1666464484
transform 1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_26
timestamp 1666464484
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1666464484
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1666464484
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_99
timestamp 1666464484
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 1666464484
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1666464484
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_202
timestamp 1666464484
transform 1 0 19688 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_214
timestamp 1666464484
transform 1 0 20792 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1666464484
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_240
timestamp 1666464484
transform 1 0 23184 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_246
timestamp 1666464484
transform 1 0 23736 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_258
timestamp 1666464484
transform 1 0 24840 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1666464484
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1666464484
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666464484
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1666464484
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1666464484
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666464484
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666464484
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666464484
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666464484
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1666464484
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666464484
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666464484
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666464484
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666464484
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666464484
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666464484
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666464484
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666464484
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666464484
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666464484
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666464484
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1666464484
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1666464484
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1666464484
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1666464484
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1666464484
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1666464484
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1666464484
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_597
timestamp 1666464484
transform 1 0 56028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_605
timestamp 1666464484
transform 1 0 56764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_608
timestamp 1666464484
transform 1 0 57040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1666464484
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_617
timestamp 1666464484
transform 1 0 57868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_623
timestamp 1666464484
transform 1 0 58420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1666464484
transform 1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_17
timestamp 1666464484
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1666464484
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_35
timestamp 1666464484
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_56
timestamp 1666464484
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_68
timestamp 1666464484
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1666464484
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_159
timestamp 1666464484
transform 1 0 15732 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_183
timestamp 1666464484
transform 1 0 17940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1666464484
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_225
timestamp 1666464484
transform 1 0 21804 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_238
timestamp 1666464484
transform 1 0 23000 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1666464484
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1666464484
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666464484
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1666464484
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666464484
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1666464484
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1666464484
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666464484
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666464484
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666464484
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1666464484
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1666464484
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666464484
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666464484
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666464484
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666464484
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666464484
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666464484
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666464484
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666464484
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666464484
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1666464484
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1666464484
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1666464484
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1666464484
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1666464484
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1666464484
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1666464484
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1666464484
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1666464484
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_601
timestamp 1666464484
transform 1 0 56396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_607
timestamp 1666464484
transform 1 0 56948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_610
timestamp 1666464484
transform 1 0 57224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_616
timestamp 1666464484
transform 1 0 57776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_623
timestamp 1666464484
transform 1 0 58420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp 1666464484
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_25
timestamp 1666464484
transform 1 0 3404 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1666464484
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1666464484
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_121
timestamp 1666464484
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_230
timestamp 1666464484
transform 1 0 22264 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_242
timestamp 1666464484
transform 1 0 23368 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_254
timestamp 1666464484
transform 1 0 24472 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_266
timestamp 1666464484
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1666464484
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1666464484
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1666464484
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1666464484
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1666464484
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1666464484
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666464484
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666464484
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1666464484
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666464484
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1666464484
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1666464484
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1666464484
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1666464484
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1666464484
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666464484
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666464484
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666464484
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666464484
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666464484
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1666464484
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1666464484
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1666464484
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1666464484
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1666464484
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1666464484
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1666464484
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_585
timestamp 1666464484
transform 1 0 54924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_593
timestamp 1666464484
transform 1 0 55660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1666464484
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_617
timestamp 1666464484
transform 1 0 57868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_623
timestamp 1666464484
transform 1 0 58420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_9
timestamp 1666464484
transform 1 0 1932 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_17
timestamp 1666464484
transform 1 0 2668 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1666464484
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1666464484
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_52
timestamp 1666464484
transform 1 0 5888 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_58
timestamp 1666464484
transform 1 0 6440 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_70
timestamp 1666464484
transform 1 0 7544 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1666464484
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_101
timestamp 1666464484
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1666464484
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_145
timestamp 1666464484
transform 1 0 14444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_157
timestamp 1666464484
transform 1 0 15548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_169
timestamp 1666464484
transform 1 0 16652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_181
timestamp 1666464484
transform 1 0 17756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1666464484
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_205
timestamp 1666464484
transform 1 0 19964 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_210
timestamp 1666464484
transform 1 0 20424 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1666464484
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1666464484
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_237
timestamp 1666464484
transform 1 0 22908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1666464484
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1666464484
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666464484
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666464484
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1666464484
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1666464484
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1666464484
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1666464484
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666464484
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1666464484
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1666464484
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1666464484
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1666464484
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666464484
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666464484
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666464484
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666464484
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666464484
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666464484
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666464484
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666464484
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666464484
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1666464484
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1666464484
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1666464484
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1666464484
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1666464484
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1666464484
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1666464484
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1666464484
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_589
timestamp 1666464484
transform 1 0 55292 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_595
timestamp 1666464484
transform 1 0 55844 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_598
timestamp 1666464484
transform 1 0 56120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_623
timestamp 1666464484
transform 1 0 58420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1666464484
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_33
timestamp 1666464484
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1666464484
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_97
timestamp 1666464484
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1666464484
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_145
timestamp 1666464484
transform 1 0 14444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_157
timestamp 1666464484
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1666464484
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1666464484
transform 1 0 19596 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_209
timestamp 1666464484
transform 1 0 20332 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1666464484
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1666464484
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1666464484
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666464484
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666464484
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666464484
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666464484
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1666464484
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666464484
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1666464484
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1666464484
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1666464484
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1666464484
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1666464484
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666464484
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666464484
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666464484
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666464484
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666464484
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1666464484
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1666464484
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1666464484
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1666464484
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1666464484
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1666464484
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1666464484
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1666464484
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_597
timestamp 1666464484
transform 1 0 56028 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_605
timestamp 1666464484
transform 1 0 56764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_608
timestamp 1666464484
transform 1 0 57040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_614
timestamp 1666464484
transform 1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_617
timestamp 1666464484
transform 1 0 57868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_623
timestamp 1666464484
transform 1 0 58420 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1666464484
transform 1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_13
timestamp 1666464484
transform 1 0 2300 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_16
timestamp 1666464484
transform 1 0 2576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1666464484
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_49
timestamp 1666464484
transform 1 0 5612 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_71
timestamp 1666464484
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_124
timestamp 1666464484
transform 1 0 12512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_130
timestamp 1666464484
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1666464484
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1666464484
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_171
timestamp 1666464484
transform 1 0 16836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_183
timestamp 1666464484
transform 1 0 17940 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1666464484
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1666464484
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_204
timestamp 1666464484
transform 1 0 19872 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_216
timestamp 1666464484
transform 1 0 20976 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_228
timestamp 1666464484
transform 1 0 22080 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_240
timestamp 1666464484
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666464484
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666464484
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1666464484
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1666464484
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1666464484
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666464484
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666464484
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1666464484
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1666464484
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1666464484
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1666464484
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1666464484
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1666464484
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1666464484
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1666464484
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666464484
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666464484
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666464484
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666464484
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1666464484
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1666464484
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1666464484
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1666464484
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1666464484
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1666464484
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1666464484
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1666464484
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1666464484
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_601
timestamp 1666464484
transform 1 0 56396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_607
timestamp 1666464484
transform 1 0 56948 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_610
timestamp 1666464484
transform 1 0 57224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_616
timestamp 1666464484
transform 1 0 57776 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_623
timestamp 1666464484
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_18
timestamp 1666464484
transform 1 0 2760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_25
timestamp 1666464484
transform 1 0 3404 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_33
timestamp 1666464484
transform 1 0 4140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1666464484
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_121
timestamp 1666464484
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_126
timestamp 1666464484
transform 1 0 12696 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_153
timestamp 1666464484
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1666464484
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_189
timestamp 1666464484
transform 1 0 18492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_202
timestamp 1666464484
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_206
timestamp 1666464484
transform 1 0 20056 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_210
timestamp 1666464484
transform 1 0 20424 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1666464484
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1666464484
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1666464484
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666464484
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666464484
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1666464484
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666464484
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666464484
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666464484
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1666464484
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1666464484
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1666464484
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1666464484
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1666464484
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666464484
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666464484
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666464484
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666464484
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666464484
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1666464484
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1666464484
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1666464484
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1666464484
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1666464484
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1666464484
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1666464484
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_597
timestamp 1666464484
transform 1 0 56028 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_605
timestamp 1666464484
transform 1 0 56764 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_608
timestamp 1666464484
transform 1 0 57040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_614
timestamp 1666464484
transform 1 0 57592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_617
timestamp 1666464484
transform 1 0 57868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_623
timestamp 1666464484
transform 1 0 58420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_18
timestamp 1666464484
transform 1 0 2760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1666464484
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1666464484
transform 1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_62
timestamp 1666464484
transform 1 0 6808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_74
timestamp 1666464484
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1666464484
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1666464484
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_208
timestamp 1666464484
transform 1 0 20240 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_214
timestamp 1666464484
transform 1 0 20792 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1666464484
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_230
timestamp 1666464484
transform 1 0 22264 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_242
timestamp 1666464484
transform 1 0 23368 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1666464484
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666464484
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666464484
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666464484
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1666464484
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1666464484
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1666464484
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666464484
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1666464484
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1666464484
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1666464484
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1666464484
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666464484
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666464484
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1666464484
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1666464484
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1666464484
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666464484
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666464484
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666464484
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666464484
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1666464484
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1666464484
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1666464484
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1666464484
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1666464484
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1666464484
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1666464484
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1666464484
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1666464484
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_601
timestamp 1666464484
transform 1 0 56396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_623
timestamp 1666464484
transform 1 0 58420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1666464484
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_19
timestamp 1666464484
transform 1 0 2852 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_22
timestamp 1666464484
transform 1 0 3128 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_28
timestamp 1666464484
transform 1 0 3680 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_40
timestamp 1666464484
transform 1 0 4784 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1666464484
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1666464484
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1666464484
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_142
timestamp 1666464484
transform 1 0 14168 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1666464484
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1666464484
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1666464484
transform 1 0 19320 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_204
timestamp 1666464484
transform 1 0 19872 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_212
timestamp 1666464484
transform 1 0 20608 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1666464484
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1666464484
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1666464484
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1666464484
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666464484
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1666464484
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1666464484
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1666464484
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1666464484
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666464484
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1666464484
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1666464484
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1666464484
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1666464484
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1666464484
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666464484
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666464484
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666464484
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666464484
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666464484
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1666464484
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1666464484
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1666464484
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1666464484
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1666464484
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1666464484
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1666464484
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1666464484
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_609
timestamp 1666464484
transform 1 0 57132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_614
timestamp 1666464484
transform 1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_617
timestamp 1666464484
transform 1 0 57868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_623
timestamp 1666464484
transform 1 0 58420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_11
timestamp 1666464484
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1666464484
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1666464484
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_108
timestamp 1666464484
transform 1 0 11040 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_120
timestamp 1666464484
transform 1 0 12144 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1666464484
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_180
timestamp 1666464484
transform 1 0 17664 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1666464484
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_201
timestamp 1666464484
transform 1 0 19596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_213
timestamp 1666464484
transform 1 0 20700 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_225
timestamp 1666464484
transform 1 0 21804 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_237
timestamp 1666464484
transform 1 0 22908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1666464484
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1666464484
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666464484
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666464484
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666464484
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666464484
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666464484
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666464484
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666464484
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666464484
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1666464484
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1666464484
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666464484
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1666464484
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1666464484
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1666464484
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1666464484
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666464484
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666464484
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666464484
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666464484
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1666464484
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1666464484
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1666464484
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1666464484
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1666464484
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1666464484
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1666464484
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1666464484
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_589
timestamp 1666464484
transform 1 0 55292 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_594
timestamp 1666464484
transform 1 0 55752 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_606
timestamp 1666464484
transform 1 0 56856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_610
timestamp 1666464484
transform 1 0 57224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_616
timestamp 1666464484
transform 1 0 57776 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_623
timestamp 1666464484
transform 1 0 58420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_9
timestamp 1666464484
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_187
timestamp 1666464484
transform 1 0 18308 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1666464484
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1666464484
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_210
timestamp 1666464484
transform 1 0 20424 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1666464484
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1666464484
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1666464484
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666464484
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666464484
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1666464484
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1666464484
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1666464484
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1666464484
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666464484
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1666464484
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1666464484
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1666464484
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1666464484
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666464484
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1666464484
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1666464484
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1666464484
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1666464484
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666464484
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1666464484
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1666464484
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1666464484
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1666464484
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1666464484
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1666464484
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1666464484
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1666464484
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1666464484
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_609
timestamp 1666464484
transform 1 0 57132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_614
timestamp 1666464484
transform 1 0 57592 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_617
timestamp 1666464484
transform 1 0 57868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_623
timestamp 1666464484
transform 1 0 58420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_9
timestamp 1666464484
transform 1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_16
timestamp 1666464484
transform 1 0 2576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1666464484
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1666464484
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666464484
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666464484
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1666464484
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666464484
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1666464484
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1666464484
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1666464484
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1666464484
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666464484
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666464484
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666464484
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1666464484
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1666464484
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666464484
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1666464484
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1666464484
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1666464484
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1666464484
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666464484
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666464484
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666464484
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666464484
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1666464484
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1666464484
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1666464484
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1666464484
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1666464484
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1666464484
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1666464484
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1666464484
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1666464484
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_601
timestamp 1666464484
transform 1 0 56396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_623
timestamp 1666464484
transform 1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1666464484
transform 1 0 2760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1666464484
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1666464484
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1666464484
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_117
timestamp 1666464484
transform 1 0 11868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_129
timestamp 1666464484
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_152
timestamp 1666464484
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1666464484
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_209
timestamp 1666464484
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1666464484
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_229
timestamp 1666464484
transform 1 0 22172 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_241
timestamp 1666464484
transform 1 0 23276 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_253
timestamp 1666464484
transform 1 0 24380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_265
timestamp 1666464484
transform 1 0 25484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1666464484
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666464484
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1666464484
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1666464484
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666464484
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1666464484
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1666464484
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1666464484
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1666464484
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666464484
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1666464484
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1666464484
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1666464484
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1666464484
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666464484
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1666464484
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1666464484
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1666464484
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1666464484
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1666464484
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1666464484
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1666464484
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1666464484
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1666464484
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1666464484
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1666464484
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1666464484
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1666464484
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1666464484
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1666464484
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_617
timestamp 1666464484
transform 1 0 57868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_623
timestamp 1666464484
transform 1 0 58420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 1666464484
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_17
timestamp 1666464484
transform 1 0 2668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1666464484
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_33
timestamp 1666464484
transform 1 0 4140 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_63
timestamp 1666464484
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1666464484
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_146
timestamp 1666464484
transform 1 0 14536 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_158
timestamp 1666464484
transform 1 0 15640 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_170
timestamp 1666464484
transform 1 0 16744 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_182
timestamp 1666464484
transform 1 0 17848 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1666464484
transform 1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1666464484
transform 1 0 20240 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_217
timestamp 1666464484
transform 1 0 21068 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_229
timestamp 1666464484
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_241
timestamp 1666464484
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1666464484
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666464484
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666464484
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1666464484
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666464484
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666464484
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1666464484
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1666464484
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1666464484
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1666464484
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666464484
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1666464484
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1666464484
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1666464484
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666464484
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666464484
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1666464484
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1666464484
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1666464484
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1666464484
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666464484
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1666464484
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666464484
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666464484
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1666464484
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1666464484
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1666464484
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1666464484
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1666464484
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1666464484
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1666464484
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1666464484
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1666464484
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1666464484
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_613
timestamp 1666464484
transform 1 0 57500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_616
timestamp 1666464484
transform 1 0 57776 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_623
timestamp 1666464484
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1666464484
transform 1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_24
timestamp 1666464484
transform 1 0 3312 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_30
timestamp 1666464484
transform 1 0 3864 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_42
timestamp 1666464484
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1666464484
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_99
timestamp 1666464484
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1666464484
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_152
timestamp 1666464484
transform 1 0 15088 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1666464484
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_194
timestamp 1666464484
transform 1 0 18952 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_200
timestamp 1666464484
transform 1 0 19504 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1666464484
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1666464484
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666464484
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666464484
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666464484
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666464484
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1666464484
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1666464484
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1666464484
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666464484
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1666464484
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1666464484
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1666464484
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1666464484
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1666464484
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1666464484
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1666464484
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1666464484
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1666464484
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1666464484
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1666464484
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1666464484
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1666464484
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1666464484
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1666464484
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1666464484
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1666464484
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1666464484
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1666464484
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1666464484
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1666464484
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1666464484
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1666464484
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_609
timestamp 1666464484
transform 1 0 57132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_614
timestamp 1666464484
transform 1 0 57592 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_617
timestamp 1666464484
transform 1 0 57868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_623
timestamp 1666464484
transform 1 0 58420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_11
timestamp 1666464484
transform 1 0 2116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_17
timestamp 1666464484
transform 1 0 2668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1666464484
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_49
timestamp 1666464484
transform 1 0 5612 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_72
timestamp 1666464484
transform 1 0 7728 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_107
timestamp 1666464484
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_119
timestamp 1666464484
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp 1666464484
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1666464484
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_202
timestamp 1666464484
transform 1 0 19688 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_208
timestamp 1666464484
transform 1 0 20240 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_220
timestamp 1666464484
transform 1 0 21344 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_232
timestamp 1666464484
transform 1 0 22448 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1666464484
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666464484
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1666464484
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666464484
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1666464484
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1666464484
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1666464484
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666464484
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666464484
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1666464484
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1666464484
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1666464484
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1666464484
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1666464484
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1666464484
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1666464484
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1666464484
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1666464484
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666464484
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1666464484
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1666464484
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1666464484
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1666464484
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1666464484
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1666464484
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1666464484
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1666464484
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1666464484
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1666464484
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1666464484
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1666464484
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1666464484
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_603
timestamp 1666464484
transform 1 0 56580 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_613
timestamp 1666464484
transform 1 0 57500 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_623
timestamp 1666464484
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1666464484
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_102
timestamp 1666464484
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_121
timestamp 1666464484
transform 1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_188
timestamp 1666464484
transform 1 0 18400 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1666464484
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_207
timestamp 1666464484
transform 1 0 20148 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1666464484
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1666464484
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1666464484
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666464484
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1666464484
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666464484
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1666464484
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1666464484
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1666464484
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1666464484
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1666464484
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1666464484
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1666464484
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1666464484
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1666464484
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1666464484
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1666464484
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1666464484
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666464484
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1666464484
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1666464484
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1666464484
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1666464484
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1666464484
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1666464484
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1666464484
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1666464484
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1666464484
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_617
timestamp 1666464484
transform 1 0 57868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_623
timestamp 1666464484
transform 1 0 58420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_9
timestamp 1666464484
transform 1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_13
timestamp 1666464484
transform 1 0 2300 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_17
timestamp 1666464484
transform 1 0 2668 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1666464484
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_184
timestamp 1666464484
transform 1 0 18032 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666464484
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666464484
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1666464484
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1666464484
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666464484
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1666464484
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1666464484
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1666464484
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1666464484
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666464484
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1666464484
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1666464484
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1666464484
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1666464484
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1666464484
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1666464484
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1666464484
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1666464484
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1666464484
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666464484
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1666464484
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1666464484
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1666464484
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1666464484
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1666464484
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1666464484
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1666464484
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1666464484
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1666464484
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1666464484
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1666464484
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1666464484
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1666464484
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_613
timestamp 1666464484
transform 1 0 57500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_616
timestamp 1666464484
transform 1 0 57776 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_623
timestamp 1666464484
transform 1 0 58420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_18
timestamp 1666464484
transform 1 0 2760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_25
timestamp 1666464484
transform 1 0 3404 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_31
timestamp 1666464484
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_43
timestamp 1666464484
transform 1 0 5060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1666464484
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_61
timestamp 1666464484
transform 1 0 6716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_73
timestamp 1666464484
transform 1 0 7820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1666464484
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1666464484
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1666464484
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_138
timestamp 1666464484
transform 1 0 13800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1666464484
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_177
timestamp 1666464484
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_182
timestamp 1666464484
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_189
timestamp 1666464484
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_196
timestamp 1666464484
transform 1 0 19136 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_208
timestamp 1666464484
transform 1 0 20240 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1666464484
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666464484
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1666464484
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666464484
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666464484
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666464484
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1666464484
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1666464484
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666464484
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666464484
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1666464484
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1666464484
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1666464484
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1666464484
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666464484
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1666464484
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1666464484
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1666464484
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1666464484
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666464484
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1666464484
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1666464484
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1666464484
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1666464484
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666464484
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1666464484
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1666464484
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1666464484
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1666464484
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1666464484
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1666464484
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1666464484
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1666464484
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1666464484
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1666464484
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_9
timestamp 1666464484
transform 1 0 1932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_17
timestamp 1666464484
transform 1 0 2668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1666464484
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1666464484
transform 1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_117
timestamp 1666464484
transform 1 0 11868 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_129
timestamp 1666464484
transform 1 0 12972 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1666464484
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_176
timestamp 1666464484
transform 1 0 17296 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_184
timestamp 1666464484
transform 1 0 18032 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_201
timestamp 1666464484
transform 1 0 19596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_213
timestamp 1666464484
transform 1 0 20700 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_225
timestamp 1666464484
transform 1 0 21804 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_237
timestamp 1666464484
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1666464484
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666464484
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666464484
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1666464484
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1666464484
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666464484
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1666464484
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1666464484
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1666464484
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1666464484
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666464484
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1666464484
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1666464484
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1666464484
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1666464484
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666464484
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1666464484
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1666464484
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1666464484
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1666464484
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1666464484
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1666464484
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666464484
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666464484
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1666464484
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1666464484
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1666464484
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1666464484
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1666464484
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1666464484
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1666464484
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1666464484
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1666464484
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1666464484
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_613
timestamp 1666464484
transform 1 0 57500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_616
timestamp 1666464484
transform 1 0 57776 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_623
timestamp 1666464484
transform 1 0 58420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_42
timestamp 1666464484
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1666464484
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_80
timestamp 1666464484
transform 1 0 8464 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_92
timestamp 1666464484
transform 1 0 9568 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_104
timestamp 1666464484
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_175
timestamp 1666464484
transform 1 0 17204 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_179
timestamp 1666464484
transform 1 0 17572 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1666464484
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_202
timestamp 1666464484
transform 1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_208
timestamp 1666464484
transform 1 0 20240 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1666464484
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1666464484
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666464484
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1666464484
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666464484
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1666464484
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1666464484
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1666464484
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1666464484
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666464484
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1666464484
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666464484
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1666464484
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1666464484
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1666464484
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1666464484
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1666464484
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1666464484
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1666464484
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1666464484
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1666464484
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1666464484
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1666464484
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1666464484
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666464484
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1666464484
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1666464484
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1666464484
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1666464484
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1666464484
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1666464484
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1666464484
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1666464484
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_609
timestamp 1666464484
transform 1 0 57132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_614
timestamp 1666464484
transform 1 0 57592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_617
timestamp 1666464484
transform 1 0 57868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_623
timestamp 1666464484
transform 1 0 58420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_9
timestamp 1666464484
transform 1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_16
timestamp 1666464484
transform 1 0 2576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1666464484
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1666464484
transform 1 0 16836 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_175
timestamp 1666464484
transform 1 0 17204 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1666464484
transform 1 0 18032 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1666464484
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_214
timestamp 1666464484
transform 1 0 20792 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_226
timestamp 1666464484
transform 1 0 21896 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_238
timestamp 1666464484
transform 1 0 23000 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666464484
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666464484
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1666464484
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1666464484
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1666464484
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1666464484
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1666464484
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1666464484
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1666464484
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1666464484
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1666464484
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1666464484
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1666464484
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1666464484
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1666464484
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1666464484
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1666464484
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1666464484
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1666464484
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1666464484
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666464484
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666464484
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666464484
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1666464484
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1666464484
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1666464484
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1666464484
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1666464484
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1666464484
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1666464484
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1666464484
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1666464484
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1666464484
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_613
timestamp 1666464484
transform 1 0 57500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_623
timestamp 1666464484
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_9
timestamp 1666464484
transform 1 0 1932 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_17
timestamp 1666464484
transform 1 0 2668 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_22
timestamp 1666464484
transform 1 0 3128 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_34
timestamp 1666464484
transform 1 0 4232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_46
timestamp 1666464484
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1666464484
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1666464484
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_146
timestamp 1666464484
transform 1 0 14536 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp 1666464484
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1666464484
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1666464484
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1666464484
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_199
timestamp 1666464484
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_211
timestamp 1666464484
transform 1 0 20516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666464484
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666464484
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666464484
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666464484
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1666464484
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1666464484
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1666464484
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1666464484
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666464484
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1666464484
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1666464484
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1666464484
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1666464484
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1666464484
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1666464484
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1666464484
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1666464484
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1666464484
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1666464484
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1666464484
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1666464484
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1666464484
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1666464484
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666464484
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1666464484
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1666464484
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1666464484
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1666464484
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1666464484
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1666464484
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1666464484
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1666464484
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1666464484
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_617
timestamp 1666464484
transform 1 0 57868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_623
timestamp 1666464484
transform 1 0 58420 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_18
timestamp 1666464484
transform 1 0 2760 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1666464484
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_47
timestamp 1666464484
transform 1 0 5428 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_71
timestamp 1666464484
transform 1 0 7636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_105
timestamp 1666464484
transform 1 0 10764 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_126
timestamp 1666464484
transform 1 0 12696 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1666464484
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_203
timestamp 1666464484
transform 1 0 19780 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_215
timestamp 1666464484
transform 1 0 20884 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_227
timestamp 1666464484
transform 1 0 21988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_239
timestamp 1666464484
transform 1 0 23092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666464484
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1666464484
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666464484
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1666464484
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1666464484
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1666464484
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1666464484
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666464484
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1666464484
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1666464484
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1666464484
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1666464484
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666464484
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1666464484
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1666464484
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1666464484
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1666464484
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1666464484
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1666464484
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1666464484
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1666464484
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1666464484
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1666464484
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1666464484
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1666464484
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1666464484
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1666464484
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1666464484
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1666464484
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1666464484
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1666464484
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_613
timestamp 1666464484
transform 1 0 57500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_616
timestamp 1666464484
transform 1 0 57776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_623
timestamp 1666464484
transform 1 0 58420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_9
timestamp 1666464484
transform 1 0 1932 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_17
timestamp 1666464484
transform 1 0 2668 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_32
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_40
timestamp 1666464484
transform 1 0 4784 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_46
timestamp 1666464484
transform 1 0 5336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1666464484
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_99
timestamp 1666464484
transform 1 0 10212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_123
timestamp 1666464484
transform 1 0 12420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1666464484
transform 1 0 13524 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1666464484
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_177
timestamp 1666464484
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_188
timestamp 1666464484
transform 1 0 18400 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_201
timestamp 1666464484
transform 1 0 19596 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1666464484
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1666464484
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666464484
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666464484
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666464484
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666464484
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666464484
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1666464484
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1666464484
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666464484
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1666464484
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1666464484
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1666464484
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1666464484
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1666464484
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1666464484
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1666464484
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1666464484
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1666464484
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666464484
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1666464484
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1666464484
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1666464484
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1666464484
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666464484
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1666464484
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1666464484
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1666464484
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1666464484
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1666464484
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1666464484
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1666464484
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1666464484
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1666464484
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1666464484
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1666464484
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1666464484
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_9
timestamp 1666464484
transform 1 0 1932 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_16
timestamp 1666464484
transform 1 0 2576 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1666464484
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_51
timestamp 1666464484
transform 1 0 5796 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_59
timestamp 1666464484
transform 1 0 6532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1666464484
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1666464484
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1666464484
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_164
timestamp 1666464484
transform 1 0 16192 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_176
timestamp 1666464484
transform 1 0 17296 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_188
timestamp 1666464484
transform 1 0 18400 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1666464484
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666464484
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666464484
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666464484
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666464484
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1666464484
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1666464484
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666464484
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1666464484
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1666464484
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1666464484
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1666464484
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666464484
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1666464484
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1666464484
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1666464484
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1666464484
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1666464484
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1666464484
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1666464484
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1666464484
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1666464484
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1666464484
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666464484
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1666464484
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1666464484
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1666464484
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1666464484
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1666464484
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1666464484
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1666464484
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1666464484
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1666464484
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1666464484
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1666464484
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1666464484
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_613
timestamp 1666464484
transform 1 0 57500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_616
timestamp 1666464484
transform 1 0 57776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_623
timestamp 1666464484
transform 1 0 58420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_18
timestamp 1666464484
transform 1 0 2760 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_24
timestamp 1666464484
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_36
timestamp 1666464484
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1666464484
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_121
timestamp 1666464484
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_187
timestamp 1666464484
transform 1 0 18308 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_190
timestamp 1666464484
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_203
timestamp 1666464484
transform 1 0 19780 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_209
timestamp 1666464484
transform 1 0 20332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1666464484
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1666464484
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1666464484
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666464484
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1666464484
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1666464484
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1666464484
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1666464484
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1666464484
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666464484
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1666464484
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1666464484
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1666464484
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1666464484
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666464484
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1666464484
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1666464484
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1666464484
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1666464484
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1666464484
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1666464484
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1666464484
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1666464484
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1666464484
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666464484
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1666464484
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1666464484
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1666464484
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1666464484
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1666464484
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1666464484
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1666464484
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1666464484
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1666464484
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_609
timestamp 1666464484
transform 1 0 57132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_614
timestamp 1666464484
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_617
timestamp 1666464484
transform 1 0 57868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1666464484
transform 1 0 58420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_9
timestamp 1666464484
transform 1 0 1932 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_17
timestamp 1666464484
transform 1 0 2668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_20
timestamp 1666464484
transform 1 0 2944 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1666464484
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_185
timestamp 1666464484
transform 1 0 18124 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_188
timestamp 1666464484
transform 1 0 18400 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_210
timestamp 1666464484
transform 1 0 20424 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_216
timestamp 1666464484
transform 1 0 20976 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_228
timestamp 1666464484
transform 1 0 22080 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_240
timestamp 1666464484
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666464484
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666464484
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1666464484
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1666464484
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666464484
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1666464484
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1666464484
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1666464484
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1666464484
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666464484
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1666464484
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1666464484
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1666464484
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1666464484
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666464484
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1666464484
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1666464484
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1666464484
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1666464484
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1666464484
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1666464484
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1666464484
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1666464484
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1666464484
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1666464484
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1666464484
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1666464484
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1666464484
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1666464484
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1666464484
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1666464484
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1666464484
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_601
timestamp 1666464484
transform 1 0 56396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_609
timestamp 1666464484
transform 1 0 57132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_622
timestamp 1666464484
transform 1 0 58328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_18
timestamp 1666464484
transform 1 0 2760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_24
timestamp 1666464484
transform 1 0 3312 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_30
timestamp 1666464484
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_42
timestamp 1666464484
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1666464484
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_77
timestamp 1666464484
transform 1 0 8188 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_98
timestamp 1666464484
transform 1 0 10120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1666464484
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_191
timestamp 1666464484
transform 1 0 18676 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_207
timestamp 1666464484
transform 1 0 20148 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1666464484
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666464484
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666464484
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666464484
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666464484
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1666464484
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1666464484
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1666464484
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1666464484
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666464484
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1666464484
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1666464484
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1666464484
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1666464484
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666464484
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1666464484
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1666464484
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1666464484
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1666464484
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666464484
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1666464484
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1666464484
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1666464484
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1666464484
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1666464484
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1666464484
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1666464484
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1666464484
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1666464484
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1666464484
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1666464484
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1666464484
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1666464484
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1666464484
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_609
timestamp 1666464484
transform 1 0 57132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_614
timestamp 1666464484
transform 1 0 57592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_617
timestamp 1666464484
transform 1 0 57868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1666464484
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_9
timestamp 1666464484
transform 1 0 1932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_16
timestamp 1666464484
transform 1 0 2576 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_22
timestamp 1666464484
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_34
timestamp 1666464484
transform 1 0 4232 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_46
timestamp 1666464484
transform 1 0 5336 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_58
timestamp 1666464484
transform 1 0 6440 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_70
timestamp 1666464484
transform 1 0 7544 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1666464484
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_182
timestamp 1666464484
transform 1 0 17848 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_190
timestamp 1666464484
transform 1 0 18584 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1666464484
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_208
timestamp 1666464484
transform 1 0 20240 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_214
timestamp 1666464484
transform 1 0 20792 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_226
timestamp 1666464484
transform 1 0 21896 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_238
timestamp 1666464484
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1666464484
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666464484
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1666464484
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1666464484
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1666464484
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666464484
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1666464484
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1666464484
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1666464484
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1666464484
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1666464484
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1666464484
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1666464484
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1666464484
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1666464484
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1666464484
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1666464484
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1666464484
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1666464484
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1666464484
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1666464484
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666464484
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666464484
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1666464484
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1666464484
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1666464484
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1666464484
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1666464484
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1666464484
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1666464484
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1666464484
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1666464484
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1666464484
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1666464484
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_613
timestamp 1666464484
transform 1 0 57500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_616
timestamp 1666464484
transform 1 0 57776 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_623
timestamp 1666464484
transform 1 0 58420 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_18
timestamp 1666464484
transform 1 0 2760 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_28
timestamp 1666464484
transform 1 0 3680 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_34
timestamp 1666464484
transform 1 0 4232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_46
timestamp 1666464484
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1666464484
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_187
timestamp 1666464484
transform 1 0 18308 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_191
timestamp 1666464484
transform 1 0 18676 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_201
timestamp 1666464484
transform 1 0 19596 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_207
timestamp 1666464484
transform 1 0 20148 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_210
timestamp 1666464484
transform 1 0 20424 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1666464484
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666464484
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666464484
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666464484
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666464484
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1666464484
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1666464484
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1666464484
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666464484
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666464484
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1666464484
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1666464484
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1666464484
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1666464484
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1666464484
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1666464484
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1666464484
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1666464484
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1666464484
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1666464484
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1666464484
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1666464484
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1666464484
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666464484
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1666464484
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1666464484
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1666464484
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1666464484
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1666464484
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1666464484
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1666464484
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1666464484
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1666464484
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1666464484
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1666464484
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_617
timestamp 1666464484
transform 1 0 57868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_623
timestamp 1666464484
transform 1 0 58420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_9
timestamp 1666464484
transform 1 0 1932 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1666464484
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_33
timestamp 1666464484
transform 1 0 4140 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_39
timestamp 1666464484
transform 1 0 4692 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_51
timestamp 1666464484
transform 1 0 5796 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_63
timestamp 1666464484
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_75
timestamp 1666464484
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_122
timestamp 1666464484
transform 1 0 12328 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1666464484
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_177
timestamp 1666464484
transform 1 0 17388 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_185
timestamp 1666464484
transform 1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_210
timestamp 1666464484
transform 1 0 20424 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_216
timestamp 1666464484
transform 1 0 20976 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_228
timestamp 1666464484
transform 1 0 22080 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_240
timestamp 1666464484
transform 1 0 23184 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1666464484
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666464484
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666464484
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1666464484
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1666464484
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1666464484
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1666464484
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1666464484
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1666464484
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1666464484
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1666464484
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1666464484
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1666464484
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1666464484
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1666464484
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1666464484
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1666464484
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666464484
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666464484
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666464484
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666464484
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1666464484
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1666464484
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1666464484
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1666464484
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1666464484
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1666464484
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1666464484
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1666464484
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1666464484
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_601
timestamp 1666464484
transform 1 0 56396 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_607
timestamp 1666464484
transform 1 0 56948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_610
timestamp 1666464484
transform 1 0 57224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_616
timestamp 1666464484
transform 1 0 57776 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_623
timestamp 1666464484
transform 1 0 58420 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1666464484
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_21
timestamp 1666464484
transform 1 0 3036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_77
timestamp 1666464484
transform 1 0 8188 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_98
timestamp 1666464484
transform 1 0 10120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1666464484
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_133
timestamp 1666464484
transform 1 0 13340 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_156
timestamp 1666464484
transform 1 0 15456 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_187
timestamp 1666464484
transform 1 0 18308 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_190
timestamp 1666464484
transform 1 0 18584 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_197
timestamp 1666464484
transform 1 0 19228 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_203
timestamp 1666464484
transform 1 0 19780 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_215
timestamp 1666464484
transform 1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666464484
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666464484
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1666464484
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1666464484
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1666464484
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666464484
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1666464484
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1666464484
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1666464484
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666464484
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1666464484
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1666464484
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1666464484
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1666464484
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666464484
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1666464484
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1666464484
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1666464484
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1666464484
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1666464484
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1666464484
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1666464484
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1666464484
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1666464484
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1666464484
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1666464484
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_597
timestamp 1666464484
transform 1 0 56028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_605
timestamp 1666464484
transform 1 0 56764 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_608
timestamp 1666464484
transform 1 0 57040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_614
timestamp 1666464484
transform 1 0 57592 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_617
timestamp 1666464484
transform 1 0 57868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1666464484
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_9
timestamp 1666464484
transform 1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_19
timestamp 1666464484
transform 1 0 2852 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1666464484
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_49
timestamp 1666464484
transform 1 0 5612 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_72
timestamp 1666464484
transform 1 0 7728 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_105
timestamp 1666464484
transform 1 0 10764 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_126
timestamp 1666464484
transform 1 0 12696 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1666464484
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666464484
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1666464484
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_202
timestamp 1666464484
transform 1 0 19688 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_214
timestamp 1666464484
transform 1 0 20792 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_226
timestamp 1666464484
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_238
timestamp 1666464484
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1666464484
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1666464484
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1666464484
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666464484
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1666464484
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1666464484
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1666464484
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1666464484
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1666464484
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666464484
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1666464484
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1666464484
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1666464484
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666464484
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1666464484
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1666464484
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1666464484
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1666464484
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1666464484
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666464484
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666464484
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666464484
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1666464484
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1666464484
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1666464484
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1666464484
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1666464484
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1666464484
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1666464484
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1666464484
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1666464484
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1666464484
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_601
timestamp 1666464484
transform 1 0 56396 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_623
timestamp 1666464484
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_9
timestamp 1666464484
transform 1 0 1932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_22
timestamp 1666464484
transform 1 0 3128 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_28
timestamp 1666464484
transform 1 0 3680 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_34
timestamp 1666464484
transform 1 0 4232 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_46
timestamp 1666464484
transform 1 0 5336 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1666464484
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_62
timestamp 1666464484
transform 1 0 6808 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_68
timestamp 1666464484
transform 1 0 7360 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_80
timestamp 1666464484
transform 1 0 8464 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_92
timestamp 1666464484
transform 1 0 9568 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_100
timestamp 1666464484
transform 1 0 10304 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_104
timestamp 1666464484
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_129
timestamp 1666464484
transform 1 0 12972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_141
timestamp 1666464484
transform 1 0 14076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_153
timestamp 1666464484
transform 1 0 15180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1666464484
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_174
timestamp 1666464484
transform 1 0 17112 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_184
timestamp 1666464484
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_190
timestamp 1666464484
transform 1 0 18584 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_203
timestamp 1666464484
transform 1 0 19780 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_209
timestamp 1666464484
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1666464484
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1666464484
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1666464484
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1666464484
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1666464484
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666464484
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666464484
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666464484
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666464484
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1666464484
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1666464484
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1666464484
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1666464484
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666464484
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1666464484
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1666464484
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1666464484
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1666464484
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666464484
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1666464484
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1666464484
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1666464484
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1666464484
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1666464484
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1666464484
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_597
timestamp 1666464484
transform 1 0 56028 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_605
timestamp 1666464484
transform 1 0 56764 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_608
timestamp 1666464484
transform 1 0 57040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_614
timestamp 1666464484
transform 1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_617
timestamp 1666464484
transform 1 0 57868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1666464484
transform 1 0 58420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_11
timestamp 1666464484
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1666464484
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_33
timestamp 1666464484
transform 1 0 4140 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_39
timestamp 1666464484
transform 1 0 4692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_56
timestamp 1666464484
transform 1 0 6256 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_67
timestamp 1666464484
transform 1 0 7268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_73
timestamp 1666464484
transform 1 0 7820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1666464484
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_102
timestamp 1666464484
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_115
timestamp 1666464484
transform 1 0 11684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_127
timestamp 1666464484
transform 1 0 12788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_169
timestamp 1666464484
transform 1 0 16652 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_182
timestamp 1666464484
transform 1 0 17848 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_188
timestamp 1666464484
transform 1 0 18400 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666464484
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666464484
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666464484
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666464484
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1666464484
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1666464484
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666464484
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666464484
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666464484
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1666464484
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1666464484
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666464484
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666464484
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666464484
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1666464484
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1666464484
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1666464484
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666464484
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666464484
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_457
timestamp 1666464484
transform 1 0 43148 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_465
timestamp 1666464484
transform 1 0 43884 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_470
timestamp 1666464484
transform 1 0 44344 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666464484
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666464484
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666464484
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1666464484
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1666464484
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1666464484
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1666464484
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1666464484
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1666464484
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1666464484
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1666464484
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1666464484
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_601
timestamp 1666464484
transform 1 0 56396 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_607
timestamp 1666464484
transform 1 0 56948 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_610
timestamp 1666464484
transform 1 0 57224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_616
timestamp 1666464484
transform 1 0 57776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_623
timestamp 1666464484
transform 1 0 58420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_7
timestamp 1666464484
transform 1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_20
timestamp 1666464484
transform 1 0 2944 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_26
timestamp 1666464484
transform 1 0 3496 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_29
timestamp 1666464484
transform 1 0 3772 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_36
timestamp 1666464484
transform 1 0 4416 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_44
timestamp 1666464484
transform 1 0 5152 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1666464484
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_61
timestamp 1666464484
transform 1 0 6716 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_67
timestamp 1666464484
transform 1 0 7268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1666464484
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_86
timestamp 1666464484
transform 1 0 9016 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_94
timestamp 1666464484
transform 1 0 9752 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_99
timestamp 1666464484
transform 1 0 10212 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_107
timestamp 1666464484
transform 1 0 10948 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1666464484
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_117
timestamp 1666464484
transform 1 0 11868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1666464484
transform 1 0 12512 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_131
timestamp 1666464484
transform 1 0 13156 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_139
timestamp 1666464484
transform 1 0 13892 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_151
timestamp 1666464484
transform 1 0 14996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_154
timestamp 1666464484
transform 1 0 15272 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_162
timestamp 1666464484
transform 1 0 16008 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1666464484
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_187
timestamp 1666464484
transform 1 0 18308 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_199
timestamp 1666464484
transform 1 0 19412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_211
timestamp 1666464484
transform 1 0 20516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666464484
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666464484
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1666464484
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1666464484
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1666464484
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1666464484
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666464484
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666464484
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666464484
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1666464484
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666464484
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666464484
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666464484
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666464484
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666464484
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1666464484
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1666464484
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1666464484
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666464484
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666464484
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1666464484
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1666464484
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1666464484
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1666464484
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1666464484
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1666464484
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1666464484
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_597
timestamp 1666464484
transform 1 0 56028 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_605
timestamp 1666464484
transform 1 0 56764 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_608
timestamp 1666464484
transform 1 0 57040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_614
timestamp 1666464484
transform 1 0 57592 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_617
timestamp 1666464484
transform 1 0 57868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_623
timestamp 1666464484
transform 1 0 58420 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_9
timestamp 1666464484
transform 1 0 1932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 1666464484
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_33
timestamp 1666464484
transform 1 0 4140 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_47
timestamp 1666464484
transform 1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_59
timestamp 1666464484
transform 1 0 6532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_71
timestamp 1666464484
transform 1 0 7636 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1666464484
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_89
timestamp 1666464484
transform 1 0 9292 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_100
timestamp 1666464484
transform 1 0 10304 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_113
timestamp 1666464484
transform 1 0 11500 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_119
timestamp 1666464484
transform 1 0 12052 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_122
timestamp 1666464484
transform 1 0 12328 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1666464484
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_152
timestamp 1666464484
transform 1 0 15088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_158
timestamp 1666464484
transform 1 0 15640 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_164
timestamp 1666464484
transform 1 0 16192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_168
timestamp 1666464484
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_171
timestamp 1666464484
transform 1 0 16836 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_179
timestamp 1666464484
transform 1 0 17572 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_183
timestamp 1666464484
transform 1 0 17940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666464484
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666464484
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1666464484
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666464484
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1666464484
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1666464484
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1666464484
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1666464484
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666464484
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666464484
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666464484
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666464484
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666464484
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666464484
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666464484
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666464484
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666464484
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666464484
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666464484
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666464484
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666464484
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666464484
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1666464484
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1666464484
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1666464484
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1666464484
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1666464484
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1666464484
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1666464484
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1666464484
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1666464484
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1666464484
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_601
timestamp 1666464484
transform 1 0 56396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_623
timestamp 1666464484
transform 1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_9
timestamp 1666464484
transform 1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_23
timestamp 1666464484
transform 1 0 3220 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_35
timestamp 1666464484
transform 1 0 4324 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_45
timestamp 1666464484
transform 1 0 5244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_61
timestamp 1666464484
transform 1 0 6716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_65
timestamp 1666464484
transform 1 0 7084 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_71
timestamp 1666464484
transform 1 0 7636 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_88
timestamp 1666464484
transform 1 0 9200 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_94
timestamp 1666464484
transform 1 0 9752 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_100
timestamp 1666464484
transform 1 0 10304 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_106
timestamp 1666464484
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_117
timestamp 1666464484
transform 1 0 11868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_127
timestamp 1666464484
transform 1 0 12788 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_157
timestamp 1666464484
transform 1 0 15548 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1666464484
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1666464484
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_186
timestamp 1666464484
transform 1 0 18216 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_198
timestamp 1666464484
transform 1 0 19320 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_210
timestamp 1666464484
transform 1 0 20424 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1666464484
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666464484
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666464484
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666464484
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666464484
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1666464484
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1666464484
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1666464484
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1666464484
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666464484
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666464484
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666464484
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666464484
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666464484
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666464484
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666464484
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666464484
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666464484
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666464484
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666464484
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666464484
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666464484
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666464484
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1666464484
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1666464484
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1666464484
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1666464484
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1666464484
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1666464484
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1666464484
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_597
timestamp 1666464484
transform 1 0 56028 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_602
timestamp 1666464484
transform 1 0 56488 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_608
timestamp 1666464484
transform 1 0 57040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_614
timestamp 1666464484
transform 1 0 57592 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_617
timestamp 1666464484
transform 1 0 57868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_623
timestamp 1666464484
transform 1 0 58420 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_11
timestamp 1666464484
transform 1 0 2116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_23
timestamp 1666464484
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_47
timestamp 1666464484
transform 1 0 5428 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_60
timestamp 1666464484
transform 1 0 6624 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_66
timestamp 1666464484
transform 1 0 7176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_70
timestamp 1666464484
transform 1 0 7544 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_74
timestamp 1666464484
transform 1 0 7912 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1666464484
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_96
timestamp 1666464484
transform 1 0 9936 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_102
timestamp 1666464484
transform 1 0 10488 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_112
timestamp 1666464484
transform 1 0 11408 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_125
timestamp 1666464484
transform 1 0 12604 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_131
timestamp 1666464484
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666464484
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_165
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_169
timestamp 1666464484
transform 1 0 16652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_181
timestamp 1666464484
transform 1 0 17756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1666464484
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666464484
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666464484
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1666464484
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666464484
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666464484
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666464484
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666464484
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666464484
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666464484
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666464484
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666464484
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666464484
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666464484
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666464484
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666464484
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666464484
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666464484
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666464484
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666464484
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666464484
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666464484
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666464484
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1666464484
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1666464484
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1666464484
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1666464484
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1666464484
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1666464484
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1666464484
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1666464484
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_589
timestamp 1666464484
transform 1 0 55292 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_595
timestamp 1666464484
transform 1 0 55844 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_598
timestamp 1666464484
transform 1 0 56120 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_620
timestamp 1666464484
transform 1 0 58144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_624
timestamp 1666464484
transform 1 0 58512 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_9
timestamp 1666464484
transform 1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_61
timestamp 1666464484
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_64
timestamp 1666464484
transform 1 0 6992 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_70
timestamp 1666464484
transform 1 0 7544 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_74
timestamp 1666464484
transform 1 0 7912 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_84
timestamp 1666464484
transform 1 0 8832 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_90
timestamp 1666464484
transform 1 0 9384 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_98
timestamp 1666464484
transform 1 0 10120 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1666464484
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_117
timestamp 1666464484
transform 1 0 11868 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_123
timestamp 1666464484
transform 1 0 12420 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_135
timestamp 1666464484
transform 1 0 13524 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_147
timestamp 1666464484
transform 1 0 14628 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 1666464484
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666464484
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666464484
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666464484
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666464484
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666464484
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666464484
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666464484
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666464484
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666464484
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666464484
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666464484
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666464484
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666464484
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666464484
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666464484
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666464484
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666464484
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666464484
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666464484
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666464484
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666464484
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666464484
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666464484
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666464484
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666464484
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1666464484
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1666464484
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1666464484
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1666464484
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1666464484
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1666464484
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1666464484
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_597
timestamp 1666464484
transform 1 0 56028 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_601
timestamp 1666464484
transform 1 0 56396 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_607
timestamp 1666464484
transform 1 0 56948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_614
timestamp 1666464484
transform 1 0 57592 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_617
timestamp 1666464484
transform 1 0 57868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_623
timestamp 1666464484
transform 1 0 58420 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_9
timestamp 1666464484
transform 1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_89
timestamp 1666464484
transform 1 0 9292 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_95
timestamp 1666464484
transform 1 0 9844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_107
timestamp 1666464484
transform 1 0 10948 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_113
timestamp 1666464484
transform 1 0 11500 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_126
timestamp 1666464484
transform 1 0 12696 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1666464484
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666464484
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666464484
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666464484
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666464484
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666464484
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666464484
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666464484
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666464484
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666464484
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666464484
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666464484
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666464484
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666464484
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666464484
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666464484
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666464484
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666464484
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666464484
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666464484
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666464484
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666464484
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666464484
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1666464484
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1666464484
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1666464484
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1666464484
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1666464484
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1666464484
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1666464484
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1666464484
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_589
timestamp 1666464484
transform 1 0 55292 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_597
timestamp 1666464484
transform 1 0 56028 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_617
timestamp 1666464484
transform 1 0 57868 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_623
timestamp 1666464484
transform 1 0 58420 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1666464484
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_124
timestamp 1666464484
transform 1 0 12512 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_130
timestamp 1666464484
transform 1 0 13064 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_142
timestamp 1666464484
transform 1 0 14168 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_154
timestamp 1666464484
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1666464484
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666464484
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666464484
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666464484
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666464484
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666464484
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666464484
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666464484
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666464484
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666464484
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666464484
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666464484
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666464484
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666464484
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666464484
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666464484
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666464484
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666464484
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666464484
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666464484
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1666464484
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1666464484
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1666464484
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1666464484
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1666464484
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1666464484
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1666464484
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_597
timestamp 1666464484
transform 1 0 56028 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_605
timestamp 1666464484
transform 1 0 56764 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_608
timestamp 1666464484
transform 1 0 57040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_614
timestamp 1666464484
transform 1 0 57592 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_617
timestamp 1666464484
transform 1 0 57868 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_623
timestamp 1666464484
transform 1 0 58420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_9
timestamp 1666464484
transform 1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666464484
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666464484
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666464484
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666464484
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1666464484
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666464484
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666464484
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666464484
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666464484
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666464484
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666464484
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1666464484
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1666464484
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1666464484
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1666464484
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666464484
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666464484
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666464484
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666464484
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666464484
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666464484
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666464484
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666464484
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1666464484
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1666464484
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1666464484
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1666464484
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1666464484
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1666464484
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1666464484
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1666464484
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1666464484
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1666464484
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_613
timestamp 1666464484
transform 1 0 57500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_616
timestamp 1666464484
transform 1 0 57776 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_623
timestamp 1666464484
transform 1 0 58420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_9
timestamp 1666464484
transform 1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666464484
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666464484
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666464484
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666464484
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666464484
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666464484
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1666464484
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1666464484
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1666464484
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1666464484
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666464484
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666464484
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666464484
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666464484
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666464484
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666464484
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666464484
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666464484
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666464484
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666464484
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666464484
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666464484
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666464484
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666464484
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666464484
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666464484
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666464484
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666464484
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666464484
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1666464484
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_561
timestamp 1666464484
transform 1 0 52716 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1666464484
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1666464484
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_599
timestamp 1666464484
transform 1 0 56212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_611
timestamp 1666464484
transform 1 0 57316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_614
timestamp 1666464484
transform 1 0 57592 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_617
timestamp 1666464484
transform 1 0 57868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1666464484
transform 1 0 58420 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666464484
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666464484
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666464484
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666464484
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666464484
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666464484
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666464484
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1666464484
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1666464484
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1666464484
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666464484
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666464484
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666464484
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666464484
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666464484
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666464484
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666464484
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666464484
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666464484
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666464484
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666464484
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666464484
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666464484
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666464484
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1666464484
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1666464484
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1666464484
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1666464484
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1666464484
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1666464484
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1666464484
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1666464484
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_589
timestamp 1666464484
transform 1 0 55292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_595
timestamp 1666464484
transform 1 0 55844 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_620
timestamp 1666464484
transform 1 0 58144 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_624
timestamp 1666464484
transform 1 0 58512 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_9
timestamp 1666464484
transform 1 0 1932 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666464484
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666464484
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666464484
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666464484
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666464484
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1666464484
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1666464484
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1666464484
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666464484
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666464484
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666464484
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1666464484
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666464484
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666464484
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666464484
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666464484
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666464484
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1666464484
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666464484
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666464484
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666464484
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666464484
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666464484
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666464484
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666464484
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666464484
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666464484
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666464484
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666464484
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1666464484
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1666464484
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1666464484
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1666464484
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_597
timestamp 1666464484
transform 1 0 56028 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_600
timestamp 1666464484
transform 1 0 56304 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_614
timestamp 1666464484
transform 1 0 57592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_617
timestamp 1666464484
transform 1 0 57868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_623
timestamp 1666464484
transform 1 0 58420 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_9
timestamp 1666464484
transform 1 0 1932 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666464484
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666464484
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666464484
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666464484
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666464484
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666464484
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666464484
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666464484
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666464484
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666464484
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666464484
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666464484
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666464484
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666464484
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666464484
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666464484
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666464484
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666464484
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1666464484
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1666464484
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1666464484
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666464484
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666464484
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666464484
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666464484
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1666464484
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1666464484
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1666464484
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1666464484
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1666464484
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1666464484
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1666464484
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1666464484
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_589
timestamp 1666464484
transform 1 0 55292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_593
timestamp 1666464484
transform 1 0 55660 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_596
timestamp 1666464484
transform 1 0 55936 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_618
timestamp 1666464484
transform 1 0 57960 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_624
timestamp 1666464484
transform 1 0 58512 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666464484
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666464484
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666464484
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666464484
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666464484
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666464484
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666464484
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666464484
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1666464484
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1666464484
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1666464484
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1666464484
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666464484
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1666464484
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1666464484
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1666464484
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1666464484
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666464484
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1666464484
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666464484
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666464484
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1666464484
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666464484
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666464484
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666464484
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666464484
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666464484
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666464484
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666464484
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666464484
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666464484
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666464484
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1666464484
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1666464484
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_573
timestamp 1666464484
transform 1 0 53820 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_587
timestamp 1666464484
transform 1 0 55108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_599
timestamp 1666464484
transform 1 0 56212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_611
timestamp 1666464484
transform 1 0 57316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_614
timestamp 1666464484
transform 1 0 57592 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_617
timestamp 1666464484
transform 1 0 57868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_623
timestamp 1666464484
transform 1 0 58420 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_9
timestamp 1666464484
transform 1 0 1932 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666464484
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1666464484
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1666464484
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666464484
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1666464484
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1666464484
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1666464484
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1666464484
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666464484
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1666464484
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1666464484
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1666464484
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1666464484
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666464484
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666464484
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1666464484
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1666464484
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1666464484
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666464484
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666464484
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666464484
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666464484
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666464484
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666464484
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666464484
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666464484
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666464484
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666464484
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666464484
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666464484
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666464484
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666464484
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1666464484
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1666464484
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1666464484
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1666464484
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_569
timestamp 1666464484
transform 1 0 53452 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_579
timestamp 1666464484
transform 1 0 54372 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1666464484
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1666464484
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_601
timestamp 1666464484
transform 1 0 56396 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_607
timestamp 1666464484
transform 1 0 56948 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_610
timestamp 1666464484
transform 1 0 57224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_616
timestamp 1666464484
transform 1 0 57776 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_623
timestamp 1666464484
transform 1 0 58420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1666464484
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666464484
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666464484
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666464484
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666464484
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1666464484
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666464484
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1666464484
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1666464484
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666464484
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1666464484
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666464484
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666464484
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1666464484
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1666464484
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1666464484
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666464484
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1666464484
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666464484
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666464484
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1666464484
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666464484
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666464484
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666464484
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666464484
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666464484
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666464484
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666464484
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666464484
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666464484
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666464484
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1666464484
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_547
timestamp 1666464484
transform 1 0 51428 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_558
timestamp 1666464484
transform 1 0 52440 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1666464484
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_575
timestamp 1666464484
transform 1 0 54004 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_600
timestamp 1666464484
transform 1 0 56304 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_606
timestamp 1666464484
transform 1 0 56856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_614
timestamp 1666464484
transform 1 0 57592 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_617
timestamp 1666464484
transform 1 0 57868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1666464484
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666464484
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666464484
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666464484
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666464484
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1666464484
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1666464484
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666464484
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1666464484
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1666464484
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1666464484
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1666464484
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666464484
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1666464484
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1666464484
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1666464484
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1666464484
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666464484
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666464484
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666464484
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1666464484
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1666464484
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666464484
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1666464484
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1666464484
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1666464484
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1666464484
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666464484
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666464484
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666464484
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666464484
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666464484
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666464484
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666464484
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666464484
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666464484
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1666464484
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1666464484
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1666464484
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1666464484
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1666464484
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1666464484
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1666464484
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1666464484
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1666464484
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_589
timestamp 1666464484
transform 1 0 55292 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_593
timestamp 1666464484
transform 1 0 55660 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_596
timestamp 1666464484
transform 1 0 55936 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1666464484
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1666464484
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666464484
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666464484
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666464484
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666464484
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666464484
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1666464484
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1666464484
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666464484
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1666464484
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1666464484
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1666464484
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1666464484
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1666464484
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1666464484
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1666464484
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1666464484
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1666464484
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666464484
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1666464484
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1666464484
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1666464484
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1666464484
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666464484
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666464484
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666464484
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666464484
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666464484
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666464484
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666464484
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666464484
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666464484
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666464484
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1666464484
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1666464484
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1666464484
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1666464484
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1666464484
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1666464484
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1666464484
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_597
timestamp 1666464484
transform 1 0 56028 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_600
timestamp 1666464484
transform 1 0 56304 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_608
timestamp 1666464484
transform 1 0 57040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_614
timestamp 1666464484
transform 1 0 57592 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_617
timestamp 1666464484
transform 1 0 57868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_623
timestamp 1666464484
transform 1 0 58420 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1666464484
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666464484
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666464484
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666464484
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666464484
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1666464484
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666464484
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666464484
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1666464484
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1666464484
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1666464484
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1666464484
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666464484
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1666464484
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1666464484
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1666464484
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1666464484
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666464484
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1666464484
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1666464484
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1666464484
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1666464484
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666464484
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666464484
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1666464484
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1666464484
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1666464484
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666464484
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666464484
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666464484
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666464484
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666464484
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666464484
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666464484
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666464484
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666464484
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1666464484
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1666464484
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1666464484
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1666464484
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1666464484
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1666464484
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1666464484
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1666464484
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_589
timestamp 1666464484
transform 1 0 55292 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_597
timestamp 1666464484
transform 1 0 56028 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_601
timestamp 1666464484
transform 1 0 56396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_623
timestamp 1666464484
transform 1 0 58420 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666464484
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666464484
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666464484
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666464484
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666464484
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666464484
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666464484
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666464484
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666464484
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666464484
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666464484
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666464484
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1666464484
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1666464484
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666464484
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1666464484
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1666464484
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1666464484
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1666464484
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1666464484
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1666464484
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1666464484
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1666464484
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1666464484
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1666464484
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1666464484
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666464484
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666464484
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1666464484
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666464484
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666464484
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666464484
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666464484
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666464484
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666464484
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666464484
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666464484
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666464484
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666464484
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666464484
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1666464484
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1666464484
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1666464484
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1666464484
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1666464484
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1666464484
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1666464484
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_597
timestamp 1666464484
transform 1 0 56028 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_605
timestamp 1666464484
transform 1 0 56764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_611
timestamp 1666464484
transform 1 0 57316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_614
timestamp 1666464484
transform 1 0 57592 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_617
timestamp 1666464484
transform 1 0 57868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_623
timestamp 1666464484
transform 1 0 58420 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1666464484
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666464484
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666464484
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666464484
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666464484
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666464484
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666464484
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666464484
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666464484
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666464484
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666464484
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666464484
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666464484
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666464484
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666464484
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666464484
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666464484
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1666464484
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1666464484
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1666464484
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666464484
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1666464484
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1666464484
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1666464484
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1666464484
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666464484
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1666464484
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1666464484
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1666464484
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1666464484
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666464484
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1666464484
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1666464484
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1666464484
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1666464484
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666464484
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666464484
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666464484
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666464484
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666464484
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666464484
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666464484
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666464484
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666464484
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1666464484
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1666464484
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1666464484
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1666464484
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1666464484
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1666464484
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_569
timestamp 1666464484
transform 1 0 53452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_579
timestamp 1666464484
transform 1 0 54372 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1666464484
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1666464484
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_601
timestamp 1666464484
transform 1 0 56396 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_607
timestamp 1666464484
transform 1 0 56948 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_610
timestamp 1666464484
transform 1 0 57224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_616
timestamp 1666464484
transform 1 0 57776 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_623
timestamp 1666464484
transform 1 0 58420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_9
timestamp 1666464484
transform 1 0 1932 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666464484
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666464484
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666464484
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1666464484
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1666464484
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666464484
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666464484
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666464484
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666464484
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666464484
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666464484
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666464484
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666464484
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666464484
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1666464484
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1666464484
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666464484
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666464484
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666464484
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666464484
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1666464484
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1666464484
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666464484
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1666464484
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1666464484
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1666464484
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1666464484
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1666464484
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666464484
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1666464484
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1666464484
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1666464484
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1666464484
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1666464484
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666464484
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1666464484
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1666464484
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1666464484
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1666464484
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1666464484
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666464484
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666464484
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666464484
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666464484
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666464484
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666464484
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666464484
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666464484
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666464484
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666464484
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666464484
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666464484
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666464484
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1666464484
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1666464484
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1666464484
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1666464484
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1666464484
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1666464484
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1666464484
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_575
timestamp 1666464484
transform 1 0 54004 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_597
timestamp 1666464484
transform 1 0 56028 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_603
timestamp 1666464484
transform 1 0 56580 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1666464484
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_617
timestamp 1666464484
transform 1 0 57868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_623
timestamp 1666464484
transform 1 0 58420 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666464484
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666464484
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666464484
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666464484
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666464484
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666464484
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666464484
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666464484
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666464484
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666464484
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666464484
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666464484
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666464484
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666464484
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666464484
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666464484
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666464484
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1666464484
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1666464484
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666464484
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1666464484
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1666464484
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1666464484
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1666464484
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1666464484
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1666464484
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1666464484
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1666464484
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1666464484
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1666464484
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1666464484
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1666464484
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1666464484
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1666464484
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1666464484
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1666464484
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1666464484
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666464484
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666464484
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1666464484
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1666464484
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666464484
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1666464484
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666464484
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666464484
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666464484
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666464484
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666464484
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666464484
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666464484
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666464484
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666464484
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666464484
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1666464484
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1666464484
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1666464484
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1666464484
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1666464484
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1666464484
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1666464484
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1666464484
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_589
timestamp 1666464484
transform 1 0 55292 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_595
timestamp 1666464484
transform 1 0 55844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_609
timestamp 1666464484
transform 1 0 57132 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_615
timestamp 1666464484
transform 1 0 57684 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_623
timestamp 1666464484
transform 1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_9
timestamp 1666464484
transform 1 0 1932 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666464484
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666464484
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1666464484
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1666464484
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1666464484
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666464484
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666464484
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666464484
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666464484
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666464484
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666464484
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666464484
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666464484
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666464484
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1666464484
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1666464484
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1666464484
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666464484
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666464484
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1666464484
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1666464484
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666464484
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1666464484
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1666464484
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1666464484
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1666464484
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1666464484
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1666464484
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1666464484
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1666464484
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1666464484
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1666464484
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1666464484
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666464484
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1666464484
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1666464484
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666464484
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666464484
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1666464484
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1666464484
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666464484
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666464484
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666464484
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666464484
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666464484
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666464484
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666464484
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666464484
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666464484
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666464484
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666464484
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666464484
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1666464484
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1666464484
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1666464484
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1666464484
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1666464484
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1666464484
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1666464484
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1666464484
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_585
timestamp 1666464484
transform 1 0 54924 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_591
timestamp 1666464484
transform 1 0 55476 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_613
timestamp 1666464484
transform 1 0 57500 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_617
timestamp 1666464484
transform 1 0 57868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_623
timestamp 1666464484
transform 1 0 58420 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_9
timestamp 1666464484
transform 1 0 1932 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666464484
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666464484
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666464484
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666464484
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666464484
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666464484
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666464484
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666464484
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666464484
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666464484
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666464484
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666464484
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666464484
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666464484
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666464484
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666464484
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1666464484
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1666464484
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1666464484
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666464484
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666464484
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666464484
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1666464484
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1666464484
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1666464484
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666464484
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1666464484
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1666464484
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1666464484
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1666464484
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666464484
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666464484
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1666464484
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1666464484
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1666464484
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1666464484
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1666464484
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666464484
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1666464484
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666464484
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1666464484
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1666464484
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1666464484
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666464484
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666464484
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666464484
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666464484
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666464484
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666464484
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666464484
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666464484
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666464484
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666464484
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1666464484
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1666464484
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1666464484
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1666464484
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1666464484
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1666464484
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1666464484
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1666464484
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1666464484
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_589
timestamp 1666464484
transform 1 0 55292 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_599
timestamp 1666464484
transform 1 0 56212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_621
timestamp 1666464484
transform 1 0 58236 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666464484
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1666464484
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1666464484
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666464484
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666464484
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666464484
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666464484
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666464484
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666464484
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666464484
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666464484
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666464484
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666464484
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666464484
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666464484
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666464484
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666464484
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666464484
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666464484
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666464484
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666464484
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666464484
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1666464484
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1666464484
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1666464484
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1666464484
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1666464484
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1666464484
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1666464484
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1666464484
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1666464484
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1666464484
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1666464484
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666464484
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1666464484
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1666464484
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666464484
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666464484
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1666464484
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666464484
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666464484
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666464484
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666464484
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666464484
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666464484
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666464484
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666464484
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666464484
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666464484
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666464484
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666464484
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666464484
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1666464484
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1666464484
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1666464484
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1666464484
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1666464484
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1666464484
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1666464484
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1666464484
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1666464484
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_597
timestamp 1666464484
transform 1 0 56028 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_603
timestamp 1666464484
transform 1 0 56580 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_611
timestamp 1666464484
transform 1 0 57316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_614
timestamp 1666464484
transform 1 0 57592 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_617
timestamp 1666464484
transform 1 0 57868 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_623
timestamp 1666464484
transform 1 0 58420 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_9
timestamp 1666464484
transform 1 0 1932 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666464484
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666464484
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666464484
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666464484
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666464484
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666464484
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666464484
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666464484
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666464484
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666464484
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666464484
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666464484
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666464484
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666464484
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666464484
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666464484
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666464484
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1666464484
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1666464484
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666464484
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666464484
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666464484
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1666464484
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1666464484
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1666464484
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1666464484
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1666464484
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1666464484
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1666464484
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1666464484
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1666464484
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666464484
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1666464484
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1666464484
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1666464484
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1666464484
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1666464484
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666464484
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1666464484
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1666464484
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1666464484
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1666464484
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1666464484
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666464484
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666464484
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666464484
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666464484
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666464484
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666464484
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666464484
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666464484
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666464484
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666464484
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1666464484
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1666464484
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1666464484
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1666464484
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1666464484
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1666464484
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1666464484
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1666464484
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1666464484
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1666464484
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1666464484
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_613
timestamp 1666464484
transform 1 0 57500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_616
timestamp 1666464484
transform 1 0 57776 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_623
timestamp 1666464484
transform 1 0 58420 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_9
timestamp 1666464484
transform 1 0 1932 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666464484
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1666464484
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1666464484
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666464484
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666464484
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666464484
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666464484
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666464484
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666464484
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666464484
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666464484
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666464484
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666464484
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666464484
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666464484
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666464484
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666464484
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666464484
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666464484
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666464484
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1666464484
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666464484
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1666464484
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1666464484
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1666464484
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1666464484
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1666464484
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1666464484
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1666464484
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1666464484
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1666464484
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1666464484
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1666464484
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1666464484
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1666464484
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1666464484
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1666464484
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1666464484
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1666464484
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666464484
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666464484
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666464484
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666464484
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666464484
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666464484
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666464484
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666464484
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666464484
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666464484
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666464484
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666464484
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666464484
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1666464484
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1666464484
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1666464484
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1666464484
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1666464484
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1666464484
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1666464484
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1666464484
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1666464484
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1666464484
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1666464484
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1666464484
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_617
timestamp 1666464484
transform 1 0 57868 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_623
timestamp 1666464484
transform 1 0 58420 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666464484
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666464484
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666464484
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666464484
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666464484
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666464484
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666464484
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666464484
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666464484
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666464484
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666464484
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666464484
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666464484
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666464484
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666464484
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666464484
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666464484
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666464484
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666464484
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666464484
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666464484
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1666464484
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1666464484
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1666464484
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1666464484
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1666464484
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1666464484
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1666464484
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1666464484
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1666464484
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1666464484
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1666464484
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1666464484
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1666464484
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1666464484
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1666464484
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1666464484
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1666464484
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1666464484
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1666464484
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1666464484
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1666464484
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1666464484
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1666464484
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666464484
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666464484
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666464484
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666464484
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666464484
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666464484
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666464484
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666464484
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666464484
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1666464484
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1666464484
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1666464484
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1666464484
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1666464484
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1666464484
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1666464484
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1666464484
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1666464484
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1666464484
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_613
timestamp 1666464484
transform 1 0 57500 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_623
timestamp 1666464484
transform 1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_9
timestamp 1666464484
transform 1 0 1932 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666464484
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666464484
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1666464484
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1666464484
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666464484
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666464484
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666464484
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666464484
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666464484
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666464484
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666464484
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666464484
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666464484
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666464484
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666464484
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666464484
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666464484
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666464484
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666464484
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666464484
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666464484
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1666464484
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666464484
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1666464484
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1666464484
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1666464484
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1666464484
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1666464484
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1666464484
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1666464484
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1666464484
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1666464484
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1666464484
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1666464484
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1666464484
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1666464484
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1666464484
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1666464484
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1666464484
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1666464484
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1666464484
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1666464484
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1666464484
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1666464484
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1666464484
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1666464484
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666464484
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666464484
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666464484
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666464484
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666464484
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666464484
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666464484
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1666464484
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1666464484
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1666464484
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1666464484
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1666464484
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1666464484
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1666464484
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1666464484
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1666464484
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1666464484
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_609
timestamp 1666464484
transform 1 0 57132 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_614
timestamp 1666464484
transform 1 0 57592 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_617
timestamp 1666464484
transform 1 0 57868 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_623
timestamp 1666464484
transform 1 0 58420 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_9
timestamp 1666464484
transform 1 0 1932 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666464484
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666464484
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666464484
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666464484
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666464484
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666464484
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666464484
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666464484
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666464484
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666464484
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666464484
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666464484
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666464484
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666464484
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666464484
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666464484
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666464484
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666464484
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666464484
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666464484
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666464484
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666464484
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1666464484
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1666464484
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1666464484
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1666464484
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1666464484
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1666464484
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1666464484
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1666464484
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1666464484
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1666464484
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1666464484
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1666464484
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1666464484
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1666464484
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1666464484
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1666464484
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1666464484
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1666464484
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1666464484
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1666464484
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1666464484
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1666464484
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666464484
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666464484
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666464484
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666464484
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666464484
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666464484
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666464484
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666464484
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666464484
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1666464484
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1666464484
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1666464484
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1666464484
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1666464484
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1666464484
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1666464484
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1666464484
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1666464484
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1666464484
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1666464484
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_613
timestamp 1666464484
transform 1 0 57500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_616
timestamp 1666464484
transform 1 0 57776 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_623
timestamp 1666464484
transform 1 0 58420 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666464484
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666464484
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1666464484
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1666464484
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1666464484
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666464484
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666464484
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666464484
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666464484
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666464484
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666464484
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666464484
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666464484
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666464484
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666464484
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666464484
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666464484
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666464484
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666464484
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666464484
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1666464484
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1666464484
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666464484
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1666464484
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1666464484
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1666464484
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1666464484
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1666464484
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1666464484
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1666464484
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1666464484
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1666464484
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1666464484
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1666464484
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1666464484
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1666464484
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1666464484
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1666464484
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1666464484
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1666464484
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1666464484
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1666464484
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1666464484
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1666464484
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1666464484
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1666464484
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1666464484
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666464484
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666464484
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666464484
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666464484
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666464484
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666464484
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1666464484
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1666464484
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1666464484
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1666464484
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1666464484
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1666464484
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1666464484
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1666464484
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1666464484
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1666464484
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1666464484
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1666464484
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_9
timestamp 1666464484
transform 1 0 1932 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666464484
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666464484
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666464484
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666464484
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666464484
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666464484
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666464484
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666464484
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666464484
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666464484
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666464484
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666464484
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666464484
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666464484
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666464484
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666464484
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666464484
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666464484
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666464484
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1666464484
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1666464484
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1666464484
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1666464484
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1666464484
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1666464484
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1666464484
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1666464484
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1666464484
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1666464484
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1666464484
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1666464484
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1666464484
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1666464484
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1666464484
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1666464484
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1666464484
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1666464484
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1666464484
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1666464484
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1666464484
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1666464484
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1666464484
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1666464484
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1666464484
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1666464484
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1666464484
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1666464484
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1666464484
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666464484
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666464484
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666464484
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666464484
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1666464484
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1666464484
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1666464484
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1666464484
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1666464484
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1666464484
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1666464484
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1666464484
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1666464484
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1666464484
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1666464484
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_613
timestamp 1666464484
transform 1 0 57500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_616
timestamp 1666464484
transform 1 0 57776 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_623
timestamp 1666464484
transform 1 0 58420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_9
timestamp 1666464484
transform 1 0 1932 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666464484
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666464484
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1666464484
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1666464484
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1666464484
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666464484
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666464484
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666464484
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666464484
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666464484
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666464484
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666464484
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666464484
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666464484
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666464484
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666464484
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666464484
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666464484
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666464484
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1666464484
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1666464484
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1666464484
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666464484
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1666464484
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1666464484
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1666464484
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1666464484
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1666464484
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1666464484
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1666464484
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1666464484
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1666464484
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1666464484
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1666464484
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1666464484
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1666464484
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1666464484
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1666464484
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1666464484
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1666464484
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1666464484
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1666464484
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1666464484
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1666464484
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1666464484
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1666464484
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1666464484
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1666464484
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1666464484
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1666464484
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1666464484
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1666464484
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666464484
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1666464484
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1666464484
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1666464484
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1666464484
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1666464484
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1666464484
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1666464484
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1666464484
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1666464484
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1666464484
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1666464484
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1666464484
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_617
timestamp 1666464484
transform 1 0 57868 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_623
timestamp 1666464484
transform 1 0 58420 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666464484
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666464484
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666464484
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666464484
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666464484
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666464484
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666464484
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666464484
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666464484
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666464484
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666464484
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666464484
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666464484
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666464484
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666464484
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666464484
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666464484
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666464484
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1666464484
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1666464484
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1666464484
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1666464484
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1666464484
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1666464484
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1666464484
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1666464484
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1666464484
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1666464484
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1666464484
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1666464484
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1666464484
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1666464484
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1666464484
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1666464484
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1666464484
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1666464484
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1666464484
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1666464484
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1666464484
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1666464484
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1666464484
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1666464484
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1666464484
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1666464484
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1666464484
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1666464484
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1666464484
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1666464484
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1666464484
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1666464484
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666464484
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666464484
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666464484
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1666464484
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1666464484
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1666464484
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1666464484
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1666464484
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1666464484
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1666464484
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1666464484
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1666464484
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1666464484
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_613
timestamp 1666464484
transform 1 0 57500 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_623
timestamp 1666464484
transform 1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_9
timestamp 1666464484
transform 1 0 1932 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666464484
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666464484
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666464484
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1666464484
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1666464484
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666464484
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666464484
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666464484
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666464484
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666464484
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666464484
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666464484
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666464484
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666464484
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666464484
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666464484
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666464484
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1666464484
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1666464484
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1666464484
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1666464484
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1666464484
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1666464484
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1666464484
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1666464484
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1666464484
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1666464484
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1666464484
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1666464484
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1666464484
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1666464484
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1666464484
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1666464484
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1666464484
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1666464484
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1666464484
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1666464484
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1666464484
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1666464484
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1666464484
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1666464484
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1666464484
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1666464484
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1666464484
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1666464484
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1666464484
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1666464484
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1666464484
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1666464484
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1666464484
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1666464484
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1666464484
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1666464484
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1666464484
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1666464484
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1666464484
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1666464484
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1666464484
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1666464484
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1666464484
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1666464484
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1666464484
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1666464484
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_609
timestamp 1666464484
transform 1 0 57132 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_614
timestamp 1666464484
transform 1 0 57592 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_617
timestamp 1666464484
transform 1 0 57868 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_623
timestamp 1666464484
transform 1 0 58420 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_9
timestamp 1666464484
transform 1 0 1932 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666464484
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666464484
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666464484
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1666464484
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1666464484
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666464484
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1666464484
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666464484
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666464484
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666464484
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666464484
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666464484
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666464484
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666464484
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666464484
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666464484
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1666464484
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1666464484
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1666464484
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1666464484
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1666464484
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1666464484
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1666464484
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1666464484
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1666464484
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1666464484
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1666464484
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1666464484
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1666464484
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1666464484
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1666464484
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1666464484
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1666464484
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1666464484
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1666464484
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1666464484
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1666464484
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1666464484
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1666464484
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1666464484
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1666464484
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1666464484
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1666464484
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1666464484
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1666464484
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1666464484
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1666464484
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1666464484
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1666464484
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1666464484
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1666464484
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1666464484
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1666464484
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1666464484
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1666464484
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1666464484
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1666464484
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1666464484
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1666464484
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1666464484
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1666464484
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1666464484
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1666464484
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_613
timestamp 1666464484
transform 1 0 57500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_616
timestamp 1666464484
transform 1 0 57776 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_623
timestamp 1666464484
transform 1 0 58420 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666464484
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1666464484
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666464484
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1666464484
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1666464484
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1666464484
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1666464484
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1666464484
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1666464484
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666464484
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666464484
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1666464484
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1666464484
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1666464484
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666464484
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1666464484
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1666464484
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1666464484
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1666464484
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1666464484
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1666464484
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1666464484
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1666464484
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1666464484
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1666464484
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1666464484
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1666464484
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1666464484
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1666464484
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1666464484
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1666464484
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1666464484
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1666464484
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1666464484
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1666464484
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1666464484
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1666464484
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1666464484
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666464484
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1666464484
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1666464484
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1666464484
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1666464484
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1666464484
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666464484
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1666464484
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1666464484
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1666464484
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1666464484
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1666464484
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1666464484
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1666464484
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1666464484
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1666464484
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1666464484
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1666464484
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1666464484
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1666464484
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1666464484
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1666464484
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1666464484
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1666464484
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1666464484
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1666464484
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_9
timestamp 1666464484
transform 1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666464484
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666464484
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1666464484
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1666464484
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1666464484
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1666464484
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1666464484
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1666464484
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1666464484
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1666464484
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1666464484
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1666464484
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1666464484
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1666464484
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1666464484
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1666464484
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1666464484
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1666464484
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1666464484
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1666464484
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1666464484
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1666464484
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1666464484
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1666464484
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1666464484
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1666464484
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1666464484
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1666464484
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1666464484
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1666464484
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1666464484
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1666464484
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1666464484
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1666464484
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1666464484
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1666464484
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1666464484
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666464484
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1666464484
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1666464484
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1666464484
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1666464484
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1666464484
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1666464484
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1666464484
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1666464484
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1666464484
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1666464484
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1666464484
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1666464484
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1666464484
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1666464484
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1666464484
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1666464484
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1666464484
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1666464484
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1666464484
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1666464484
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1666464484
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1666464484
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1666464484
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1666464484
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1666464484
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1666464484
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_613
timestamp 1666464484
transform 1 0 57500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_616
timestamp 1666464484
transform 1 0 57776 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_623
timestamp 1666464484
transform 1 0 58420 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_9
timestamp 1666464484
transform 1 0 1932 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1666464484
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1666464484
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1666464484
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1666464484
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1666464484
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1666464484
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1666464484
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1666464484
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1666464484
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1666464484
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1666464484
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1666464484
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1666464484
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1666464484
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1666464484
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1666464484
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1666464484
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1666464484
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1666464484
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1666464484
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1666464484
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1666464484
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1666464484
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1666464484
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1666464484
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1666464484
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1666464484
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1666464484
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1666464484
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1666464484
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1666464484
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1666464484
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1666464484
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1666464484
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1666464484
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1666464484
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1666464484
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1666464484
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1666464484
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1666464484
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1666464484
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1666464484
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1666464484
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1666464484
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1666464484
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1666464484
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1666464484
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1666464484
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1666464484
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1666464484
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1666464484
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1666464484
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1666464484
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1666464484
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1666464484
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1666464484
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1666464484
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1666464484
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1666464484
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1666464484
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1666464484
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1666464484
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1666464484
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1666464484
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1666464484
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_617
timestamp 1666464484
transform 1 0 57868 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_623
timestamp 1666464484
transform 1 0 58420 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1666464484
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1666464484
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1666464484
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1666464484
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1666464484
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1666464484
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1666464484
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1666464484
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1666464484
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1666464484
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1666464484
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1666464484
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1666464484
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1666464484
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1666464484
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1666464484
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1666464484
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1666464484
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1666464484
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1666464484
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1666464484
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1666464484
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1666464484
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1666464484
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1666464484
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1666464484
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1666464484
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1666464484
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1666464484
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1666464484
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1666464484
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1666464484
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1666464484
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1666464484
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1666464484
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1666464484
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1666464484
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1666464484
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1666464484
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1666464484
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1666464484
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1666464484
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1666464484
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1666464484
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1666464484
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1666464484
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1666464484
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1666464484
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1666464484
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1666464484
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1666464484
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1666464484
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1666464484
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1666464484
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1666464484
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1666464484
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1666464484
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1666464484
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1666464484
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1666464484
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1666464484
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1666464484
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1666464484
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_613
timestamp 1666464484
transform 1 0 57500 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_623
timestamp 1666464484
transform 1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_9
timestamp 1666464484
transform 1 0 1932 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1666464484
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1666464484
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1666464484
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1666464484
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1666464484
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1666464484
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1666464484
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1666464484
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1666464484
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1666464484
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1666464484
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1666464484
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1666464484
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1666464484
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1666464484
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1666464484
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1666464484
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1666464484
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1666464484
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1666464484
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1666464484
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1666464484
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1666464484
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1666464484
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1666464484
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1666464484
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1666464484
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1666464484
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1666464484
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1666464484
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1666464484
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1666464484
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1666464484
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1666464484
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1666464484
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1666464484
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1666464484
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1666464484
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1666464484
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1666464484
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1666464484
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1666464484
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1666464484
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1666464484
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1666464484
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1666464484
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1666464484
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1666464484
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1666464484
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1666464484
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1666464484
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1666464484
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1666464484
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1666464484
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1666464484
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1666464484
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1666464484
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1666464484
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1666464484
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1666464484
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1666464484
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1666464484
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_609
timestamp 1666464484
transform 1 0 57132 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_614
timestamp 1666464484
transform 1 0 57592 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_85_617
timestamp 1666464484
transform 1 0 57868 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_623
timestamp 1666464484
transform 1 0 58420 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_9
timestamp 1666464484
transform 1 0 1932 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1666464484
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1666464484
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1666464484
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1666464484
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1666464484
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1666464484
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1666464484
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1666464484
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1666464484
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1666464484
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1666464484
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1666464484
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1666464484
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1666464484
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1666464484
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1666464484
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1666464484
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1666464484
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1666464484
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1666464484
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1666464484
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1666464484
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1666464484
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1666464484
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1666464484
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1666464484
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1666464484
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1666464484
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1666464484
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1666464484
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1666464484
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1666464484
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1666464484
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1666464484
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1666464484
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1666464484
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1666464484
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1666464484
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1666464484
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1666464484
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1666464484
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1666464484
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1666464484
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1666464484
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1666464484
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1666464484
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1666464484
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1666464484
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1666464484
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1666464484
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1666464484
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1666464484
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1666464484
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1666464484
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1666464484
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1666464484
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1666464484
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1666464484
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1666464484
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1666464484
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1666464484
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1666464484
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_613
timestamp 1666464484
transform 1 0 57500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_616
timestamp 1666464484
transform 1 0 57776 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_623
timestamp 1666464484
transform 1 0 58420 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1666464484
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1666464484
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1666464484
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1666464484
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1666464484
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1666464484
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1666464484
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1666464484
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1666464484
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1666464484
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1666464484
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1666464484
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1666464484
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1666464484
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1666464484
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1666464484
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1666464484
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1666464484
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1666464484
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1666464484
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1666464484
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1666464484
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1666464484
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1666464484
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1666464484
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1666464484
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1666464484
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1666464484
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1666464484
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1666464484
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1666464484
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1666464484
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1666464484
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1666464484
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1666464484
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1666464484
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1666464484
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1666464484
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1666464484
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1666464484
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1666464484
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1666464484
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1666464484
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1666464484
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1666464484
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1666464484
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1666464484
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1666464484
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1666464484
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1666464484
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1666464484
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1666464484
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1666464484
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1666464484
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1666464484
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1666464484
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1666464484
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1666464484
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1666464484
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1666464484
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1666464484
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1666464484
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1666464484
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_9
timestamp 1666464484
transform 1 0 1932 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1666464484
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1666464484
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1666464484
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1666464484
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1666464484
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1666464484
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1666464484
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1666464484
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1666464484
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1666464484
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1666464484
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1666464484
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1666464484
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1666464484
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1666464484
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1666464484
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1666464484
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1666464484
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1666464484
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1666464484
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1666464484
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1666464484
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1666464484
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1666464484
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1666464484
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1666464484
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1666464484
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1666464484
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1666464484
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1666464484
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1666464484
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1666464484
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1666464484
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1666464484
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1666464484
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1666464484
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1666464484
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1666464484
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1666464484
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1666464484
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1666464484
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1666464484
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1666464484
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1666464484
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1666464484
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1666464484
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1666464484
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1666464484
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1666464484
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1666464484
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1666464484
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1666464484
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1666464484
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1666464484
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1666464484
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1666464484
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1666464484
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1666464484
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1666464484
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1666464484
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1666464484
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1666464484
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1666464484
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_613
timestamp 1666464484
transform 1 0 57500 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_616
timestamp 1666464484
transform 1 0 57776 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_623
timestamp 1666464484
transform 1 0 58420 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_9
timestamp 1666464484
transform 1 0 1932 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1666464484
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1666464484
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1666464484
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1666464484
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1666464484
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1666464484
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1666464484
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1666464484
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1666464484
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1666464484
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1666464484
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1666464484
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1666464484
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1666464484
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1666464484
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1666464484
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1666464484
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1666464484
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1666464484
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1666464484
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1666464484
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1666464484
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1666464484
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1666464484
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1666464484
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1666464484
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1666464484
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1666464484
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1666464484
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1666464484
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1666464484
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1666464484
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1666464484
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1666464484
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1666464484
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1666464484
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1666464484
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1666464484
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1666464484
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1666464484
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1666464484
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1666464484
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1666464484
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1666464484
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1666464484
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1666464484
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1666464484
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1666464484
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1666464484
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1666464484
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1666464484
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1666464484
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1666464484
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1666464484
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1666464484
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1666464484
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1666464484
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1666464484
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1666464484
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1666464484
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1666464484
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1666464484
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1666464484
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_89_617
timestamp 1666464484
transform 1 0 57868 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_623
timestamp 1666464484
transform 1 0 58420 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1666464484
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1666464484
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1666464484
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1666464484
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1666464484
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1666464484
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1666464484
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1666464484
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1666464484
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1666464484
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1666464484
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1666464484
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1666464484
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1666464484
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1666464484
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1666464484
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1666464484
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1666464484
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1666464484
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1666464484
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1666464484
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1666464484
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1666464484
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1666464484
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1666464484
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1666464484
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1666464484
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1666464484
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1666464484
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1666464484
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1666464484
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1666464484
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1666464484
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1666464484
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1666464484
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1666464484
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1666464484
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1666464484
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1666464484
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1666464484
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1666464484
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1666464484
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1666464484
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1666464484
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1666464484
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1666464484
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1666464484
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1666464484
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1666464484
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1666464484
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1666464484
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1666464484
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1666464484
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1666464484
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1666464484
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1666464484
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1666464484
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1666464484
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1666464484
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1666464484
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1666464484
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1666464484
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1666464484
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_613
timestamp 1666464484
transform 1 0 57500 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_623
timestamp 1666464484
transform 1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_9
timestamp 1666464484
transform 1 0 1932 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1666464484
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1666464484
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1666464484
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1666464484
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1666464484
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1666464484
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1666464484
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1666464484
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1666464484
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1666464484
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1666464484
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1666464484
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1666464484
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1666464484
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1666464484
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1666464484
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1666464484
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1666464484
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1666464484
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1666464484
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1666464484
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1666464484
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1666464484
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1666464484
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1666464484
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1666464484
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1666464484
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1666464484
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1666464484
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1666464484
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1666464484
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1666464484
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1666464484
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1666464484
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1666464484
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1666464484
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1666464484
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1666464484
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1666464484
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1666464484
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1666464484
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1666464484
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1666464484
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1666464484
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1666464484
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1666464484
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1666464484
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1666464484
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1666464484
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1666464484
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1666464484
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1666464484
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1666464484
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1666464484
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1666464484
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1666464484
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1666464484
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1666464484
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1666464484
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1666464484
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1666464484
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_609
timestamp 1666464484
transform 1 0 57132 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_614
timestamp 1666464484
transform 1 0 57592 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_91_617
timestamp 1666464484
transform 1 0 57868 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_623
timestamp 1666464484
transform 1 0 58420 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_9
timestamp 1666464484
transform 1 0 1932 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1666464484
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1666464484
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1666464484
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1666464484
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1666464484
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1666464484
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1666464484
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1666464484
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1666464484
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1666464484
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1666464484
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1666464484
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1666464484
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1666464484
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1666464484
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1666464484
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1666464484
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1666464484
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1666464484
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1666464484
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1666464484
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1666464484
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1666464484
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1666464484
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1666464484
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1666464484
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1666464484
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1666464484
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1666464484
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1666464484
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_92_301
timestamp 1666464484
transform 1 0 28796 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_305
timestamp 1666464484
transform 1 0 29164 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1666464484
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1666464484
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1666464484
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1666464484
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1666464484
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1666464484
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1666464484
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1666464484
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1666464484
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1666464484
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1666464484
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1666464484
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1666464484
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1666464484
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1666464484
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1666464484
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1666464484
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1666464484
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1666464484
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1666464484
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1666464484
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1666464484
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1666464484
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1666464484
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1666464484
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1666464484
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1666464484
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1666464484
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1666464484
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1666464484
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1666464484
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1666464484
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_613
timestamp 1666464484
transform 1 0 57500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_616
timestamp 1666464484
transform 1 0 57776 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_623
timestamp 1666464484
transform 1 0 58420 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1666464484
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1666464484
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1666464484
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1666464484
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1666464484
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1666464484
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1666464484
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1666464484
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1666464484
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1666464484
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1666464484
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1666464484
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1666464484
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1666464484
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1666464484
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1666464484
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1666464484
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1666464484
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1666464484
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1666464484
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1666464484
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1666464484
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1666464484
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1666464484
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1666464484
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1666464484
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1666464484
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1666464484
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1666464484
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1666464484
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_293
timestamp 1666464484
transform 1 0 28060 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_303
timestamp 1666464484
transform 1 0 28980 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_316
timestamp 1666464484
transform 1 0 30176 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_328
timestamp 1666464484
transform 1 0 31280 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_337
timestamp 1666464484
transform 1 0 32108 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_344
timestamp 1666464484
transform 1 0 32752 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_356
timestamp 1666464484
transform 1 0 33856 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_368
timestamp 1666464484
transform 1 0 34960 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_380
timestamp 1666464484
transform 1 0 36064 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1666464484
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1666464484
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_417
timestamp 1666464484
transform 1 0 39468 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_421
timestamp 1666464484
transform 1 0 39836 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_427
timestamp 1666464484
transform 1 0 40388 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_439
timestamp 1666464484
transform 1 0 41492 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1666464484
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1666464484
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1666464484
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1666464484
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1666464484
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1666464484
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1666464484
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1666464484
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1666464484
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1666464484
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1666464484
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1666464484
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1666464484
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1666464484
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1666464484
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1666464484
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1666464484
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1666464484
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1666464484
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_9
timestamp 1666464484
transform 1 0 1932 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1666464484
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1666464484
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1666464484
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1666464484
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1666464484
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1666464484
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1666464484
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1666464484
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1666464484
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1666464484
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1666464484
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1666464484
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1666464484
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1666464484
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1666464484
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1666464484
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1666464484
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1666464484
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1666464484
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1666464484
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1666464484
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1666464484
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1666464484
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1666464484
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_245
timestamp 1666464484
transform 1 0 23644 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1666464484
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_253
timestamp 1666464484
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_263
timestamp 1666464484
transform 1 0 25300 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_275
timestamp 1666464484
transform 1 0 26404 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_287
timestamp 1666464484
transform 1 0 27508 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_299
timestamp 1666464484
transform 1 0 28612 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_303
timestamp 1666464484
transform 1 0 28980 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_306
timestamp 1666464484
transform 1 0 29256 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_309
timestamp 1666464484
transform 1 0 29532 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_324
timestamp 1666464484
transform 1 0 30912 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_328
timestamp 1666464484
transform 1 0 31280 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_335
timestamp 1666464484
transform 1 0 31924 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_352
timestamp 1666464484
transform 1 0 33488 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_358
timestamp 1666464484
transform 1 0 34040 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1666464484
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1666464484
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_389
timestamp 1666464484
transform 1 0 36892 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_395
timestamp 1666464484
transform 1 0 37444 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_398
timestamp 1666464484
transform 1 0 37720 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_408
timestamp 1666464484
transform 1 0 38640 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_418
timestamp 1666464484
transform 1 0 39560 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_421
timestamp 1666464484
transform 1 0 39836 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_430
timestamp 1666464484
transform 1 0 40664 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_436
timestamp 1666464484
transform 1 0 41216 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_448
timestamp 1666464484
transform 1 0 42320 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_460
timestamp 1666464484
transform 1 0 43424 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_472
timestamp 1666464484
transform 1 0 44528 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1666464484
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1666464484
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1666464484
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1666464484
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1666464484
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1666464484
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1666464484
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1666464484
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1666464484
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1666464484
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1666464484
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1666464484
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1666464484
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1666464484
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_613
timestamp 1666464484
transform 1 0 57500 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_616
timestamp 1666464484
transform 1 0 57776 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_623
timestamp 1666464484
transform 1 0 58420 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_9
timestamp 1666464484
transform 1 0 1932 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1666464484
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1666464484
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1666464484
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1666464484
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1666464484
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1666464484
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1666464484
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1666464484
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1666464484
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1666464484
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1666464484
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1666464484
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1666464484
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1666464484
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1666464484
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1666464484
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1666464484
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1666464484
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1666464484
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1666464484
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1666464484
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1666464484
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1666464484
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1666464484
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1666464484
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_249
timestamp 1666464484
transform 1 0 24012 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_259
timestamp 1666464484
transform 1 0 24932 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_269
timestamp 1666464484
transform 1 0 25852 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_275
timestamp 1666464484
transform 1 0 26404 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_278
timestamp 1666464484
transform 1 0 26680 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_281
timestamp 1666464484
transform 1 0 26956 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_291
timestamp 1666464484
transform 1 0 27876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_303
timestamp 1666464484
transform 1 0 28980 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_307
timestamp 1666464484
transform 1 0 29348 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1666464484
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_329
timestamp 1666464484
transform 1 0 31372 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_334
timestamp 1666464484
transform 1 0 31832 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_337
timestamp 1666464484
transform 1 0 32108 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_346
timestamp 1666464484
transform 1 0 32936 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_354
timestamp 1666464484
transform 1 0 33672 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_359
timestamp 1666464484
transform 1 0 34132 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_368
timestamp 1666464484
transform 1 0 34960 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_380
timestamp 1666464484
transform 1 0 36064 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_389
timestamp 1666464484
transform 1 0 36892 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_393
timestamp 1666464484
transform 1 0 37260 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_401
timestamp 1666464484
transform 1 0 37996 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_405
timestamp 1666464484
transform 1 0 38364 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_415
timestamp 1666464484
transform 1 0 39284 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_419
timestamp 1666464484
transform 1 0 39652 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_427
timestamp 1666464484
transform 1 0 40388 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_436
timestamp 1666464484
transform 1 0 41216 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_442
timestamp 1666464484
transform 1 0 41768 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1666464484
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1666464484
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1666464484
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1666464484
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1666464484
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1666464484
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1666464484
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1666464484
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1666464484
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1666464484
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1666464484
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1666464484
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1666464484
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1666464484
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1666464484
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1666464484
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1666464484
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1666464484
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_95_617
timestamp 1666464484
transform 1 0 57868 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_623
timestamp 1666464484
transform 1 0 58420 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1666464484
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1666464484
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1666464484
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1666464484
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1666464484
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1666464484
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1666464484
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1666464484
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1666464484
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1666464484
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1666464484
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1666464484
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1666464484
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1666464484
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1666464484
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1666464484
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1666464484
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1666464484
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1666464484
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1666464484
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1666464484
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1666464484
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_221
timestamp 1666464484
transform 1 0 21436 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_228
timestamp 1666464484
transform 1 0 22080 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_240
timestamp 1666464484
transform 1 0 23184 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1666464484
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_265
timestamp 1666464484
transform 1 0 25484 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_273
timestamp 1666464484
transform 1 0 26220 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_285
timestamp 1666464484
transform 1 0 27324 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_297
timestamp 1666464484
transform 1 0 28428 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_305
timestamp 1666464484
transform 1 0 29164 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1666464484
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1666464484
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_333
timestamp 1666464484
transform 1 0 31740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_336
timestamp 1666464484
transform 1 0 32016 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_347
timestamp 1666464484
transform 1 0 33028 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_359
timestamp 1666464484
transform 1 0 34132 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1666464484
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_365
timestamp 1666464484
transform 1 0 34684 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_375
timestamp 1666464484
transform 1 0 35604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_387
timestamp 1666464484
transform 1 0 36708 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_391
timestamp 1666464484
transform 1 0 37076 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_402
timestamp 1666464484
transform 1 0 38088 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_406
timestamp 1666464484
transform 1 0 38456 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_411
timestamp 1666464484
transform 1 0 38916 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_96_417
timestamp 1666464484
transform 1 0 39468 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_421
timestamp 1666464484
transform 1 0 39836 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_425
timestamp 1666464484
transform 1 0 40204 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_431
timestamp 1666464484
transform 1 0 40756 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_443
timestamp 1666464484
transform 1 0 41860 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_455
timestamp 1666464484
transform 1 0 42964 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_467
timestamp 1666464484
transform 1 0 44068 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1666464484
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1666464484
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1666464484
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1666464484
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1666464484
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1666464484
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1666464484
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1666464484
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1666464484
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1666464484
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1666464484
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1666464484
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1666464484
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1666464484
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1666464484
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_613
timestamp 1666464484
transform 1 0 57500 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_623
timestamp 1666464484
transform 1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_9
timestamp 1666464484
transform 1 0 1932 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1666464484
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1666464484
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1666464484
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1666464484
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1666464484
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1666464484
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1666464484
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1666464484
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1666464484
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1666464484
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1666464484
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1666464484
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1666464484
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1666464484
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1666464484
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1666464484
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1666464484
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1666464484
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1666464484
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1666464484
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1666464484
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1666464484
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1666464484
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_225
timestamp 1666464484
transform 1 0 21804 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_232
timestamp 1666464484
transform 1 0 22448 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_244
timestamp 1666464484
transform 1 0 23552 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_256
timestamp 1666464484
transform 1 0 24656 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_268
timestamp 1666464484
transform 1 0 25760 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1666464484
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1666464484
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_305
timestamp 1666464484
transform 1 0 29164 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_311
timestamp 1666464484
transform 1 0 29716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_323
timestamp 1666464484
transform 1 0 30820 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1666464484
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_337
timestamp 1666464484
transform 1 0 32108 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_341
timestamp 1666464484
transform 1 0 32476 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_353
timestamp 1666464484
transform 1 0 33580 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_365
timestamp 1666464484
transform 1 0 34684 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_377
timestamp 1666464484
transform 1 0 35788 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_389
timestamp 1666464484
transform 1 0 36892 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1666464484
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_407
timestamp 1666464484
transform 1 0 38548 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_415
timestamp 1666464484
transform 1 0 39284 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_420
timestamp 1666464484
transform 1 0 39744 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_432
timestamp 1666464484
transform 1 0 40848 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_444
timestamp 1666464484
transform 1 0 41952 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_449
timestamp 1666464484
transform 1 0 42412 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_459
timestamp 1666464484
transform 1 0 43332 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_471
timestamp 1666464484
transform 1 0 44436 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_483
timestamp 1666464484
transform 1 0 45540 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_495
timestamp 1666464484
transform 1 0 46644 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1666464484
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1666464484
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1666464484
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1666464484
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1666464484
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1666464484
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1666464484
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1666464484
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1666464484
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1666464484
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1666464484
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_609
timestamp 1666464484
transform 1 0 57132 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_614
timestamp 1666464484
transform 1 0 57592 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_97_617
timestamp 1666464484
transform 1 0 57868 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_623
timestamp 1666464484
transform 1 0 58420 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_9
timestamp 1666464484
transform 1 0 1932 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1666464484
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1666464484
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1666464484
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1666464484
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1666464484
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1666464484
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1666464484
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1666464484
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1666464484
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1666464484
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1666464484
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1666464484
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1666464484
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1666464484
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1666464484
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1666464484
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1666464484
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1666464484
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1666464484
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1666464484
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1666464484
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_209
timestamp 1666464484
transform 1 0 20332 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_217
timestamp 1666464484
transform 1 0 21068 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_223
timestamp 1666464484
transform 1 0 21620 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_235
timestamp 1666464484
transform 1 0 22724 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_238
timestamp 1666464484
transform 1 0 23000 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_250
timestamp 1666464484
transform 1 0 24104 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_253
timestamp 1666464484
transform 1 0 24380 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_261
timestamp 1666464484
transform 1 0 25116 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_273
timestamp 1666464484
transform 1 0 26220 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_283
timestamp 1666464484
transform 1 0 27140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_295
timestamp 1666464484
transform 1 0 28244 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_302
timestamp 1666464484
transform 1 0 28888 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_98_309
timestamp 1666464484
transform 1 0 29532 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_319
timestamp 1666464484
transform 1 0 30452 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_323
timestamp 1666464484
transform 1 0 30820 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_326
timestamp 1666464484
transform 1 0 31096 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_338
timestamp 1666464484
transform 1 0 32200 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_342
timestamp 1666464484
transform 1 0 32568 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_351
timestamp 1666464484
transform 1 0 33396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1666464484
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_365
timestamp 1666464484
transform 1 0 34684 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_373
timestamp 1666464484
transform 1 0 35420 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_383
timestamp 1666464484
transform 1 0 36340 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_395
timestamp 1666464484
transform 1 0 37444 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_403
timestamp 1666464484
transform 1 0 38180 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1666464484
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1666464484
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1666464484
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_433
timestamp 1666464484
transform 1 0 40940 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_443
timestamp 1666464484
transform 1 0 41860 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_455
timestamp 1666464484
transform 1 0 42964 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_98_466
timestamp 1666464484
transform 1 0 43976 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_474
timestamp 1666464484
transform 1 0 44712 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1666464484
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1666464484
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1666464484
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1666464484
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1666464484
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1666464484
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1666464484
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1666464484
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1666464484
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1666464484
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1666464484
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1666464484
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1666464484
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_601
timestamp 1666464484
transform 1 0 56396 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_607
timestamp 1666464484
transform 1 0 56948 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_610
timestamp 1666464484
transform 1 0 57224 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_616
timestamp 1666464484
transform 1 0 57776 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_623
timestamp 1666464484
transform 1 0 58420 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1666464484
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1666464484
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1666464484
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1666464484
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1666464484
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1666464484
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1666464484
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1666464484
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1666464484
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1666464484
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1666464484
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1666464484
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1666464484
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1666464484
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1666464484
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1666464484
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1666464484
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1666464484
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1666464484
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1666464484
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1666464484
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_222
timestamp 1666464484
transform 1 0 21528 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_225
timestamp 1666464484
transform 1 0 21804 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_232
timestamp 1666464484
transform 1 0 22448 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_252
timestamp 1666464484
transform 1 0 24288 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_258
timestamp 1666464484
transform 1 0 24840 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_265
timestamp 1666464484
transform 1 0 25484 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_99_277
timestamp 1666464484
transform 1 0 26588 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_281
timestamp 1666464484
transform 1 0 26956 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_291
timestamp 1666464484
transform 1 0 27876 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_299
timestamp 1666464484
transform 1 0 28612 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_308
timestamp 1666464484
transform 1 0 29440 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_322
timestamp 1666464484
transform 1 0 30728 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_334
timestamp 1666464484
transform 1 0 31832 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_337
timestamp 1666464484
transform 1 0 32108 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_341
timestamp 1666464484
transform 1 0 32476 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_350
timestamp 1666464484
transform 1 0 33304 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_370
timestamp 1666464484
transform 1 0 35144 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_382
timestamp 1666464484
transform 1 0 36248 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_390
timestamp 1666464484
transform 1 0 36984 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_393
timestamp 1666464484
transform 1 0 37260 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_402
timestamp 1666464484
transform 1 0 38088 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_413
timestamp 1666464484
transform 1 0 39100 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_425
timestamp 1666464484
transform 1 0 40204 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_437
timestamp 1666464484
transform 1 0 41308 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_445
timestamp 1666464484
transform 1 0 42044 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_449
timestamp 1666464484
transform 1 0 42412 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_465
timestamp 1666464484
transform 1 0 43884 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_477
timestamp 1666464484
transform 1 0 44988 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_489
timestamp 1666464484
transform 1 0 46092 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_501
timestamp 1666464484
transform 1 0 47196 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1666464484
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1666464484
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1666464484
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1666464484
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1666464484
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1666464484
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1666464484
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1666464484
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_599
timestamp 1666464484
transform 1 0 56212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_605
timestamp 1666464484
transform 1 0 56764 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_611
timestamp 1666464484
transform 1 0 57316 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1666464484
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_617
timestamp 1666464484
transform 1 0 57868 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1666464484
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_9
timestamp 1666464484
transform 1 0 1932 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_21
timestamp 1666464484
transform 1 0 3036 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_26
timestamp 1666464484
transform 1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_29
timestamp 1666464484
transform 1 0 3772 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_35
timestamp 1666464484
transform 1 0 4324 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_47
timestamp 1666464484
transform 1 0 5428 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_100_57
timestamp 1666464484
transform 1 0 6348 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_71
timestamp 1666464484
transform 1 0 7636 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_79
timestamp 1666464484
transform 1 0 8372 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_82
timestamp 1666464484
transform 1 0 8648 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_85
timestamp 1666464484
transform 1 0 8924 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_89
timestamp 1666464484
transform 1 0 9292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_101
timestamp 1666464484
transform 1 0 10396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_113
timestamp 1666464484
transform 1 0 11500 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_121
timestamp 1666464484
transform 1 0 12236 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_126
timestamp 1666464484
transform 1 0 12696 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_138
timestamp 1666464484
transform 1 0 13800 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_141
timestamp 1666464484
transform 1 0 14076 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_149
timestamp 1666464484
transform 1 0 14812 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_152
timestamp 1666464484
transform 1 0 15088 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_164
timestamp 1666464484
transform 1 0 16192 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_178
timestamp 1666464484
transform 1 0 17480 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_190
timestamp 1666464484
transform 1 0 18584 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_197
timestamp 1666464484
transform 1 0 19228 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_201
timestamp 1666464484
transform 1 0 19596 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_204
timestamp 1666464484
transform 1 0 19872 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_216
timestamp 1666464484
transform 1 0 20976 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_223
timestamp 1666464484
transform 1 0 21620 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_227
timestamp 1666464484
transform 1 0 21988 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_230
timestamp 1666464484
transform 1 0 22264 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_242
timestamp 1666464484
transform 1 0 23368 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_250
timestamp 1666464484
transform 1 0 24104 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_253
timestamp 1666464484
transform 1 0 24380 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_257
timestamp 1666464484
transform 1 0 24748 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_269
timestamp 1666464484
transform 1 0 25852 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_281
timestamp 1666464484
transform 1 0 26956 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_295
timestamp 1666464484
transform 1 0 28244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1666464484
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_309
timestamp 1666464484
transform 1 0 29532 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_317
timestamp 1666464484
transform 1 0 30268 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_329
timestamp 1666464484
transform 1 0 31372 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_339
timestamp 1666464484
transform 1 0 32292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_351
timestamp 1666464484
transform 1 0 33396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1666464484
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_365
timestamp 1666464484
transform 1 0 34684 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_371
timestamp 1666464484
transform 1 0 35236 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_374
timestamp 1666464484
transform 1 0 35512 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_382
timestamp 1666464484
transform 1 0 36248 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_386
timestamp 1666464484
transform 1 0 36616 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_398
timestamp 1666464484
transform 1 0 37720 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_403
timestamp 1666464484
transform 1 0 38180 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_414
timestamp 1666464484
transform 1 0 39192 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1666464484
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_433
timestamp 1666464484
transform 1 0 40940 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_438
timestamp 1666464484
transform 1 0 41400 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_450
timestamp 1666464484
transform 1 0 42504 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_100_466
timestamp 1666464484
transform 1 0 43976 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_474
timestamp 1666464484
transform 1 0 44712 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_477
timestamp 1666464484
transform 1 0 44988 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_481
timestamp 1666464484
transform 1 0 45356 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_493
timestamp 1666464484
transform 1 0 46460 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_507
timestamp 1666464484
transform 1 0 47748 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_519
timestamp 1666464484
transform 1 0 48852 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1666464484
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_533
timestamp 1666464484
transform 1 0 50140 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_537
timestamp 1666464484
transform 1 0 50508 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_549
timestamp 1666464484
transform 1 0 51612 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_555
timestamp 1666464484
transform 1 0 52164 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_567
timestamp 1666464484
transform 1 0 53268 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1666464484
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1666464484
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_589
timestamp 1666464484
transform 1 0 55292 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_593
timestamp 1666464484
transform 1 0 55660 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_596
timestamp 1666464484
transform 1 0 55936 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_602
timestamp 1666464484
transform 1 0 56488 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_609
timestamp 1666464484
transform 1 0 57132 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_616
timestamp 1666464484
transform 1 0 57776 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_623
timestamp 1666464484
transform 1 0 58420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_12
timestamp 1666464484
transform 1 0 2208 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_26
timestamp 1666464484
transform 1 0 3496 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_29
timestamp 1666464484
transform 1 0 3772 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_38
timestamp 1666464484
transform 1 0 4600 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1666464484
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_57
timestamp 1666464484
transform 1 0 6348 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_61
timestamp 1666464484
transform 1 0 6716 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_69
timestamp 1666464484
transform 1 0 7452 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_82
timestamp 1666464484
transform 1 0 8648 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_85
timestamp 1666464484
transform 1 0 8924 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_90
timestamp 1666464484
transform 1 0 9384 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_96
timestamp 1666464484
transform 1 0 9936 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_103
timestamp 1666464484
transform 1 0 10580 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_107
timestamp 1666464484
transform 1 0 10948 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_110
timestamp 1666464484
transform 1 0 11224 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_113
timestamp 1666464484
transform 1 0 11500 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_118
timestamp 1666464484
transform 1 0 11960 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_101_129
timestamp 1666464484
transform 1 0 12972 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_135
timestamp 1666464484
transform 1 0 13524 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_138
timestamp 1666464484
transform 1 0 13800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_141
timestamp 1666464484
transform 1 0 14076 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_146
timestamp 1666464484
transform 1 0 14536 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_155
timestamp 1666464484
transform 1 0 15364 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_163
timestamp 1666464484
transform 1 0 16100 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_166
timestamp 1666464484
transform 1 0 16376 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_169
timestamp 1666464484
transform 1 0 16652 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_174
timestamp 1666464484
transform 1 0 17112 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_181
timestamp 1666464484
transform 1 0 17756 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_187
timestamp 1666464484
transform 1 0 18308 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_194
timestamp 1666464484
transform 1 0 18952 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_197
timestamp 1666464484
transform 1 0 19228 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_203
timestamp 1666464484
transform 1 0 19780 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_207
timestamp 1666464484
transform 1 0 20148 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_213
timestamp 1666464484
transform 1 0 20700 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_220
timestamp 1666464484
transform 1 0 21344 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_225
timestamp 1666464484
transform 1 0 21804 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_229
timestamp 1666464484
transform 1 0 22172 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_233
timestamp 1666464484
transform 1 0 22540 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_239
timestamp 1666464484
transform 1 0 23092 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_246
timestamp 1666464484
transform 1 0 23736 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_101_253
timestamp 1666464484
transform 1 0 24380 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_259
timestamp 1666464484
transform 1 0 24932 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_265
timestamp 1666464484
transform 1 0 25484 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_272
timestamp 1666464484
transform 1 0 26128 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_278
timestamp 1666464484
transform 1 0 26680 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_281
timestamp 1666464484
transform 1 0 26956 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_286
timestamp 1666464484
transform 1 0 27416 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_294
timestamp 1666464484
transform 1 0 28152 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_298
timestamp 1666464484
transform 1 0 28520 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_306
timestamp 1666464484
transform 1 0 29256 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_309
timestamp 1666464484
transform 1 0 29532 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_314
timestamp 1666464484
transform 1 0 29992 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_320
timestamp 1666464484
transform 1 0 30544 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_324
timestamp 1666464484
transform 1 0 30912 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_330
timestamp 1666464484
transform 1 0 31464 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_337
timestamp 1666464484
transform 1 0 32108 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_342
timestamp 1666464484
transform 1 0 32568 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_346
timestamp 1666464484
transform 1 0 32936 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_350
timestamp 1666464484
transform 1 0 33304 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_356
timestamp 1666464484
transform 1 0 33856 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_362
timestamp 1666464484
transform 1 0 34408 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_365
timestamp 1666464484
transform 1 0 34684 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_370
timestamp 1666464484
transform 1 0 35144 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_377
timestamp 1666464484
transform 1 0 35788 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_385
timestamp 1666464484
transform 1 0 36524 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1666464484
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_393
timestamp 1666464484
transform 1 0 37260 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_402
timestamp 1666464484
transform 1 0 38088 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_408
timestamp 1666464484
transform 1 0 38640 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_415
timestamp 1666464484
transform 1 0 39284 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_419
timestamp 1666464484
transform 1 0 39652 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_421
timestamp 1666464484
transform 1 0 39836 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_428
timestamp 1666464484
transform 1 0 40480 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_434
timestamp 1666464484
transform 1 0 41032 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1666464484
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1666464484
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_449
timestamp 1666464484
transform 1 0 42412 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_454
timestamp 1666464484
transform 1 0 42872 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_460
timestamp 1666464484
transform 1 0 43424 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_467
timestamp 1666464484
transform 1 0 44068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1666464484
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_477
timestamp 1666464484
transform 1 0 44988 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_482
timestamp 1666464484
transform 1 0 45448 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_493
timestamp 1666464484
transform 1 0 46460 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_499
timestamp 1666464484
transform 1 0 47012 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1666464484
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_505
timestamp 1666464484
transform 1 0 47564 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_510
timestamp 1666464484
transform 1 0 48024 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_519
timestamp 1666464484
transform 1 0 48852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_525
timestamp 1666464484
transform 1 0 49404 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_531
timestamp 1666464484
transform 1 0 49956 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1666464484
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_538
timestamp 1666464484
transform 1 0 50600 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_545
timestamp 1666464484
transform 1 0 51244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_551
timestamp 1666464484
transform 1 0 51796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_558
timestamp 1666464484
transform 1 0 52440 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_561
timestamp 1666464484
transform 1 0 52716 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_567
timestamp 1666464484
transform 1 0 53268 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_571
timestamp 1666464484
transform 1 0 53636 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_577
timestamp 1666464484
transform 1 0 54188 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_584
timestamp 1666464484
transform 1 0 54832 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_589
timestamp 1666464484
transform 1 0 55292 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_593
timestamp 1666464484
transform 1 0 55660 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_597
timestamp 1666464484
transform 1 0 56028 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_603
timestamp 1666464484
transform 1 0 56580 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_610
timestamp 1666464484
transform 1 0 57224 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_101_617
timestamp 1666464484
transform 1 0 57868 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_623
timestamp 1666464484
transform 1 0 58420 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _208_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3036 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _209_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3220 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 1666464484
transform -1 0 6624 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1666464484
transform -1 0 7084 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 1666464484
transform 1 0 11776 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1666464484
transform -1 0 9016 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 1666464484
transform 1 0 8004 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1666464484
transform -1 0 7912 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1666464484
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1666464484
transform 1 0 15732 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1666464484
transform -1 0 19780 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1666464484
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1666464484
transform 1 0 19596 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _221_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19228 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1666464484
transform 1 0 18768 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1666464484
transform 1 0 17756 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1666464484
transform 1 0 19412 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1666464484
transform 1 0 18400 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _226_
timestamp 1666464484
transform 1 0 19596 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1666464484
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1666464484
transform -1 0 22356 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1666464484
transform 1 0 21988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1666464484
transform 1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1666464484
transform 1 0 18400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _232_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 38732 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _233_
timestamp 1666464484
transform 1 0 38088 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _234_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33488 0 1 53312
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _235_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 32752 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _236_
timestamp 1666464484
transform 1 0 29716 0 1 53312
box -38 -48 1234 592
use sky130_fd_sc_hd__or3b_4  _237_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29348 0 -1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _238_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30268 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _239_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _240_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32384 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _241_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 38548 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _242_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37444 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _243_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 40756 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _244_
timestamp 1666464484
transform 1 0 40020 0 1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _245_
timestamp 1666464484
transform 1 0 39744 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _246_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 41860 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _247_
timestamp 1666464484
transform -1 0 34960 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _248_
timestamp 1666464484
transform -1 0 33304 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _249_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31924 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _250_
timestamp 1666464484
transform -1 0 24288 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _251_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _252_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _253_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23368 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _254_
timestamp 1666464484
transform -1 0 41308 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _255_
timestamp 1666464484
transform 1 0 38456 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _256_
timestamp 1666464484
transform -1 0 33396 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _257_
timestamp 1666464484
transform -1 0 25484 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _258_
timestamp 1666464484
transform 1 0 25852 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _259_
timestamp 1666464484
transform 1 0 21068 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _260_
timestamp 1666464484
transform 1 0 27140 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _261_
timestamp 1666464484
transform -1 0 43332 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _262_
timestamp 1666464484
transform 1 0 36248 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _263_
timestamp 1666464484
transform -1 0 35604 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _264_
timestamp 1666464484
transform 1 0 25300 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1666464484
transform -1 0 24932 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _266_
timestamp 1666464484
transform 1 0 21620 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _267_
timestamp 1666464484
transform 1 0 24564 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _268_
timestamp 1666464484
transform -1 0 43976 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _269_
timestamp 1666464484
transform 1 0 38548 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _270_
timestamp 1666464484
transform -1 0 35144 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _271_
timestamp 1666464484
transform 1 0 25668 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _272_
timestamp 1666464484
transform 1 0 26588 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _273_
timestamp 1666464484
transform 1 0 21988 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _274_
timestamp 1666464484
transform 1 0 27140 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _275_
timestamp 1666464484
transform -1 0 43976 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _276_
timestamp 1666464484
transform 1 0 38456 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _277_
timestamp 1666464484
transform -1 0 36248 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _278_
timestamp 1666464484
transform -1 0 28888 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _279_
timestamp 1666464484
transform 1 0 28704 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _280_
timestamp 1666464484
transform 1 0 21160 0 1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _281_
timestamp 1666464484
transform 1 0 29716 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _282_
timestamp 1666464484
transform -1 0 43884 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _283_
timestamp 1666464484
transform 1 0 37444 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _284_
timestamp 1666464484
transform -1 0 36340 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _285_
timestamp 1666464484
transform -1 0 30268 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _286_
timestamp 1666464484
transform 1 0 29992 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _287_
timestamp 1666464484
transform 1 0 21160 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _288_
timestamp 1666464484
transform 1 0 31096 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _289_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 56948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _290_
timestamp 1666464484
transform 1 0 56120 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _291_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 56488 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1666464484
transform 1 0 58052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _293_
timestamp 1666464484
transform 1 0 55660 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1666464484
transform 1 0 56948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 57592 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1666464484
transform 1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _297_
timestamp 1666464484
transform -1 0 58420 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1666464484
transform 1 0 57316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _299_
timestamp 1666464484
transform -1 0 58420 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1666464484
transform 1 0 58052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _301_
timestamp 1666464484
transform -1 0 58420 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1666464484
transform 1 0 55476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _303_
timestamp 1666464484
transform -1 0 58420 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1666464484
transform 1 0 44068 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _305_
timestamp 1666464484
transform -1 0 58420 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _306_
timestamp 1666464484
transform -1 0 58328 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_2  _307_
timestamp 1666464484
transform -1 0 57868 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp 1666464484
transform 1 0 46276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _309_
timestamp 1666464484
transform -1 0 58144 0 1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1666464484
transform 1 0 57132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _311_
timestamp 1666464484
transform -1 0 57960 0 1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1666464484
transform 1 0 48300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _313_
timestamp 1666464484
transform -1 0 58144 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _314_
timestamp 1666464484
transform -1 0 53820 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _315_
timestamp 1666464484
transform -1 0 56304 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _316_
timestamp 1666464484
transform -1 0 55108 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _317_
timestamp 1666464484
transform -1 0 58236 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _318_
timestamp 1666464484
transform -1 0 52440 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_2  _319_
timestamp 1666464484
transform -1 0 58420 0 1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1666464484
transform 1 0 52900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _321_
timestamp 1666464484
transform -1 0 56028 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1666464484
transform 1 0 54372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _323_
timestamp 1666464484
transform -1 0 57500 0 -1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1666464484
transform 1 0 55476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _325_
timestamp 1666464484
transform -1 0 58236 0 1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1666464484
transform 1 0 56304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _327_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23000 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _328_
timestamp 1666464484
transform -1 0 18952 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1666464484
transform -1 0 3496 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1666464484
transform -1 0 4232 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1666464484
transform -1 0 8556 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1666464484
transform -1 0 9200 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1666464484
transform 1 0 9108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1666464484
transform -1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1666464484
transform -1 0 3404 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1666464484
transform -1 0 4416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1666464484
transform -1 0 6072 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1666464484
transform -1 0 6808 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1666464484
transform -1 0 5244 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1666464484
transform -1 0 5428 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1666464484
transform -1 0 6256 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1666464484
transform -1 0 7268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1666464484
transform 1 0 10212 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1666464484
transform -1 0 10212 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1666464484
transform 1 0 10672 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1666464484
transform -1 0 11132 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1666464484
transform 1 0 16928 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1666464484
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1666464484
transform 1 0 19596 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp 1666464484
transform 1 0 18952 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1666464484
transform 1 0 18952 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1666464484
transform 1 0 18124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1666464484
transform 1 0 18584 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1666464484
transform 1 0 17388 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1666464484
transform 1 0 18768 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1666464484
transform 1 0 17756 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1666464484
transform 1 0 20884 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1666464484
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1666464484
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _360_
timestamp 1666464484
transform 1 0 20792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _361_
timestamp 1666464484
transform 1 0 22172 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _362_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _363_
timestamp 1666464484
transform -1 0 20976 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1666464484
transform -1 0 2760 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _365_
timestamp 1666464484
transform -1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _366_
timestamp 1666464484
transform -1 0 2760 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp 1666464484
transform -1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1666464484
transform -1 0 2852 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _369_
timestamp 1666464484
transform -1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1666464484
transform -1 0 2760 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _371_
timestamp 1666464484
transform -1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1666464484
transform -1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1666464484
transform -1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1666464484
transform -1 0 2760 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1666464484
transform -1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1666464484
transform -1 0 2760 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1666464484
transform -1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1666464484
transform 1 0 11684 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1666464484
transform -1 0 10396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1666464484
transform 1 0 19688 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1666464484
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1666464484
transform -1 0 19688 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _383_
timestamp 1666464484
transform 1 0 19044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1666464484
transform 1 0 19228 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1666464484
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1666464484
transform 1 0 19688 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _387_
timestamp 1666464484
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1666464484
transform -1 0 18952 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _389_
timestamp 1666464484
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _391_
timestamp 1666464484
transform 1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1666464484
transform -1 0 22816 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _393_
timestamp 1666464484
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1666464484
transform 1 0 22172 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _395_
timestamp 1666464484
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _396_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23000 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  _397_
timestamp 1666464484
transform -1 0 18952 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1666464484
transform -1 0 2760 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1666464484
transform -1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1666464484
transform -1 0 2760 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _401_
timestamp 1666464484
transform -1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1666464484
transform -1 0 2760 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1666464484
transform -1 0 2576 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1666464484
transform -1 0 2484 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp 1666464484
transform -1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1666464484
transform -1 0 2760 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1666464484
transform -1 0 2576 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1666464484
transform -1 0 2760 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1666464484
transform -1 0 2576 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1666464484
transform 1 0 12696 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1666464484
transform -1 0 12512 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1666464484
transform -1 0 10488 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1666464484
transform -1 0 12972 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1666464484
transform 1 0 14260 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1666464484
transform 1 0 12880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _416_
timestamp 1666464484
transform 1 0 17020 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _417_
timestamp 1666464484
transform -1 0 16652 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp 1666464484
transform 1 0 18124 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _419_
timestamp 1666464484
transform 1 0 17296 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp 1666464484
transform 1 0 19412 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _421_
timestamp 1666464484
transform 1 0 18216 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp 1666464484
transform 1 0 18308 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _423_
timestamp 1666464484
transform 1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _424_
timestamp 1666464484
transform 1 0 19412 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _425_
timestamp 1666464484
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _426_
timestamp 1666464484
transform 1 0 20424 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _427_
timestamp 1666464484
transform 1 0 19688 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _428_
timestamp 1666464484
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 1666464484
transform 1 0 18124 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _430_
timestamp 1666464484
transform 1 0 22172 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  _431_
timestamp 1666464484
transform -1 0 20700 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _432_
timestamp 1666464484
transform -1 0 2760 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _433_
timestamp 1666464484
transform -1 0 3312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _434_
timestamp 1666464484
transform -1 0 2760 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1666464484
transform -1 0 2668 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1666464484
transform 1 0 11684 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1666464484
transform 1 0 11224 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _438_
timestamp 1666464484
transform -1 0 2944 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _439_
timestamp 1666464484
transform -1 0 3128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _440_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5980 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _441_
timestamp 1666464484
transform -1 0 12696 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _442_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8740 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _443_
timestamp 1666464484
transform -1 0 11040 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _444_
timestamp 1666464484
transform -1 0 8464 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _445_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8556 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _446_
timestamp 1666464484
transform -1 0 10120 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _447_
timestamp 1666464484
transform 1 0 10396 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _448_
timestamp 1666464484
transform -1 0 11868 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _449_
timestamp 1666464484
transform -1 0 7728 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _450_
timestamp 1666464484
transform -1 0 7636 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _451_
timestamp 1666464484
transform 1 0 16836 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _452_
timestamp 1666464484
transform -1 0 4968 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _453_
timestamp 1666464484
transform -1 0 17296 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _454_
timestamp 1666464484
transform -1 0 15180 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _455_
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _456_
timestamp 1666464484
transform -1 0 5980 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _457_
timestamp 1666464484
transform -1 0 5888 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _458_
timestamp 1666464484
transform -1 0 8648 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _459_
timestamp 1666464484
transform -1 0 6256 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _460_
timestamp 1666464484
transform -1 0 6072 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _461_
timestamp 1666464484
transform -1 0 10028 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _462_
timestamp 1666464484
transform -1 0 6072 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _463_
timestamp 1666464484
transform 1 0 10764 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _464_
timestamp 1666464484
transform -1 0 14444 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1666464484
transform -1 0 14168 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 1666464484
transform -1 0 15732 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _467_
timestamp 1666464484
transform -1 0 15640 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _468_
timestamp 1666464484
transform -1 0 16376 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 1666464484
transform -1 0 16560 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _470_
timestamp 1666464484
transform -1 0 9844 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _471_
timestamp 1666464484
transform -1 0 10396 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1666464484
transform 1 0 9108 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _473_
timestamp 1666464484
transform -1 0 6072 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _474_
timestamp 1666464484
transform 1 0 9292 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _475_
timestamp 1666464484
transform -1 0 5796 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1666464484
transform -1 0 5796 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1666464484
transform -1 0 7636 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _478_
timestamp 1666464484
transform -1 0 12972 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _479_
timestamp 1666464484
transform -1 0 14536 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _480_
timestamp 1666464484
transform 1 0 13156 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _481_
timestamp 1666464484
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 1666464484
transform -1 0 16100 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _483_
timestamp 1666464484
transform 1 0 9476 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1666464484
transform -1 0 16192 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _485_
timestamp 1666464484
transform -1 0 17664 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _486_
timestamp 1666464484
transform -1 0 16836 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _487_
timestamp 1666464484
transform -1 0 16008 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1666464484
transform 1 0 8648 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1666464484
transform -1 0 6900 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1666464484
transform 1 0 10856 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 1666464484
transform -1 0 7728 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 1666464484
transform -1 0 8648 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 1666464484
transform -1 0 13340 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _494_
timestamp 1666464484
transform 1 0 9292 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1666464484
transform -1 0 10120 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _496_
timestamp 1666464484
transform -1 0 15088 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _497_
timestamp 1666464484
transform -1 0 15456 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _498_
timestamp 1666464484
transform -1 0 6256 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _499_
timestamp 1666464484
transform -1 0 13800 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _500_
timestamp 1666464484
transform -1 0 17848 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _501_
timestamp 1666464484
transform -1 0 14168 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _502_
timestamp 1666464484
transform -1 0 17940 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _503_
timestamp 1666464484
transform 1 0 16652 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1666464484
transform -1 0 57868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_reg_wr_i dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11500 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_reg_wr_i
timestamp 1666464484
transform -1 0 9660 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_reg_wr_i
timestamp 1666464484
transform -1 0 9660 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_reg_wr_i
timestamp 1666464484
transform 1 0 12972 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_reg_wr_i
timestamp 1666464484
transform 1 0 12972 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_reg_wr_i
timestamp 1666464484
transform -1 0 9660 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_reg_wr_i
timestamp 1666464484
transform -1 0 9660 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_reg_wr_i
timestamp 1666464484
transform 1 0 12972 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_reg_wr_i
timestamp 1666464484
transform 1 0 12972 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout235
timestamp 1666464484
transform 1 0 6348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout236
timestamp 1666464484
transform -1 0 5888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout237
timestamp 1666464484
transform -1 0 12788 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout238
timestamp 1666464484
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout239
timestamp 1666464484
transform 1 0 5336 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout240 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout241
timestamp 1666464484
transform 1 0 14536 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout242
timestamp 1666464484
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout243
timestamp 1666464484
transform 1 0 5336 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform -1 0 56764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 2208 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1666464484
transform -1 0 3496 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1666464484
transform -1 0 4600 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1666464484
transform -1 0 6072 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1666464484
transform 1 0 6716 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1666464484
transform -1 0 8648 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1666464484
transform -1 0 9384 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1666464484
transform -1 0 10580 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform -1 0 11960 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform -1 0 12972 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1666464484
transform -1 0 14536 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform -1 0 15364 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1666464484
transform -1 0 17112 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1666464484
transform -1 0 17756 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1666464484
transform -1 0 18952 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1666464484
transform -1 0 20148 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1666464484
transform -1 0 21344 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1666464484
transform -1 0 22540 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1666464484
transform -1 0 23736 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1666464484
transform -1 0 24932 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1666464484
transform 1 0 25852 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1666464484
transform 1 0 27140 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1666464484
transform -1 0 28520 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1666464484
transform 1 0 29716 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1666464484
transform -1 0 30912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1666464484
transform -1 0 32568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1666464484
transform -1 0 33304 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1666464484
transform 1 0 34868 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1666464484
transform -1 0 35788 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1666464484
transform 1 0 36616 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1666464484
transform 1 0 37812 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1666464484
transform 1 0 39008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1666464484
transform 1 0 40204 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1666464484
transform 1 0 41400 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1666464484
transform 1 0 42596 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1666464484
transform 1 0 43792 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1666464484
transform 1 0 45172 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1666464484
transform 1 0 46184 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1666464484
transform 1 0 47748 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1666464484
transform 1 0 48576 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1666464484
transform 1 0 50324 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1666464484
transform 1 0 50968 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1666464484
transform 1 0 52164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1666464484
transform 1 0 53360 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1666464484
transform 1 0 54556 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1666464484
transform 1 0 55752 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1666464484
transform 1 0 56948 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1666464484
transform 1 0 58144 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input50
timestamp 1666464484
transform 1 0 24564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1666464484
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  input52 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  input53
timestamp 1666464484
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1666464484
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1666464484
transform -1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1666464484
transform 1 0 17848 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1666464484
transform -1 0 18952 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1666464484
transform 1 0 20056 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1666464484
transform 1 0 20608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1666464484
transform -1 0 22540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1666464484
transform 1 0 23184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1666464484
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1666464484
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1666464484
transform -1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1666464484
transform -1 0 11224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1666464484
transform -1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1666464484
transform 1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1666464484
transform -1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1666464484
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1666464484
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1666464484
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1666464484
transform 1 0 56488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1666464484
transform 1 0 55844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1666464484
transform 1 0 57316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1666464484
transform -1 0 57776 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1666464484
transform 1 0 58144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1666464484
transform 1 0 58144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1666464484
transform 1 0 58144 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1666464484
transform 1 0 57316 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1666464484
transform 1 0 58144 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1666464484
transform 1 0 58144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1666464484
transform 1 0 58144 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1666464484
transform 1 0 58144 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1666464484
transform 1 0 58144 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1666464484
transform 1 0 58144 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1666464484
transform 1 0 58144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1666464484
transform 1 0 58144 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1666464484
transform 1 0 58144 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1666464484
transform 1 0 58144 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1666464484
transform 1 0 58144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1666464484
transform 1 0 58144 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1666464484
transform 1 0 58144 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1666464484
transform -1 0 58420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1666464484
transform -1 0 58420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1666464484
transform -1 0 58420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1666464484
transform -1 0 58420 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1666464484
transform 1 0 58144 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1666464484
transform 1 0 58144 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1666464484
transform -1 0 58420 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1666464484
transform 1 0 58144 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1666464484
transform 1 0 58144 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1666464484
transform 1 0 58144 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1666464484
transform 1 0 58144 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1666464484
transform 1 0 58144 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1666464484
transform 1 0 58144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1666464484
transform 1 0 58144 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1666464484
transform 1 0 58144 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1666464484
transform 1 0 58144 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1666464484
transform 1 0 58144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1666464484
transform 1 0 58144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1666464484
transform 1 0 58144 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1666464484
transform 1 0 58144 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1666464484
transform 1 0 58144 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1666464484
transform 1 0 58144 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1666464484
transform 1 0 58144 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1666464484
transform 1 0 58144 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1666464484
transform 1 0 58144 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1666464484
transform 1 0 58144 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1666464484
transform 1 0 58144 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1666464484
transform 1 0 58144 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1666464484
transform 1 0 58144 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1666464484
transform 1 0 58144 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1666464484
transform 1 0 58144 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1666464484
transform 1 0 58144 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1666464484
transform 1 0 58144 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1666464484
transform 1 0 58144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1666464484
transform 1 0 58144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1666464484
transform 1 0 58144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1666464484
transform 1 0 58144 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1666464484
transform 1 0 58144 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1666464484
transform 1 0 58144 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1666464484
transform 1 0 58144 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1666464484
transform 1 0 58144 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1666464484
transform -1 0 57776 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1666464484
transform 1 0 58144 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1666464484
transform 1 0 58144 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1666464484
transform 1 0 58144 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input138
timestamp 1666464484
transform 1 0 58144 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1666464484
transform 1 0 58144 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1666464484
transform 1 0 58144 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1666464484
transform 1 0 58144 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1666464484
transform 1 0 58144 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1666464484
transform 1 0 56856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input144 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34868 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input145
timestamp 1666464484
transform 1 0 36064 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1666464484
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1666464484
transform 1 0 27784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1666464484
transform 1 0 28888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1666464484
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1666464484
transform 1 0 31096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1666464484
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1666464484
transform 1 0 33304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1666464484
transform -1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1666464484
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1666464484
transform -1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1666464484
transform -1 0 2668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1666464484
transform -1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1666464484
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1666464484
transform -1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1666464484
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1666464484
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1666464484
transform -1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1666464484
transform -1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1666464484
transform -1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1666464484
transform -1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1666464484
transform -1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1666464484
transform -1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1666464484
transform -1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1666464484
transform -1 0 2668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1666464484
transform -1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1666464484
transform -1 0 1932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1666464484
transform -1 0 1932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1666464484
transform -1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1666464484
transform -1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1666464484
transform -1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1666464484
transform -1 0 1932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1666464484
transform -1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1666464484
transform -1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1666464484
transform -1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1666464484
transform -1 0 1932 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1666464484
transform -1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1666464484
transform -1 0 1932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1666464484
transform -1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1666464484
transform -1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1666464484
transform -1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1666464484
transform -1 0 1932 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1666464484
transform -1 0 1932 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1666464484
transform -1 0 1932 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1666464484
transform -1 0 1932 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1666464484
transform -1 0 1932 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1666464484
transform -1 0 1932 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1666464484
transform -1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1666464484
transform -1 0 1932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1666464484
transform -1 0 1932 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1666464484
transform -1 0 1932 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1666464484
transform -1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1666464484
transform -1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1666464484
transform -1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1666464484
transform -1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1666464484
transform -1 0 1932 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1666464484
transform -1 0 1932 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1666464484
transform -1 0 1932 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1666464484
transform -1 0 1932 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1666464484
transform -1 0 1932 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1666464484
transform -1 0 1932 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1666464484
transform -1 0 1932 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1666464484
transform -1 0 1932 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1666464484
transform -1 0 1932 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1666464484
transform -1 0 1932 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1666464484
transform -1 0 1932 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1666464484
transform -1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1666464484
transform -1 0 1932 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1666464484
transform -1 0 1932 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1666464484
transform -1 0 1932 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1666464484
transform -1 0 1932 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1666464484
transform -1 0 1932 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1666464484
transform -1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1666464484
transform -1 0 38548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1666464484
transform 1 0 38916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1666464484
transform -1 0 40388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1666464484
transform -1 0 41400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1666464484
transform -1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1666464484
transform -1 0 43700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1666464484
transform -1 0 54648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1666464484
transform -1 0 55844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1666464484
transform -1 0 44712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1666464484
transform -1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1666464484
transform -1 0 46920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1666464484
transform -1 0 48116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1666464484
transform -1 0 49128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1666464484
transform -1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1666464484
transform -1 0 51428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1666464484
transform -1 0 52440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1666464484
transform -1 0 53544 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 56414 0 56470 800 0 FreeSans 224 90 0 0 loopback_i
port 0 nsew signal input
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 loopback_o
port 1 nsew signal tristate
flabel metal2 s 1858 59200 1914 60000 0 FreeSans 224 90 0 0 mux0_i[0]
port 2 nsew signal input
flabel metal2 s 3054 59200 3110 60000 0 FreeSans 224 90 0 0 mux0_i[1]
port 3 nsew signal input
flabel metal2 s 4250 59200 4306 60000 0 FreeSans 224 90 0 0 mux0_i[2]
port 4 nsew signal input
flabel metal2 s 5446 59200 5502 60000 0 FreeSans 224 90 0 0 mux0_i[3]
port 5 nsew signal input
flabel metal2 s 6642 59200 6698 60000 0 FreeSans 224 90 0 0 mux0_i[4]
port 6 nsew signal input
flabel metal2 s 7838 59200 7894 60000 0 FreeSans 224 90 0 0 mux0_i[5]
port 7 nsew signal input
flabel metal2 s 9034 59200 9090 60000 0 FreeSans 224 90 0 0 mux1_i[0]
port 8 nsew signal input
flabel metal2 s 10230 59200 10286 60000 0 FreeSans 224 90 0 0 mux1_i[1]
port 9 nsew signal input
flabel metal2 s 11426 59200 11482 60000 0 FreeSans 224 90 0 0 mux1_i[2]
port 10 nsew signal input
flabel metal2 s 12622 59200 12678 60000 0 FreeSans 224 90 0 0 mux1_i[3]
port 11 nsew signal input
flabel metal2 s 13818 59200 13874 60000 0 FreeSans 224 90 0 0 mux1_i[4]
port 12 nsew signal input
flabel metal2 s 15014 59200 15070 60000 0 FreeSans 224 90 0 0 mux1_i[5]
port 13 nsew signal input
flabel metal2 s 16210 59200 16266 60000 0 FreeSans 224 90 0 0 mux2_i[0]
port 14 nsew signal input
flabel metal2 s 17406 59200 17462 60000 0 FreeSans 224 90 0 0 mux2_i[1]
port 15 nsew signal input
flabel metal2 s 18602 59200 18658 60000 0 FreeSans 224 90 0 0 mux2_i[2]
port 16 nsew signal input
flabel metal2 s 19798 59200 19854 60000 0 FreeSans 224 90 0 0 mux2_i[3]
port 17 nsew signal input
flabel metal2 s 20994 59200 21050 60000 0 FreeSans 224 90 0 0 mux2_i[4]
port 18 nsew signal input
flabel metal2 s 22190 59200 22246 60000 0 FreeSans 224 90 0 0 mux2_i[5]
port 19 nsew signal input
flabel metal2 s 23386 59200 23442 60000 0 FreeSans 224 90 0 0 mux3_i[0]
port 20 nsew signal input
flabel metal2 s 24582 59200 24638 60000 0 FreeSans 224 90 0 0 mux3_i[1]
port 21 nsew signal input
flabel metal2 s 25778 59200 25834 60000 0 FreeSans 224 90 0 0 mux3_i[2]
port 22 nsew signal input
flabel metal2 s 26974 59200 27030 60000 0 FreeSans 224 90 0 0 mux3_i[3]
port 23 nsew signal input
flabel metal2 s 28170 59200 28226 60000 0 FreeSans 224 90 0 0 mux3_i[4]
port 24 nsew signal input
flabel metal2 s 29366 59200 29422 60000 0 FreeSans 224 90 0 0 mux3_i[5]
port 25 nsew signal input
flabel metal2 s 30562 59200 30618 60000 0 FreeSans 224 90 0 0 mux4_i[0]
port 26 nsew signal input
flabel metal2 s 31758 59200 31814 60000 0 FreeSans 224 90 0 0 mux4_i[1]
port 27 nsew signal input
flabel metal2 s 32954 59200 33010 60000 0 FreeSans 224 90 0 0 mux4_i[2]
port 28 nsew signal input
flabel metal2 s 34150 59200 34206 60000 0 FreeSans 224 90 0 0 mux4_i[3]
port 29 nsew signal input
flabel metal2 s 35346 59200 35402 60000 0 FreeSans 224 90 0 0 mux4_i[4]
port 30 nsew signal input
flabel metal2 s 36542 59200 36598 60000 0 FreeSans 224 90 0 0 mux4_i[5]
port 31 nsew signal input
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 mux5_i[0]
port 32 nsew signal input
flabel metal2 s 38934 59200 38990 60000 0 FreeSans 224 90 0 0 mux5_i[1]
port 33 nsew signal input
flabel metal2 s 40130 59200 40186 60000 0 FreeSans 224 90 0 0 mux5_i[2]
port 34 nsew signal input
flabel metal2 s 41326 59200 41382 60000 0 FreeSans 224 90 0 0 mux5_i[3]
port 35 nsew signal input
flabel metal2 s 42522 59200 42578 60000 0 FreeSans 224 90 0 0 mux5_i[4]
port 36 nsew signal input
flabel metal2 s 43718 59200 43774 60000 0 FreeSans 224 90 0 0 mux5_i[5]
port 37 nsew signal input
flabel metal2 s 44914 59200 44970 60000 0 FreeSans 224 90 0 0 mux6_i[0]
port 38 nsew signal input
flabel metal2 s 46110 59200 46166 60000 0 FreeSans 224 90 0 0 mux6_i[1]
port 39 nsew signal input
flabel metal2 s 47306 59200 47362 60000 0 FreeSans 224 90 0 0 mux6_i[2]
port 40 nsew signal input
flabel metal2 s 48502 59200 48558 60000 0 FreeSans 224 90 0 0 mux6_i[3]
port 41 nsew signal input
flabel metal2 s 49698 59200 49754 60000 0 FreeSans 224 90 0 0 mux6_i[4]
port 42 nsew signal input
flabel metal2 s 50894 59200 50950 60000 0 FreeSans 224 90 0 0 mux6_i[5]
port 43 nsew signal input
flabel metal2 s 52090 59200 52146 60000 0 FreeSans 224 90 0 0 mux7_i[0]
port 44 nsew signal input
flabel metal2 s 53286 59200 53342 60000 0 FreeSans 224 90 0 0 mux7_i[1]
port 45 nsew signal input
flabel metal2 s 54482 59200 54538 60000 0 FreeSans 224 90 0 0 mux7_i[2]
port 46 nsew signal input
flabel metal2 s 55678 59200 55734 60000 0 FreeSans 224 90 0 0 mux7_i[3]
port 47 nsew signal input
flabel metal2 s 56874 59200 56930 60000 0 FreeSans 224 90 0 0 mux7_i[4]
port 48 nsew signal input
flabel metal2 s 58070 59200 58126 60000 0 FreeSans 224 90 0 0 mux7_i[5]
port 49 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 mux_adr_i[0]
port 50 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 mux_adr_i[1]
port 51 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 mux_adr_i[2]
port 52 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 mux_o[0]
port 53 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 mux_o[1]
port 54 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 mux_o[2]
port 55 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 mux_o[3]
port 56 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 mux_o[4]
port 57 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 mux_o[5]
port 58 nsew signal tristate
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 reg0_o[0]
port 59 nsew signal tristate
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 reg0_o[10]
port 60 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 reg0_o[11]
port 61 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 reg0_o[12]
port 62 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 reg0_o[13]
port 63 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 reg0_o[14]
port 64 nsew signal tristate
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 reg0_o[15]
port 65 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 reg0_o[1]
port 66 nsew signal tristate
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 reg0_o[2]
port 67 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 reg0_o[3]
port 68 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 reg0_o[4]
port 69 nsew signal tristate
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 reg0_o[5]
port 70 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 reg0_o[6]
port 71 nsew signal tristate
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 reg0_o[7]
port 72 nsew signal tristate
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 reg0_o[8]
port 73 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 reg0_o[9]
port 74 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 reg1_o[0]
port 75 nsew signal tristate
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 reg1_o[10]
port 76 nsew signal tristate
flabel metal3 s 0 26256 800 26376 0 FreeSans 480 0 0 0 reg1_o[11]
port 77 nsew signal tristate
flabel metal3 s 0 27072 800 27192 0 FreeSans 480 0 0 0 reg1_o[12]
port 78 nsew signal tristate
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 reg1_o[13]
port 79 nsew signal tristate
flabel metal3 s 0 28704 800 28824 0 FreeSans 480 0 0 0 reg1_o[14]
port 80 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 reg1_o[15]
port 81 nsew signal tristate
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 reg1_o[1]
port 82 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 reg1_o[2]
port 83 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 reg1_o[3]
port 84 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 reg1_o[4]
port 85 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 reg1_o[5]
port 86 nsew signal tristate
flabel metal3 s 0 22176 800 22296 0 FreeSans 480 0 0 0 reg1_o[6]
port 87 nsew signal tristate
flabel metal3 s 0 22992 800 23112 0 FreeSans 480 0 0 0 reg1_o[7]
port 88 nsew signal tristate
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 reg1_o[8]
port 89 nsew signal tristate
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 reg1_o[9]
port 90 nsew signal tristate
flabel metal3 s 0 30336 800 30456 0 FreeSans 480 0 0 0 reg2_o[0]
port 91 nsew signal tristate
flabel metal3 s 0 38496 800 38616 0 FreeSans 480 0 0 0 reg2_o[10]
port 92 nsew signal tristate
flabel metal3 s 0 39312 800 39432 0 FreeSans 480 0 0 0 reg2_o[11]
port 93 nsew signal tristate
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 reg2_o[12]
port 94 nsew signal tristate
flabel metal3 s 0 40944 800 41064 0 FreeSans 480 0 0 0 reg2_o[13]
port 95 nsew signal tristate
flabel metal3 s 0 41760 800 41880 0 FreeSans 480 0 0 0 reg2_o[14]
port 96 nsew signal tristate
flabel metal3 s 0 42576 800 42696 0 FreeSans 480 0 0 0 reg2_o[15]
port 97 nsew signal tristate
flabel metal3 s 0 31152 800 31272 0 FreeSans 480 0 0 0 reg2_o[1]
port 98 nsew signal tristate
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 reg2_o[2]
port 99 nsew signal tristate
flabel metal3 s 0 32784 800 32904 0 FreeSans 480 0 0 0 reg2_o[3]
port 100 nsew signal tristate
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 reg2_o[4]
port 101 nsew signal tristate
flabel metal3 s 0 34416 800 34536 0 FreeSans 480 0 0 0 reg2_o[5]
port 102 nsew signal tristate
flabel metal3 s 0 35232 800 35352 0 FreeSans 480 0 0 0 reg2_o[6]
port 103 nsew signal tristate
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 reg2_o[7]
port 104 nsew signal tristate
flabel metal3 s 0 36864 800 36984 0 FreeSans 480 0 0 0 reg2_o[8]
port 105 nsew signal tristate
flabel metal3 s 0 37680 800 37800 0 FreeSans 480 0 0 0 reg2_o[9]
port 106 nsew signal tristate
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 reg3_o[0]
port 107 nsew signal tristate
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 reg3_o[10]
port 108 nsew signal tristate
flabel metal3 s 0 52368 800 52488 0 FreeSans 480 0 0 0 reg3_o[11]
port 109 nsew signal tristate
flabel metal3 s 0 53184 800 53304 0 FreeSans 480 0 0 0 reg3_o[12]
port 110 nsew signal tristate
flabel metal3 s 0 54000 800 54120 0 FreeSans 480 0 0 0 reg3_o[13]
port 111 nsew signal tristate
flabel metal3 s 0 54816 800 54936 0 FreeSans 480 0 0 0 reg3_o[14]
port 112 nsew signal tristate
flabel metal3 s 0 55632 800 55752 0 FreeSans 480 0 0 0 reg3_o[15]
port 113 nsew signal tristate
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 reg3_o[1]
port 114 nsew signal tristate
flabel metal3 s 0 45024 800 45144 0 FreeSans 480 0 0 0 reg3_o[2]
port 115 nsew signal tristate
flabel metal3 s 0 45840 800 45960 0 FreeSans 480 0 0 0 reg3_o[3]
port 116 nsew signal tristate
flabel metal3 s 0 46656 800 46776 0 FreeSans 480 0 0 0 reg3_o[4]
port 117 nsew signal tristate
flabel metal3 s 0 47472 800 47592 0 FreeSans 480 0 0 0 reg3_o[5]
port 118 nsew signal tristate
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 reg3_o[6]
port 119 nsew signal tristate
flabel metal3 s 0 49104 800 49224 0 FreeSans 480 0 0 0 reg3_o[7]
port 120 nsew signal tristate
flabel metal3 s 0 49920 800 50040 0 FreeSans 480 0 0 0 reg3_o[8]
port 121 nsew signal tristate
flabel metal3 s 0 50736 800 50856 0 FreeSans 480 0 0 0 reg3_o[9]
port 122 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 reg_adr_i[0]
port 123 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 reg_adr_i[1]
port 124 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 reg_dat_i[0]
port 125 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 reg_dat_i[10]
port 126 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 reg_dat_i[11]
port 127 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 reg_dat_i[12]
port 128 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 reg_dat_i[13]
port 129 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 reg_dat_i[14]
port 130 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 reg_dat_i[15]
port 131 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 reg_dat_i[1]
port 132 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 reg_dat_i[2]
port 133 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 reg_dat_i[3]
port 134 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 reg_dat_i[4]
port 135 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 reg_dat_i[5]
port 136 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 reg_dat_i[6]
port 137 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 reg_dat_i[7]
port 138 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 reg_dat_i[8]
port 139 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 reg_dat_i[9]
port 140 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 reg_wr_i
port 141 nsew signal input
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 rst_n_i
port 142 nsew signal input
flabel metal3 s 59200 960 60000 1080 0 FreeSans 480 0 0 0 temp0_dac_i[0]
port 143 nsew signal input
flabel metal3 s 59200 1776 60000 1896 0 FreeSans 480 0 0 0 temp0_dac_i[1]
port 144 nsew signal input
flabel metal3 s 59200 2592 60000 2712 0 FreeSans 480 0 0 0 temp0_dac_i[2]
port 145 nsew signal input
flabel metal3 s 59200 3408 60000 3528 0 FreeSans 480 0 0 0 temp0_dac_i[3]
port 146 nsew signal input
flabel metal3 s 59200 4224 60000 4344 0 FreeSans 480 0 0 0 temp0_dac_i[4]
port 147 nsew signal input
flabel metal3 s 59200 5040 60000 5160 0 FreeSans 480 0 0 0 temp0_dac_i[5]
port 148 nsew signal input
flabel metal3 s 59200 20544 60000 20664 0 FreeSans 480 0 0 0 temp0_ticks_i[0]
port 149 nsew signal input
flabel metal3 s 59200 28704 60000 28824 0 FreeSans 480 0 0 0 temp0_ticks_i[10]
port 150 nsew signal input
flabel metal3 s 59200 29520 60000 29640 0 FreeSans 480 0 0 0 temp0_ticks_i[11]
port 151 nsew signal input
flabel metal3 s 59200 21360 60000 21480 0 FreeSans 480 0 0 0 temp0_ticks_i[1]
port 152 nsew signal input
flabel metal3 s 59200 22176 60000 22296 0 FreeSans 480 0 0 0 temp0_ticks_i[2]
port 153 nsew signal input
flabel metal3 s 59200 22992 60000 23112 0 FreeSans 480 0 0 0 temp0_ticks_i[3]
port 154 nsew signal input
flabel metal3 s 59200 23808 60000 23928 0 FreeSans 480 0 0 0 temp0_ticks_i[4]
port 155 nsew signal input
flabel metal3 s 59200 24624 60000 24744 0 FreeSans 480 0 0 0 temp0_ticks_i[5]
port 156 nsew signal input
flabel metal3 s 59200 25440 60000 25560 0 FreeSans 480 0 0 0 temp0_ticks_i[6]
port 157 nsew signal input
flabel metal3 s 59200 26256 60000 26376 0 FreeSans 480 0 0 0 temp0_ticks_i[7]
port 158 nsew signal input
flabel metal3 s 59200 27072 60000 27192 0 FreeSans 480 0 0 0 temp0_ticks_i[8]
port 159 nsew signal input
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 temp0_ticks_i[9]
port 160 nsew signal input
flabel metal3 s 59200 5856 60000 5976 0 FreeSans 480 0 0 0 temp1_dac_i[0]
port 161 nsew signal input
flabel metal3 s 59200 6672 60000 6792 0 FreeSans 480 0 0 0 temp1_dac_i[1]
port 162 nsew signal input
flabel metal3 s 59200 7488 60000 7608 0 FreeSans 480 0 0 0 temp1_dac_i[2]
port 163 nsew signal input
flabel metal3 s 59200 8304 60000 8424 0 FreeSans 480 0 0 0 temp1_dac_i[3]
port 164 nsew signal input
flabel metal3 s 59200 9120 60000 9240 0 FreeSans 480 0 0 0 temp1_dac_i[4]
port 165 nsew signal input
flabel metal3 s 59200 9936 60000 10056 0 FreeSans 480 0 0 0 temp1_dac_i[5]
port 166 nsew signal input
flabel metal3 s 59200 30336 60000 30456 0 FreeSans 480 0 0 0 temp1_ticks_i[0]
port 167 nsew signal input
flabel metal3 s 59200 38496 60000 38616 0 FreeSans 480 0 0 0 temp1_ticks_i[10]
port 168 nsew signal input
flabel metal3 s 59200 39312 60000 39432 0 FreeSans 480 0 0 0 temp1_ticks_i[11]
port 169 nsew signal input
flabel metal3 s 59200 31152 60000 31272 0 FreeSans 480 0 0 0 temp1_ticks_i[1]
port 170 nsew signal input
flabel metal3 s 59200 31968 60000 32088 0 FreeSans 480 0 0 0 temp1_ticks_i[2]
port 171 nsew signal input
flabel metal3 s 59200 32784 60000 32904 0 FreeSans 480 0 0 0 temp1_ticks_i[3]
port 172 nsew signal input
flabel metal3 s 59200 33600 60000 33720 0 FreeSans 480 0 0 0 temp1_ticks_i[4]
port 173 nsew signal input
flabel metal3 s 59200 34416 60000 34536 0 FreeSans 480 0 0 0 temp1_ticks_i[5]
port 174 nsew signal input
flabel metal3 s 59200 35232 60000 35352 0 FreeSans 480 0 0 0 temp1_ticks_i[6]
port 175 nsew signal input
flabel metal3 s 59200 36048 60000 36168 0 FreeSans 480 0 0 0 temp1_ticks_i[7]
port 176 nsew signal input
flabel metal3 s 59200 36864 60000 36984 0 FreeSans 480 0 0 0 temp1_ticks_i[8]
port 177 nsew signal input
flabel metal3 s 59200 37680 60000 37800 0 FreeSans 480 0 0 0 temp1_ticks_i[9]
port 178 nsew signal input
flabel metal3 s 59200 10752 60000 10872 0 FreeSans 480 0 0 0 temp2_dac_i[0]
port 179 nsew signal input
flabel metal3 s 59200 11568 60000 11688 0 FreeSans 480 0 0 0 temp2_dac_i[1]
port 180 nsew signal input
flabel metal3 s 59200 12384 60000 12504 0 FreeSans 480 0 0 0 temp2_dac_i[2]
port 181 nsew signal input
flabel metal3 s 59200 13200 60000 13320 0 FreeSans 480 0 0 0 temp2_dac_i[3]
port 182 nsew signal input
flabel metal3 s 59200 14016 60000 14136 0 FreeSans 480 0 0 0 temp2_dac_i[4]
port 183 nsew signal input
flabel metal3 s 59200 14832 60000 14952 0 FreeSans 480 0 0 0 temp2_dac_i[5]
port 184 nsew signal input
flabel metal3 s 59200 40128 60000 40248 0 FreeSans 480 0 0 0 temp2_ticks_i[0]
port 185 nsew signal input
flabel metal3 s 59200 48288 60000 48408 0 FreeSans 480 0 0 0 temp2_ticks_i[10]
port 186 nsew signal input
flabel metal3 s 59200 49104 60000 49224 0 FreeSans 480 0 0 0 temp2_ticks_i[11]
port 187 nsew signal input
flabel metal3 s 59200 40944 60000 41064 0 FreeSans 480 0 0 0 temp2_ticks_i[1]
port 188 nsew signal input
flabel metal3 s 59200 41760 60000 41880 0 FreeSans 480 0 0 0 temp2_ticks_i[2]
port 189 nsew signal input
flabel metal3 s 59200 42576 60000 42696 0 FreeSans 480 0 0 0 temp2_ticks_i[3]
port 190 nsew signal input
flabel metal3 s 59200 43392 60000 43512 0 FreeSans 480 0 0 0 temp2_ticks_i[4]
port 191 nsew signal input
flabel metal3 s 59200 44208 60000 44328 0 FreeSans 480 0 0 0 temp2_ticks_i[5]
port 192 nsew signal input
flabel metal3 s 59200 45024 60000 45144 0 FreeSans 480 0 0 0 temp2_ticks_i[6]
port 193 nsew signal input
flabel metal3 s 59200 45840 60000 45960 0 FreeSans 480 0 0 0 temp2_ticks_i[7]
port 194 nsew signal input
flabel metal3 s 59200 46656 60000 46776 0 FreeSans 480 0 0 0 temp2_ticks_i[8]
port 195 nsew signal input
flabel metal3 s 59200 47472 60000 47592 0 FreeSans 480 0 0 0 temp2_ticks_i[9]
port 196 nsew signal input
flabel metal3 s 59200 15648 60000 15768 0 FreeSans 480 0 0 0 temp3_dac_i[0]
port 197 nsew signal input
flabel metal3 s 59200 16464 60000 16584 0 FreeSans 480 0 0 0 temp3_dac_i[1]
port 198 nsew signal input
flabel metal3 s 59200 17280 60000 17400 0 FreeSans 480 0 0 0 temp3_dac_i[2]
port 199 nsew signal input
flabel metal3 s 59200 18096 60000 18216 0 FreeSans 480 0 0 0 temp3_dac_i[3]
port 200 nsew signal input
flabel metal3 s 59200 18912 60000 19032 0 FreeSans 480 0 0 0 temp3_dac_i[4]
port 201 nsew signal input
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 temp3_dac_i[5]
port 202 nsew signal input
flabel metal3 s 59200 49920 60000 50040 0 FreeSans 480 0 0 0 temp3_ticks_i[0]
port 203 nsew signal input
flabel metal3 s 59200 58080 60000 58200 0 FreeSans 480 0 0 0 temp3_ticks_i[10]
port 204 nsew signal input
flabel metal3 s 59200 58896 60000 59016 0 FreeSans 480 0 0 0 temp3_ticks_i[11]
port 205 nsew signal input
flabel metal3 s 59200 50736 60000 50856 0 FreeSans 480 0 0 0 temp3_ticks_i[1]
port 206 nsew signal input
flabel metal3 s 59200 51552 60000 51672 0 FreeSans 480 0 0 0 temp3_ticks_i[2]
port 207 nsew signal input
flabel metal3 s 59200 52368 60000 52488 0 FreeSans 480 0 0 0 temp3_ticks_i[3]
port 208 nsew signal input
flabel metal3 s 59200 53184 60000 53304 0 FreeSans 480 0 0 0 temp3_ticks_i[4]
port 209 nsew signal input
flabel metal3 s 59200 54000 60000 54120 0 FreeSans 480 0 0 0 temp3_ticks_i[5]
port 210 nsew signal input
flabel metal3 s 59200 54816 60000 54936 0 FreeSans 480 0 0 0 temp3_ticks_i[6]
port 211 nsew signal input
flabel metal3 s 59200 55632 60000 55752 0 FreeSans 480 0 0 0 temp3_ticks_i[7]
port 212 nsew signal input
flabel metal3 s 59200 56448 60000 56568 0 FreeSans 480 0 0 0 temp3_ticks_i[8]
port 213 nsew signal input
flabel metal3 s 59200 57264 60000 57384 0 FreeSans 480 0 0 0 temp3_ticks_i[9]
port 214 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 temp_dac_o[0]
port 215 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 temp_dac_o[1]
port 216 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 temp_dac_o[2]
port 217 nsew signal tristate
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 temp_dac_o[3]
port 218 nsew signal tristate
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 temp_dac_o[4]
port 219 nsew signal tristate
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 temp_dac_o[5]
port 220 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 temp_sel_i[0]
port 221 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 temp_sel_i[1]
port 222 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 temp_ticks_o[0]
port 223 nsew signal tristate
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 temp_ticks_o[10]
port 224 nsew signal tristate
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 temp_ticks_o[11]
port 225 nsew signal tristate
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 temp_ticks_o[1]
port 226 nsew signal tristate
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 temp_ticks_o[2]
port 227 nsew signal tristate
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 temp_ticks_o[3]
port 228 nsew signal tristate
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 temp_ticks_o[4]
port 229 nsew signal tristate
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 temp_ticks_o[5]
port 230 nsew signal tristate
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 temp_ticks_o[6]
port 231 nsew signal tristate
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 temp_ticks_o[7]
port 232 nsew signal tristate
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 temp_ticks_o[8]
port 233 nsew signal tristate
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 temp_ticks_o[9]
port 234 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 235 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 235 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 236 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 236 nsew ground bidirectional
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal1 5382 16626 5382 16626 0 _000_
rlabel metal1 12236 25194 12236 25194 0 _001_
rlabel metal1 8740 27302 8740 27302 0 _002_
rlabel metal3 4876 16524 4876 16524 0 _003_
rlabel metal2 6854 22134 6854 22134 0 _004_
rlabel metal1 5704 4794 5704 4794 0 _005_
rlabel metal1 8510 26350 8510 26350 0 _006_
rlabel metal1 10442 26758 10442 26758 0 _007_
rlabel metal1 11500 17714 11500 17714 0 _008_
rlabel metal2 16882 25500 16882 25500 0 _009_
rlabel metal2 17250 22440 17250 22440 0 _010_
rlabel metal1 18124 20230 18124 20230 0 _011_
rlabel metal2 6762 18258 6762 18258 0 _012_
rlabel metal2 17802 17170 17802 17170 0 _013_
rlabel metal1 20194 10744 20194 10744 0 _014_
rlabel metal1 20378 14586 20378 14586 0 _015_
rlabel metal1 4514 3706 4514 3706 0 _016_
rlabel metal1 4002 2958 4002 2958 0 _017_
rlabel metal2 3450 7072 3450 7072 0 _018_
rlabel metal2 5934 8126 5934 8126 0 _019_
rlabel metal1 4278 6222 4278 6222 0 _020_
rlabel metal1 4738 10472 4738 10472 0 _021_
rlabel metal1 5796 9622 5796 9622 0 _022_
rlabel metal1 11086 8840 11086 8840 0 _023_
rlabel metal1 18676 6630 18676 6630 0 _024_
rlabel metal1 13846 11832 13846 11832 0 _025_
rlabel metal1 15410 3128 15410 3128 0 _026_
rlabel metal1 15318 7480 15318 7480 0 _027_
rlabel metal1 16054 4216 16054 4216 0 _028_
rlabel metal1 17986 3434 17986 3434 0 _029_
rlabel metal2 9522 3536 9522 3536 0 _030_
rlabel metal1 12374 5168 12374 5168 0 _031_
rlabel metal1 6394 17034 6394 17034 0 _032_
rlabel metal1 5520 10574 5520 10574 0 _033_
rlabel metal2 9614 13906 9614 13906 0 _034_
rlabel metal2 2530 21828 2530 21828 0 _035_
rlabel metal1 2530 21012 2530 21012 0 _036_
rlabel metal1 3726 23222 3726 23222 0 _037_
rlabel metal1 12926 26826 12926 26826 0 _038_
rlabel metal2 14214 22474 14214 22474 0 _039_
rlabel metal1 13202 26758 13202 26758 0 _040_
rlabel metal2 16606 24344 16606 24344 0 _041_
rlabel metal2 17342 19244 17342 19244 0 _042_
rlabel metal2 17342 16898 17342 16898 0 _043_
rlabel metal2 16974 19890 16974 19890 0 _044_
rlabel metal2 18722 11730 18722 11730 0 _045_
rlabel metal1 18814 9418 18814 9418 0 _046_
rlabel metal1 17940 16218 17940 16218 0 _047_
rlabel metal1 3956 14518 3956 14518 0 _048_
rlabel metal1 2668 16422 2668 16422 0 _049_
rlabel metal1 11224 19890 11224 19890 0 _050_
rlabel metal2 3082 20604 3082 20604 0 _051_
rlabel metal2 8326 23290 8326 23290 0 _052_
rlabel metal1 10816 22202 10816 22202 0 _053_
rlabel metal1 9384 11662 9384 11662 0 _054_
rlabel metal1 9292 22542 9292 22542 0 _055_
rlabel metal1 15281 13702 15281 13702 0 _056_
rlabel metal2 18722 24922 18722 24922 0 _057_
rlabel metal2 18170 22338 18170 22338 0 _058_
rlabel metal2 17066 17782 17066 17782 0 _059_
rlabel metal1 17986 23018 17986 23018 0 _060_
rlabel metal2 18722 15232 18722 15232 0 _061_
rlabel metal1 19826 7922 19826 7922 0 _062_
rlabel metal1 17710 12954 17710 12954 0 _063_
rlabel metal2 39054 55318 39054 55318 0 _064_
rlabel metal2 38778 56066 38778 56066 0 _065_
rlabel metal2 31786 54706 31786 54706 0 _066_
rlabel metal1 32706 53210 32706 53210 0 _067_
rlabel viali 27096 54638 27096 54638 0 _068_
rlabel metal2 28474 55556 28474 55556 0 _069_
rlabel metal1 28658 55692 28658 55692 0 _070_
rlabel metal2 24610 56100 24610 56100 0 _071_
rlabel via1 32887 55726 32887 55726 0 _072_
rlabel metal2 38962 55420 38962 55420 0 _073_
rlabel metal1 33028 56338 33028 56338 0 _074_
rlabel via1 40799 56338 40799 56338 0 _075_
rlabel metal2 41538 54706 41538 54706 0 _076_
rlabel metal2 41814 55522 41814 55522 0 _077_
rlabel metal2 38318 55624 38318 55624 0 _078_
rlabel metal2 33350 56032 33350 56032 0 _079_
rlabel metal1 27278 56168 27278 56168 0 _080_
rlabel metal2 26634 54944 26634 54944 0 _081_
rlabel metal2 23598 55930 23598 55930 0 _082_
rlabel metal1 21988 55250 21988 55250 0 _083_
rlabel metal2 23414 55930 23414 55930 0 _084_
rlabel metal1 34362 55658 34362 55658 0 _085_
rlabel viali 33257 55726 33257 55726 0 _086_
rlabel via2 28934 55947 28934 55947 0 _087_
rlabel viali 25990 56338 25990 56338 0 _088_
rlabel metal1 27370 56440 27370 56440 0 _089_
rlabel metal1 27186 56338 27186 56338 0 _090_
rlabel metal1 35466 54570 35466 54570 0 _091_
rlabel metal1 35880 54298 35880 54298 0 _092_
rlabel metal2 34914 54264 34914 54264 0 _093_
rlabel viali 24793 54162 24793 54162 0 _094_
rlabel metal2 24794 53754 24794 53754 0 _095_
rlabel metal2 22954 54026 22954 54026 0 _096_
rlabel metal1 35650 56338 35650 56338 0 _097_
rlabel via1 35005 56338 35005 56338 0 _098_
rlabel metal1 26910 54672 26910 54672 0 _099_
rlabel viali 26726 54638 26726 54638 0 _100_
rlabel metal2 27370 54366 27370 54366 0 _101_
rlabel metal1 26634 54162 26634 54162 0 _102_
rlabel metal1 36892 56406 36892 56406 0 _103_
rlabel metal1 37306 55930 37306 55930 0 _104_
rlabel via1 28980 56341 28980 56341 0 _105_
rlabel metal2 28842 56134 28842 56134 0 _106_
rlabel metal2 29946 55930 29946 55930 0 _107_
rlabel metal2 29210 56338 29210 56338 0 _108_
rlabel metal1 38502 55624 38502 55624 0 _109_
rlabel metal2 37490 55250 37490 55250 0 _110_
rlabel metal2 31050 56134 31050 56134 0 _111_
rlabel via1 30204 56338 30204 56338 0 _112_
rlabel metal1 31326 56440 31326 56440 0 _113_
rlabel via2 28382 55675 28382 55675 0 _114_
rlabel metal1 57362 24582 57362 24582 0 _115_
rlabel metal1 57086 24582 57086 24582 0 _116_
rlabel metal2 58282 4284 58282 4284 0 _117_
rlabel metal1 57224 3502 57224 3502 0 _118_
rlabel metal1 39652 3502 39652 3502 0 _119_
rlabel metal1 57546 4080 57546 4080 0 _120_
rlabel metal1 57960 4114 57960 4114 0 _121_
rlabel metal1 56120 13158 56120 13158 0 _122_
rlabel metal2 56534 26826 56534 26826 0 _123_
rlabel metal1 57408 22066 57408 22066 0 _124_
rlabel metal1 55982 29478 55982 29478 0 _125_
rlabel metal2 57408 16560 57408 16560 0 _126_
rlabel metal1 48760 3502 48760 3502 0 _127_
rlabel metal2 54510 31552 54510 31552 0 _128_
rlabel metal1 54740 33490 54740 33490 0 _129_
rlabel metal2 52394 34782 52394 34782 0 _130_
rlabel metal1 55016 36278 55016 36278 0 _131_
rlabel metal1 54556 37638 54556 37638 0 _132_
rlabel metal1 55936 4114 55936 4114 0 _133_
rlabel metal1 56672 39270 56672 39270 0 _134_
rlabel metal1 20562 19142 20562 19142 0 _135_
rlabel metal1 3174 23834 3174 23834 0 _136_
rlabel metal1 3726 23086 3726 23086 0 _137_
rlabel metal1 8740 28050 8740 28050 0 _138_
rlabel metal1 8694 27438 8694 27438 0 _139_
rlabel metal1 3772 26962 3772 26962 0 _140_
rlabel metal1 6302 25874 6302 25874 0 _141_
rlabel metal2 5198 27642 5198 27642 0 _142_
rlabel metal1 6210 26418 6210 26418 0 _143_
rlabel metal2 9982 27982 9982 27982 0 _144_
rlabel metal2 10902 26826 10902 26826 0 _145_
rlabel metal1 17020 26758 17020 26758 0 _146_
rlabel metal2 19642 24582 19642 24582 0 _147_
rlabel metal1 18676 20434 18676 20434 0 _148_
rlabel metal1 18124 19346 18124 19346 0 _149_
rlabel metal2 18814 16388 18814 16388 0 _150_
rlabel metal1 20654 10642 20654 10642 0 _151_
rlabel metal2 20746 14212 20746 14212 0 _152_
rlabel metal2 22586 3332 22586 3332 0 _153_
rlabel metal1 22770 4624 22770 4624 0 _154_
rlabel metal1 2162 3536 2162 3536 0 _155_
rlabel metal1 3174 3434 3174 3434 0 _156_
rlabel metal2 2254 3468 2254 3468 0 _157_
rlabel metal1 3036 7378 3036 7378 0 _158_
rlabel metal1 2944 8466 2944 8466 0 _159_
rlabel metal2 2806 6460 2806 6460 0 _160_
rlabel metal1 2944 10642 2944 10642 0 _161_
rlabel metal1 2944 11118 2944 11118 0 _162_
rlabel metal1 10166 8908 10166 8908 0 _163_
rlabel metal1 19596 6426 19596 6426 0 _164_
rlabel metal1 19550 10778 19550 10778 0 _165_
rlabel metal2 19366 3468 19366 3468 0 _166_
rlabel metal1 19872 5882 19872 5882 0 _167_
rlabel metal2 18906 3910 18906 3910 0 _168_
rlabel metal1 20148 3502 20148 3502 0 _169_
rlabel metal2 22770 3910 22770 3910 0 _170_
rlabel metal2 22402 4284 22402 4284 0 _171_
rlabel metal1 20332 18802 20332 18802 0 _172_
rlabel metal1 5060 23562 5060 23562 0 _173_
rlabel metal1 2944 17170 2944 17170 0 _174_
rlabel metal1 2944 13906 2944 13906 0 _175_
rlabel metal2 2346 13498 2346 13498 0 _176_
rlabel metal2 2438 18564 2438 18564 0 _177_
rlabel metal2 2346 21114 2346 21114 0 _178_
rlabel metal2 2346 23290 2346 23290 0 _179_
rlabel metal2 12282 27132 12282 27132 0 _180_
rlabel metal1 12558 25874 12558 25874 0 _181_
rlabel metal1 13708 26962 13708 26962 0 _182_
rlabel metal1 16813 26486 16813 26486 0 _183_
rlabel metal2 18170 18054 18170 18054 0 _184_
rlabel metal1 18952 17170 18952 17170 0 _185_
rlabel metal1 17756 18394 17756 18394 0 _186_
rlabel metal1 19182 11118 19182 11118 0 _187_
rlabel metal1 20194 9554 20194 9554 0 _188_
rlabel metal1 19412 14586 19412 14586 0 _189_
rlabel metal1 19964 19686 19964 19686 0 _190_
rlabel metal2 2162 24276 2162 24276 0 _191_
rlabel metal1 2668 22406 2668 22406 0 _192_
rlabel metal2 2392 18836 2392 18836 0 _193_
rlabel metal2 11454 29818 11454 29818 0 _194_
rlabel metal2 2898 26316 2898 26316 0 _195_
rlabel metal2 2990 25738 2990 25738 0 _196_
rlabel metal2 6854 28220 6854 28220 0 _197_
rlabel metal1 9292 26962 9292 26962 0 _198_
rlabel metal2 7682 28730 7682 28730 0 _199_
rlabel metal1 16721 27914 16721 27914 0 _200_
rlabel metal2 19642 25466 19642 25466 0 _201_
rlabel metal1 19550 22202 19550 22202 0 _202_
rlabel metal1 18400 18734 18400 18734 0 _203_
rlabel metal2 19458 23494 19458 23494 0 _204_
rlabel metal1 19550 15130 19550 15130 0 _205_
rlabel metal2 22218 8636 22218 8636 0 _206_
rlabel metal1 18860 12818 18860 12818 0 _207_
rlabel metal1 9844 6358 9844 6358 0 clknet_0_reg_wr_i
rlabel metal2 5934 3264 5934 3264 0 clknet_3_0__leaf_reg_wr_i
rlabel metal2 6026 10336 6026 10336 0 clknet_3_1__leaf_reg_wr_i
rlabel metal1 16744 7378 16744 7378 0 clknet_3_2__leaf_reg_wr_i
rlabel metal1 14444 9486 14444 9486 0 clknet_3_3__leaf_reg_wr_i
rlabel metal2 5934 17408 5934 17408 0 clknet_3_4__leaf_reg_wr_i
rlabel metal2 5750 25058 5750 25058 0 clknet_3_5__leaf_reg_wr_i
rlabel metal2 17250 17476 17250 17476 0 clknet_3_6__leaf_reg_wr_i
rlabel metal2 15410 25024 15410 25024 0 clknet_3_7__leaf_reg_wr_i
rlabel metal1 56488 2414 56488 2414 0 loopback_i
rlabel metal2 57546 1520 57546 1520 0 loopback_o
rlabel metal1 1932 57426 1932 57426 0 mux0_i[0]
rlabel metal1 3266 57426 3266 57426 0 mux0_i[1]
rlabel metal1 4324 57426 4324 57426 0 mux0_i[2]
rlabel metal1 5796 57426 5796 57426 0 mux0_i[3]
rlabel metal1 6716 56882 6716 56882 0 mux0_i[4]
rlabel metal1 8234 57426 8234 57426 0 mux0_i[5]
rlabel metal1 9108 57426 9108 57426 0 mux1_i[0]
rlabel metal1 10304 57426 10304 57426 0 mux1_i[1]
rlabel metal1 11316 57562 11316 57562 0 mux1_i[2]
rlabel metal1 12696 57426 12696 57426 0 mux1_i[3]
rlabel metal1 13800 57562 13800 57562 0 mux1_i[4]
rlabel metal1 15088 57426 15088 57426 0 mux1_i[5]
rlabel metal2 16238 58388 16238 58388 0 mux2_i[0]
rlabel metal1 17480 57426 17480 57426 0 mux2_i[1]
rlabel metal1 18676 57426 18676 57426 0 mux2_i[2]
rlabel metal1 19964 57426 19964 57426 0 mux2_i[3]
rlabel metal1 21068 57426 21068 57426 0 mux2_i[4]
rlabel metal1 22264 57426 22264 57426 0 mux2_i[5]
rlabel metal1 23460 57426 23460 57426 0 mux3_i[0]
rlabel metal1 24656 57426 24656 57426 0 mux3_i[1]
rlabel metal1 25622 57562 25622 57562 0 mux3_i[2]
rlabel metal1 26818 57562 26818 57562 0 mux3_i[3]
rlabel metal1 28244 57426 28244 57426 0 mux3_i[4]
rlabel metal1 29302 57562 29302 57562 0 mux3_i[5]
rlabel metal1 30636 57426 30636 57426 0 mux4_i[0]
rlabel metal1 32062 57426 32062 57426 0 mux4_i[1]
rlabel metal1 33028 57426 33028 57426 0 mux4_i[2]
rlabel metal1 34224 57562 34224 57562 0 mux4_i[3]
rlabel metal1 35466 57426 35466 57426 0 mux4_i[4]
rlabel metal1 36708 57426 36708 57426 0 mux4_i[5]
rlabel metal1 37904 57426 37904 57426 0 mux5_i[0]
rlabel metal1 39100 57426 39100 57426 0 mux5_i[1]
rlabel metal1 40296 57426 40296 57426 0 mux5_i[2]
rlabel metal2 41354 58320 41354 58320 0 mux5_i[3]
rlabel metal2 42826 57647 42826 57647 0 mux5_i[4]
rlabel metal1 43884 57426 43884 57426 0 mux5_i[5]
rlabel metal1 45172 57426 45172 57426 0 mux6_i[0]
rlabel metal1 46276 57426 46276 57426 0 mux6_i[1]
rlabel metal1 47656 57426 47656 57426 0 mux6_i[2]
rlabel metal1 48668 57426 48668 57426 0 mux6_i[3]
rlabel metal1 50140 57426 50140 57426 0 mux6_i[4]
rlabel metal1 51152 57426 51152 57426 0 mux6_i[5]
rlabel metal1 52256 57426 52256 57426 0 mux7_i[0]
rlabel metal1 53452 57426 53452 57426 0 mux7_i[1]
rlabel metal1 54648 57426 54648 57426 0 mux7_i[2]
rlabel metal1 55844 57426 55844 57426 0 mux7_i[3]
rlabel metal1 57040 57426 57040 57426 0 mux7_i[4]
rlabel metal1 58236 57426 58236 57426 0 mux7_i[5]
rlabel metal1 24564 2346 24564 2346 0 mux_adr_i[0]
rlabel metal1 25576 2414 25576 2414 0 mux_adr_i[1]
rlabel metal2 26634 1520 26634 1520 0 mux_adr_i[2]
rlabel metal2 27738 1792 27738 1792 0 mux_o[0]
rlabel metal2 28842 1520 28842 1520 0 mux_o[1]
rlabel metal2 29946 1520 29946 1520 0 mux_o[2]
rlabel metal2 31050 1520 31050 1520 0 mux_o[3]
rlabel metal2 32154 1520 32154 1520 0 mux_o[4]
rlabel metal2 33258 1520 33258 1520 0 mux_o[5]
rlabel metal1 57178 2618 57178 2618 0 net1
rlabel metal2 11914 57018 11914 57018 0 net10
rlabel metal1 57592 29614 57592 29614 0 net100
rlabel metal1 57270 28526 57270 28526 0 net101
rlabel metal2 56994 33490 56994 33490 0 net102
rlabel metal1 58144 31858 58144 31858 0 net103
rlabel metal1 56258 34612 56258 34612 0 net104
rlabel metal1 58144 36550 58144 36550 0 net105
rlabel metal2 57454 36618 57454 36618 0 net106
rlabel metal1 56695 37978 56695 37978 0 net107
rlabel via1 57615 5746 57615 5746 0 net108
rlabel via1 56730 6290 56730 6290 0 net109
rlabel metal1 21850 55216 21850 55216 0 net11
rlabel metal1 57730 8602 57730 8602 0 net110
rlabel metal1 57776 12682 57776 12682 0 net111
rlabel metal1 57487 11186 57487 11186 0 net112
rlabel via1 57349 13362 57349 13362 0 net113
rlabel metal2 57040 38692 57040 38692 0 net114
rlabel metal1 57316 39066 57316 39066 0 net115
rlabel metal1 58098 49062 58098 49062 0 net116
rlabel metal1 57487 25330 57487 25330 0 net117
rlabel metal1 58604 41990 58604 41990 0 net118
rlabel metal2 57868 35972 57868 35972 0 net119
rlabel metal1 21390 56712 21390 56712 0 net12
rlabel metal1 57500 43622 57500 43622 0 net120
rlabel metal1 58788 44166 58788 44166 0 net121
rlabel metal1 58742 45254 58742 45254 0 net122
rlabel via1 57165 35122 57165 35122 0 net123
rlabel metal1 58420 36006 58420 36006 0 net124
rlabel metal1 55798 37876 55798 37876 0 net125
rlabel metal1 58006 15878 58006 15878 0 net126
rlabel metal1 58512 16422 58512 16422 0 net127
rlabel metal1 58236 17510 58236 17510 0 net128
rlabel metal1 58512 18054 58512 18054 0 net129
rlabel metal1 20976 55726 20976 55726 0 net13
rlabel metal1 58328 19482 58328 19482 0 net130
rlabel metal1 58420 19686 58420 19686 0 net131
rlabel metal1 57546 27506 57546 27506 0 net132
rlabel metal1 57914 38522 57914 38522 0 net133
rlabel metal2 57730 48042 57730 48042 0 net134
rlabel metal2 57454 25364 57454 25364 0 net135
rlabel metal2 56994 30838 56994 30838 0 net136
rlabel metal1 58190 28526 58190 28526 0 net137
rlabel metal1 58052 33626 58052 33626 0 net138
rlabel metal1 57270 31858 57270 31858 0 net139
rlabel metal2 20746 56916 20746 56916 0 net14
rlabel metal1 57454 55386 57454 55386 0 net140
rlabel metal1 58880 55590 58880 55590 0 net141
rlabel metal1 58374 36890 58374 36890 0 net142
rlabel metal1 56166 37910 56166 37910 0 net143
rlabel metal1 41998 2414 41998 2414 0 net144
rlabel metal1 57086 36074 57086 36074 0 net145
rlabel metal1 57960 2414 57960 2414 0 net146
rlabel metal1 27554 3026 27554 3026 0 net147
rlabel metal1 28842 2414 28842 2414 0 net148
rlabel metal1 29946 2414 29946 2414 0 net149
rlabel metal1 19895 57290 19895 57290 0 net15
rlabel metal1 31050 2414 31050 2414 0 net150
rlabel metal1 31326 3094 31326 3094 0 net151
rlabel metal1 33258 2414 33258 2414 0 net152
rlabel metal1 2254 3604 2254 3604 0 net153
rlabel metal1 2254 2822 2254 2822 0 net154
rlabel metal2 1886 12988 1886 12988 0 net155
rlabel metal1 2622 14348 2622 14348 0 net156
rlabel metal1 4554 14790 4554 14790 0 net157
rlabel metal1 22310 3604 22310 3604 0 net158
rlabel metal1 22678 4726 22678 4726 0 net159
rlabel metal2 18906 55726 18906 55726 0 net16
rlabel metal1 2346 4046 2346 4046 0 net160
rlabel metal1 4692 6766 4692 6766 0 net161
rlabel metal1 2070 6290 2070 6290 0 net162
rlabel metal2 2346 6528 2346 6528 0 net163
rlabel metal1 2392 10574 2392 10574 0 net164
rlabel metal1 2070 8942 2070 8942 0 net165
rlabel metal2 4094 9282 4094 9282 0 net166
rlabel metal1 4186 9486 4186 9486 0 net167
rlabel metal2 2438 11424 2438 11424 0 net168
rlabel metal1 2668 17646 2668 17646 0 net169
rlabel metal2 20102 57052 20102 57052 0 net17
rlabel metal2 2438 24174 2438 24174 0 net170
rlabel metal1 4186 25194 4186 25194 0 net171
rlabel metal1 19458 18326 19458 18326 0 net172
rlabel metal1 3864 27914 3864 27914 0 net173
rlabel metal1 1886 29172 1886 29172 0 net174
rlabel metal1 1886 29580 1886 29580 0 net175
rlabel metal1 2208 17646 2208 17646 0 net176
rlabel metal1 2070 18734 2070 18734 0 net177
rlabel metal2 1886 21998 1886 21998 0 net178
rlabel metal2 2254 21284 2254 21284 0 net179
rlabel metal2 21298 57018 21298 57018 0 net18
rlabel metal1 1978 20910 1978 20910 0 net180
rlabel metal1 1886 21964 1886 21964 0 net181
rlabel metal1 1886 23052 1886 23052 0 net182
rlabel metal2 3542 24480 3542 24480 0 net183
rlabel metal1 3358 24786 3358 24786 0 net184
rlabel metal1 2438 22678 2438 22678 0 net185
rlabel metal1 2622 38726 2622 38726 0 net186
rlabel metal1 2162 39406 2162 39406 0 net187
rlabel metal1 4370 40358 4370 40358 0 net188
rlabel metal1 2162 41106 2162 41106 0 net189
rlabel metal2 30406 56848 30406 56848 0 net19
rlabel metal1 2162 42194 2162 42194 0 net190
rlabel metal1 2162 42670 2162 42670 0 net191
rlabel metal1 2208 19754 2208 19754 0 net192
rlabel metal1 2162 32402 2162 32402 0 net193
rlabel metal2 5612 21420 5612 21420 0 net194
rlabel metal1 6348 21114 6348 21114 0 net195
rlabel metal1 1886 34544 1886 34544 0 net196
rlabel metal1 2162 35666 2162 35666 0 net197
rlabel metal1 2162 36142 2162 36142 0 net198
rlabel metal2 2438 36992 2438 36992 0 net199
rlabel metal1 4531 57562 4531 57562 0 net2
rlabel metal2 25070 56542 25070 56542 0 net20
rlabel metal2 2438 37536 2438 37536 0 net200
rlabel metal1 4646 24038 4646 24038 0 net201
rlabel metal1 5566 19924 5566 19924 0 net202
rlabel metal1 19274 21658 19274 21658 0 net203
rlabel metal1 3266 18190 3266 18190 0 net204
rlabel metal2 18538 17459 18538 17459 0 net205
rlabel metal1 2162 55250 2162 55250 0 net206
rlabel metal1 2116 55726 2116 55726 0 net207
rlabel metal1 4324 44166 4324 44166 0 net208
rlabel metal1 2162 45458 2162 45458 0 net209
rlabel metal1 24932 56338 24932 56338 0 net21
rlabel metal1 2990 27506 2990 27506 0 net210
rlabel metal1 3956 27098 3956 27098 0 net211
rlabel metal1 5198 28186 5198 28186 0 net212
rlabel metal1 5750 26486 5750 26486 0 net213
rlabel metal1 2162 49198 2162 49198 0 net214
rlabel metal2 2024 31620 2024 31620 0 net215
rlabel metal1 4278 25398 4278 25398 0 net216
rlabel metal1 37858 3094 37858 3094 0 net217
rlabel metal1 38594 2414 38594 2414 0 net218
rlabel metal2 38962 2890 38962 2890 0 net219
rlabel metal1 25852 54162 25852 54162 0 net22
rlabel metal1 40434 2958 40434 2958 0 net220
rlabel metal2 41906 2176 41906 2176 0 net221
rlabel metal1 42964 2414 42964 2414 0 net222
rlabel metal1 43700 2414 43700 2414 0 net223
rlabel metal1 55062 2414 55062 2414 0 net224
rlabel metal1 56074 3366 56074 3366 0 net225
rlabel metal2 44850 3366 44850 3366 0 net226
rlabel metal2 45770 2890 45770 2890 0 net227
rlabel metal1 46874 2448 46874 2448 0 net228
rlabel metal1 48208 2414 48208 2414 0 net229
rlabel metal2 26174 55930 26174 55930 0 net23
rlabel metal1 49312 2414 49312 2414 0 net230
rlabel metal2 50646 2686 50646 2686 0 net231
rlabel metal1 51428 2414 51428 2414 0 net232
rlabel metal1 52670 2414 52670 2414 0 net233
rlabel metal1 53958 2414 53958 2414 0 net234
rlabel metal1 5665 3434 5665 3434 0 net235
rlabel metal2 5198 13090 5198 13090 0 net236
rlabel metal1 12236 3094 12236 3094 0 net237
rlabel metal1 17066 13192 17066 13192 0 net238
rlabel metal1 5290 18292 5290 18292 0 net239
rlabel metal2 28382 56508 28382 56508 0 net24
rlabel metal2 5014 22848 5014 22848 0 net240
rlabel metal2 11822 24684 11822 24684 0 net241
rlabel metal2 14858 21930 14858 21930 0 net242
rlabel metal1 6440 3434 6440 3434 0 net243
rlabel metal2 29762 57052 29762 57052 0 net25
rlabel metal2 32338 56814 32338 56814 0 net26
rlabel metal2 32982 56474 32982 56474 0 net27
rlabel metal1 34224 54570 34224 54570 0 net28
rlabel metal2 34730 56814 34730 56814 0 net29
rlabel metal2 3174 56525 3174 56525 0 net3
rlabel metal2 35834 56814 35834 56814 0 net30
rlabel metal2 35926 56474 35926 56474 0 net31
rlabel metal2 37674 56780 37674 56780 0 net32
rlabel metal2 38686 56780 38686 56780 0 net33
rlabel metal1 39146 57256 39146 57256 0 net34
rlabel via1 38779 56814 38779 56814 0 net35
rlabel viali 38682 55726 38682 55726 0 net36
rlabel metal1 42734 57290 42734 57290 0 net37
rlabel viali 41721 55726 41721 55726 0 net38
rlabel metal2 42734 56984 42734 56984 0 net39
rlabel metal1 5014 57222 5014 57222 0 net4
rlabel viali 43193 55250 43193 55250 0 net40
rlabel metal2 44758 56304 44758 56304 0 net41
rlabel metal1 43838 56848 43838 56848 0 net42
rlabel metal2 44666 56882 44666 56882 0 net43
rlabel metal2 52210 56508 52210 56508 0 net44
rlabel metal2 53406 56712 53406 56712 0 net45
rlabel metal2 54602 56270 54602 56270 0 net46
rlabel metal1 43562 55624 43562 55624 0 net47
rlabel metal1 43746 56780 43746 56780 0 net48
rlabel metal1 43470 56304 43470 56304 0 net49
rlabel metal2 5750 55658 5750 55658 0 net5
rlabel metal1 26956 2618 26956 2618 0 net50
rlabel metal1 32752 2550 32752 2550 0 net51
rlabel metal1 28888 2482 28888 2482 0 net52
rlabel metal2 22402 2550 22402 2550 0 net53
rlabel metal1 22172 6086 22172 6086 0 net54
rlabel metal1 3818 24106 3818 24106 0 net55
rlabel metal1 19780 23834 19780 23834 0 net56
rlabel metal1 19044 2414 19044 2414 0 net57
rlabel metal1 20240 22950 20240 22950 0 net58
rlabel metal1 20976 2414 20976 2414 0 net59
rlabel metal2 7038 56066 7038 56066 0 net6
rlabel metal1 22448 3502 22448 3502 0 net60
rlabel metal1 22632 4454 22632 4454 0 net61
rlabel metal1 2806 4182 2806 4182 0 net62
rlabel metal2 3910 15267 3910 15267 0 net63
rlabel metal1 3450 26010 3450 26010 0 net64
rlabel metal1 3450 6630 3450 6630 0 net65
rlabel metal1 3542 22950 3542 22950 0 net66
rlabel metal2 6348 22780 6348 22780 0 net67
rlabel metal1 12144 10030 12144 10030 0 net68
rlabel metal1 18032 27370 18032 27370 0 net69
rlabel metal2 8326 56576 8326 56576 0 net7
rlabel metal1 17710 2550 17710 2550 0 net70
rlabel metal1 5060 4182 5060 4182 0 net71
rlabel metal1 56626 3162 56626 3162 0 net72
rlabel metal2 55890 4692 55890 4692 0 net73
rlabel metal1 56764 2550 56764 2550 0 net74
rlabel metal1 57776 4794 57776 4794 0 net75
rlabel metal1 58098 4794 58098 4794 0 net76
rlabel metal1 58466 13362 58466 13362 0 net77
rlabel metal1 58236 21114 58236 21114 0 net78
rlabel metal2 57270 37468 57270 37468 0 net79
rlabel metal2 9338 57086 9338 57086 0 net8
rlabel metal1 57914 29274 57914 29274 0 net80
rlabel metal2 58190 23460 58190 23460 0 net81
rlabel metal1 57178 22746 57178 22746 0 net82
rlabel metal1 58466 23290 58466 23290 0 net83
rlabel metal1 57638 24310 57638 24310 0 net84
rlabel metal1 58144 24650 58144 24650 0 net85
rlabel metal1 57040 25738 57040 25738 0 net86
rlabel metal1 58144 26486 58144 26486 0 net87
rlabel metal1 58788 36074 58788 36074 0 net88
rlabel metal1 54786 37910 54786 37910 0 net89
rlabel metal2 10534 57052 10534 57052 0 net9
rlabel metal1 56534 5814 56534 5814 0 net90
rlabel metal1 55706 6358 55706 6358 0 net91
rlabel metal1 58236 8058 58236 8058 0 net92
rlabel metal2 58374 8772 58374 8772 0 net93
rlabel metal2 58374 10268 58374 10268 0 net94
rlabel metal1 58328 13294 58328 13294 0 net95
rlabel metal2 58374 29036 58374 29036 0 net96
rlabel metal1 57362 38998 57362 38998 0 net97
rlabel metal2 57270 39780 57270 39780 0 net98
rlabel metal1 58466 25330 58466 25330 0 net99
rlabel metal3 1188 4284 1188 4284 0 reg0_o[0]
rlabel metal3 1188 12444 1188 12444 0 reg0_o[10]
rlabel metal3 1188 13260 1188 13260 0 reg0_o[11]
rlabel metal3 1556 14076 1556 14076 0 reg0_o[12]
rlabel metal2 1702 14739 1702 14739 0 reg0_o[13]
rlabel metal3 1188 15708 1188 15708 0 reg0_o[14]
rlabel metal2 1702 16473 1702 16473 0 reg0_o[15]
rlabel metal3 1188 5100 1188 5100 0 reg0_o[1]
rlabel via2 1702 5899 1702 5899 0 reg0_o[2]
rlabel metal2 1702 6579 1702 6579 0 reg0_o[3]
rlabel metal3 1556 7548 1556 7548 0 reg0_o[4]
rlabel metal2 1702 8211 1702 8211 0 reg0_o[5]
rlabel via2 1702 9163 1702 9163 0 reg0_o[6]
rlabel metal2 1702 9707 1702 9707 0 reg0_o[7]
rlabel metal2 1702 10523 1702 10523 0 reg0_o[8]
rlabel metal3 1188 11628 1188 11628 0 reg0_o[9]
rlabel metal3 1556 17340 1556 17340 0 reg1_o[0]
rlabel via2 1702 25483 1702 25483 0 reg1_o[10]
rlabel metal3 1188 26316 1188 26316 0 reg1_o[11]
rlabel metal3 1188 27132 1188 27132 0 reg1_o[12]
rlabel metal3 1188 27948 1188 27948 0 reg1_o[13]
rlabel metal3 1188 28764 1188 28764 0 reg1_o[14]
rlabel metal3 1188 29580 1188 29580 0 reg1_o[15]
rlabel metal2 1702 18003 1702 18003 0 reg1_o[1]
rlabel via2 1702 18955 1702 18955 0 reg1_o[2]
rlabel metal2 1702 19635 1702 19635 0 reg1_o[3]
rlabel via2 1702 20587 1702 20587 0 reg1_o[4]
rlabel metal2 1702 21267 1702 21267 0 reg1_o[5]
rlabel via2 1702 22219 1702 22219 0 reg1_o[6]
rlabel metal3 1188 23052 1188 23052 0 reg1_o[7]
rlabel metal3 1188 23868 1188 23868 0 reg1_o[8]
rlabel metal3 1188 24684 1188 24684 0 reg1_o[9]
rlabel metal3 1188 30396 1188 30396 0 reg2_o[0]
rlabel metal3 1188 38556 1188 38556 0 reg2_o[10]
rlabel metal3 1188 39372 1188 39372 0 reg2_o[11]
rlabel metal3 1188 40188 1188 40188 0 reg2_o[12]
rlabel metal3 1188 41004 1188 41004 0 reg2_o[13]
rlabel metal3 1188 41820 1188 41820 0 reg2_o[14]
rlabel metal3 1188 42636 1188 42636 0 reg2_o[15]
rlabel metal3 1188 31212 1188 31212 0 reg2_o[1]
rlabel metal3 1188 32028 1188 32028 0 reg2_o[2]
rlabel metal3 1188 32844 1188 32844 0 reg2_o[3]
rlabel metal3 1188 33660 1188 33660 0 reg2_o[4]
rlabel metal3 1188 34476 1188 34476 0 reg2_o[5]
rlabel metal3 1188 35292 1188 35292 0 reg2_o[6]
rlabel metal3 1188 36108 1188 36108 0 reg2_o[7]
rlabel metal3 1188 36924 1188 36924 0 reg2_o[8]
rlabel metal3 1188 37740 1188 37740 0 reg2_o[9]
rlabel metal3 1188 43452 1188 43452 0 reg3_o[0]
rlabel metal3 1188 51612 1188 51612 0 reg3_o[10]
rlabel metal3 1188 52428 1188 52428 0 reg3_o[11]
rlabel metal3 1188 53244 1188 53244 0 reg3_o[12]
rlabel metal3 1188 54060 1188 54060 0 reg3_o[13]
rlabel metal3 1188 54876 1188 54876 0 reg3_o[14]
rlabel metal3 1188 55692 1188 55692 0 reg3_o[15]
rlabel metal3 1188 44268 1188 44268 0 reg3_o[1]
rlabel metal3 1188 45084 1188 45084 0 reg3_o[2]
rlabel metal3 1188 45900 1188 45900 0 reg3_o[3]
rlabel metal3 1188 46716 1188 46716 0 reg3_o[4]
rlabel metal3 1188 47532 1188 47532 0 reg3_o[5]
rlabel metal3 1188 48348 1188 48348 0 reg3_o[6]
rlabel metal3 1188 49164 1188 49164 0 reg3_o[7]
rlabel metal3 1188 49980 1188 49980 0 reg3_o[8]
rlabel metal3 1188 50796 1188 50796 0 reg3_o[9]
rlabel metal1 4600 2414 4600 2414 0 reg_adr_i[0]
rlabel metal1 5704 2414 5704 2414 0 reg_adr_i[1]
rlabel metal1 6992 2414 6992 2414 0 reg_dat_i[0]
rlabel metal1 17112 2958 17112 2958 0 reg_dat_i[10]
rlabel metal2 18906 1622 18906 1622 0 reg_dat_i[11]
rlabel metal2 20010 1761 20010 1761 0 reg_dat_i[12]
rlabel metal1 20884 2482 20884 2482 0 reg_dat_i[13]
rlabel metal1 22310 2380 22310 2380 0 reg_dat_i[14]
rlabel metal1 23276 2414 23276 2414 0 reg_dat_i[15]
rlabel metal1 7682 2822 7682 2822 0 reg_dat_i[1]
rlabel metal1 9062 3366 9062 3366 0 reg_dat_i[2]
rlabel metal1 10166 2822 10166 2822 0 reg_dat_i[3]
rlabel metal1 11132 2346 11132 2346 0 reg_dat_i[4]
rlabel metal1 12512 2414 12512 2414 0 reg_dat_i[5]
rlabel metal1 13432 2414 13432 2414 0 reg_dat_i[6]
rlabel metal1 14306 2414 14306 2414 0 reg_dat_i[7]
rlabel metal1 15686 2414 15686 2414 0 reg_dat_i[8]
rlabel metal1 16836 2346 16836 2346 0 reg_dat_i[9]
rlabel metal1 7544 3570 7544 3570 0 reg_wr_i
rlabel metal1 2392 2414 2392 2414 0 rst_n_i
rlabel metal3 58842 1020 58842 1020 0 temp0_dac_i[0]
rlabel metal3 57692 1836 57692 1836 0 temp0_dac_i[1]
rlabel metal1 57546 2380 57546 2380 0 temp0_dac_i[2]
rlabel metal2 57546 4029 57546 4029 0 temp0_dac_i[3]
rlabel metal2 58374 4437 58374 4437 0 temp0_dac_i[4]
rlabel metal2 58374 5151 58374 5151 0 temp0_dac_i[5]
rlabel metal2 58374 20757 58374 20757 0 temp0_ticks_i[0]
rlabel metal1 57040 29002 57040 29002 0 temp0_ticks_i[10]
rlabel metal1 58420 29138 58420 29138 0 temp0_ticks_i[11]
rlabel metal2 58374 21471 58374 21471 0 temp0_ticks_i[1]
rlabel metal2 58374 22423 58374 22423 0 temp0_ticks_i[2]
rlabel via2 58374 23069 58374 23069 0 temp0_ticks_i[3]
rlabel metal2 58374 24021 58374 24021 0 temp0_ticks_i[4]
rlabel metal2 58374 24735 58374 24735 0 temp0_ticks_i[5]
rlabel metal2 58374 25687 58374 25687 0 temp0_ticks_i[6]
rlabel via2 58374 26333 58374 26333 0 temp0_ticks_i[7]
rlabel metal2 58374 27047 58374 27047 0 temp0_ticks_i[8]
rlabel metal1 58420 28050 58420 28050 0 temp0_ticks_i[9]
rlabel metal2 58374 6103 58374 6103 0 temp1_dac_i[0]
rlabel via2 58374 6749 58374 6749 0 temp1_dac_i[1]
rlabel metal2 58374 7701 58374 7701 0 temp1_dac_i[2]
rlabel metal2 58190 8415 58190 8415 0 temp1_dac_i[3]
rlabel metal2 58190 9367 58190 9367 0 temp1_dac_i[4]
rlabel via2 58190 10013 58190 10013 0 temp1_dac_i[5]
rlabel metal1 58420 30362 58420 30362 0 temp1_ticks_i[0]
rlabel metal2 58374 38743 58374 38743 0 temp1_ticks_i[10]
rlabel metal1 58374 40052 58374 40052 0 temp1_ticks_i[11]
rlabel metal2 58190 31263 58190 31263 0 temp1_ticks_i[1]
rlabel metal2 58374 32215 58374 32215 0 temp1_ticks_i[2]
rlabel metal1 58098 33490 58098 33490 0 temp1_ticks_i[3]
rlabel metal2 58374 33813 58374 33813 0 temp1_ticks_i[4]
rlabel metal2 58374 34527 58374 34527 0 temp1_ticks_i[5]
rlabel metal2 58374 35479 58374 35479 0 temp1_ticks_i[6]
rlabel metal1 58144 36754 58144 36754 0 temp1_ticks_i[7]
rlabel metal2 58374 37077 58374 37077 0 temp1_ticks_i[8]
rlabel metal2 58374 37791 58374 37791 0 temp1_ticks_i[9]
rlabel metal1 58420 10642 58420 10642 0 temp2_dac_i[0]
rlabel metal2 58374 11679 58374 11679 0 temp2_dac_i[1]
rlabel metal3 58842 12444 58842 12444 0 temp2_dac_i[2]
rlabel metal1 58144 12818 58144 12818 0 temp2_dac_i[3]
rlabel metal2 58374 14229 58374 14229 0 temp2_dac_i[4]
rlabel metal2 58374 14943 58374 14943 0 temp2_dac_i[5]
rlabel metal2 58374 40341 58374 40341 0 temp2_ticks_i[0]
rlabel metal2 58374 48535 58374 48535 0 temp2_ticks_i[10]
rlabel via2 58374 49181 58374 49181 0 temp2_ticks_i[11]
rlabel metal2 58374 41055 58374 41055 0 temp2_ticks_i[1]
rlabel metal2 58374 42007 58374 42007 0 temp2_ticks_i[2]
rlabel via2 58374 42653 58374 42653 0 temp2_ticks_i[3]
rlabel metal2 58374 43605 58374 43605 0 temp2_ticks_i[4]
rlabel metal2 58374 44319 58374 44319 0 temp2_ticks_i[5]
rlabel metal2 58374 45271 58374 45271 0 temp2_ticks_i[6]
rlabel via2 58374 45917 58374 45917 0 temp2_ticks_i[7]
rlabel metal2 58374 46869 58374 46869 0 temp2_ticks_i[8]
rlabel metal2 58374 47583 58374 47583 0 temp2_ticks_i[9]
rlabel via2 58374 15691 58374 15691 0 temp3_dac_i[0]
rlabel via2 58374 16541 58374 16541 0 temp3_dac_i[1]
rlabel metal2 58374 17493 58374 17493 0 temp3_dac_i[2]
rlabel metal2 58374 18207 58374 18207 0 temp3_dac_i[3]
rlabel via2 58374 18955 58374 18955 0 temp3_dac_i[4]
rlabel via2 58374 19805 58374 19805 0 temp3_dac_i[5]
rlabel metal2 58374 50133 58374 50133 0 temp3_ticks_i[0]
rlabel metal1 58420 56338 58420 56338 0 temp3_ticks_i[10]
rlabel metal2 57546 57885 57546 57885 0 temp3_ticks_i[11]
rlabel metal2 58374 50847 58374 50847 0 temp3_ticks_i[1]
rlabel metal2 58374 51799 58374 51799 0 temp3_ticks_i[2]
rlabel via2 58374 52445 58374 52445 0 temp3_ticks_i[3]
rlabel metal2 58374 53397 58374 53397 0 temp3_ticks_i[4]
rlabel metal2 58374 54111 58374 54111 0 temp3_ticks_i[5]
rlabel metal1 57960 55250 57960 55250 0 temp3_ticks_i[6]
rlabel via2 58374 55709 58374 55709 0 temp3_ticks_i[7]
rlabel metal2 58374 56661 58374 56661 0 temp3_ticks_i[8]
rlabel metal2 57086 57069 57086 57069 0 temp3_ticks_i[9]
rlabel metal2 36570 1520 36570 1520 0 temp_dac_o[0]
rlabel metal2 37674 1520 37674 1520 0 temp_dac_o[1]
rlabel metal2 38778 1520 38778 1520 0 temp_dac_o[2]
rlabel metal2 39882 1520 39882 1520 0 temp_dac_o[3]
rlabel metal2 40986 1520 40986 1520 0 temp_dac_o[4]
rlabel metal2 42090 1520 42090 1520 0 temp_dac_o[5]
rlabel metal2 34362 1520 34362 1520 0 temp_sel_i[0]
rlabel metal2 35926 1700 35926 1700 0 temp_sel_i[1]
rlabel metal2 43194 1520 43194 1520 0 temp_ticks_o[0]
rlabel metal2 54234 1520 54234 1520 0 temp_ticks_o[10]
rlabel metal2 55338 1520 55338 1520 0 temp_ticks_o[11]
rlabel metal2 44298 1520 44298 1520 0 temp_ticks_o[1]
rlabel metal2 45402 1520 45402 1520 0 temp_ticks_o[2]
rlabel metal2 46506 1520 46506 1520 0 temp_ticks_o[3]
rlabel metal2 47610 1520 47610 1520 0 temp_ticks_o[4]
rlabel metal2 48714 1520 48714 1520 0 temp_ticks_o[5]
rlabel metal2 49818 1520 49818 1520 0 temp_ticks_o[6]
rlabel metal2 50922 1520 50922 1520 0 temp_ticks_o[7]
rlabel metal2 52026 1520 52026 1520 0 temp_ticks_o[8]
rlabel metal2 53130 1520 53130 1520 0 temp_ticks_o[9]
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
