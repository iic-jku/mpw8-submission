VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO audiodac
  CLASS BLOCK ;
  FOREIGN audiodac ;
  ORIGIN 0.000 0.000 ;
  SIZE 660.140 BY 670.860 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END clk_i
  PIN ds_n_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 494.590 666.860 494.870 670.860 ;
    END
  END ds_n_o
  PIN ds_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.770 666.860 165.050 670.860 ;
    END
  END ds_o
  PIN fifo_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END fifo_ack_o
  PIN fifo_empty_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END fifo_empty_o
  PIN fifo_full_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END fifo_full_o
  PIN fifo_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END fifo_i[0]
  PIN fifo_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END fifo_i[10]
  PIN fifo_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END fifo_i[11]
  PIN fifo_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END fifo_i[12]
  PIN fifo_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END fifo_i[13]
  PIN fifo_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END fifo_i[14]
  PIN fifo_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END fifo_i[15]
  PIN fifo_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END fifo_i[1]
  PIN fifo_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END fifo_i[2]
  PIN fifo_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END fifo_i[3]
  PIN fifo_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END fifo_i[4]
  PIN fifo_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END fifo_i[5]
  PIN fifo_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END fifo_i[6]
  PIN fifo_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END fifo_i[7]
  PIN fifo_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END fifo_i[8]
  PIN fifo_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END fifo_i[9]
  PIN fifo_rdy_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END fifo_rdy_i
  PIN mode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END mode_i
  PIN osr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END osr_i[0]
  PIN osr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END osr_i[1]
  PIN rst_n_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 613.730 0.000 614.010 4.000 ;
    END
  END rst_n_i
  PIN tst_fifo_loop_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END tst_fifo_loop_i
  PIN tst_sinegen_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END tst_sinegen_en_i
  PIN tst_sinegen_step_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END tst_sinegen_step_i[0]
  PIN tst_sinegen_step_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END tst_sinegen_step_i[1]
  PIN tst_sinegen_step_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END tst_sinegen_step_i[2]
  PIN tst_sinegen_step_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END tst_sinegen_step_i[3]
  PIN tst_sinegen_step_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END tst_sinegen_step_i[4]
  PIN tst_sinegen_step_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END tst_sinegen_step_i[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 658.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 658.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 658.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 658.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 658.480 ;
    END
  END vccd1
  PIN volume_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END volume_i[0]
  PIN volume_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END volume_i[1]
  PIN volume_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END volume_i[2]
  PIN volume_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END volume_i[3]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 658.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 658.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 658.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 658.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 654.580 658.325 ;
      LAYER met1 ;
        RECT 4.670 10.640 654.580 658.480 ;
      LAYER met2 ;
        RECT 4.690 666.580 164.490 667.490 ;
        RECT 165.330 666.580 494.310 667.490 ;
        RECT 495.150 666.580 653.100 667.490 ;
        RECT 4.690 4.280 653.100 666.580 ;
        RECT 4.690 4.000 15.450 4.280 ;
        RECT 16.290 4.000 45.350 4.280 ;
        RECT 46.190 4.000 75.250 4.280 ;
        RECT 76.090 4.000 105.150 4.280 ;
        RECT 105.990 4.000 135.050 4.280 ;
        RECT 135.890 4.000 164.950 4.280 ;
        RECT 165.790 4.000 194.850 4.280 ;
        RECT 195.690 4.000 224.750 4.280 ;
        RECT 225.590 4.000 254.650 4.280 ;
        RECT 255.490 4.000 284.550 4.280 ;
        RECT 285.390 4.000 314.450 4.280 ;
        RECT 315.290 4.000 344.350 4.280 ;
        RECT 345.190 4.000 374.250 4.280 ;
        RECT 375.090 4.000 404.150 4.280 ;
        RECT 404.990 4.000 434.050 4.280 ;
        RECT 434.890 4.000 463.950 4.280 ;
        RECT 464.790 4.000 493.850 4.280 ;
        RECT 494.690 4.000 523.750 4.280 ;
        RECT 524.590 4.000 553.650 4.280 ;
        RECT 554.490 4.000 583.550 4.280 ;
        RECT 584.390 4.000 613.450 4.280 ;
        RECT 614.290 4.000 643.350 4.280 ;
        RECT 644.190 4.000 653.100 4.280 ;
      LAYER met3 ;
        RECT 3.990 640.240 644.855 658.405 ;
        RECT 4.400 638.840 644.855 640.240 ;
        RECT 3.990 596.720 644.855 638.840 ;
        RECT 4.400 595.320 644.855 596.720 ;
        RECT 3.990 553.200 644.855 595.320 ;
        RECT 4.400 551.800 644.855 553.200 ;
        RECT 3.990 509.680 644.855 551.800 ;
        RECT 4.400 508.280 644.855 509.680 ;
        RECT 3.990 466.160 644.855 508.280 ;
        RECT 4.400 464.760 644.855 466.160 ;
        RECT 3.990 422.640 644.855 464.760 ;
        RECT 4.400 421.240 644.855 422.640 ;
        RECT 3.990 379.120 644.855 421.240 ;
        RECT 4.400 377.720 644.855 379.120 ;
        RECT 3.990 335.600 644.855 377.720 ;
        RECT 4.400 334.200 644.855 335.600 ;
        RECT 3.990 292.080 644.855 334.200 ;
        RECT 4.400 290.680 644.855 292.080 ;
        RECT 3.990 248.560 644.855 290.680 ;
        RECT 4.400 247.160 644.855 248.560 ;
        RECT 3.990 205.040 644.855 247.160 ;
        RECT 4.400 203.640 644.855 205.040 ;
        RECT 3.990 161.520 644.855 203.640 ;
        RECT 4.400 160.120 644.855 161.520 ;
        RECT 3.990 118.000 644.855 160.120 ;
        RECT 4.400 116.600 644.855 118.000 ;
        RECT 3.990 74.480 644.855 116.600 ;
        RECT 4.400 73.080 644.855 74.480 ;
        RECT 3.990 30.960 644.855 73.080 ;
        RECT 4.400 29.560 644.855 30.960 ;
        RECT 3.990 10.715 644.855 29.560 ;
      LAYER met4 ;
        RECT 24.215 47.775 97.440 550.625 ;
        RECT 99.840 47.775 174.240 550.625 ;
        RECT 176.640 47.775 251.040 550.625 ;
        RECT 253.440 47.775 327.840 550.625 ;
        RECT 330.240 47.775 404.640 550.625 ;
        RECT 407.040 47.775 481.440 550.625 ;
        RECT 483.840 47.775 511.225 550.625 ;
  END
END audiodac
END LIBRARY

