magic
tech sky130A
magscale 1 2
timestamp 1672093665
<< obsli1 >>
rect 1104 2159 131100 132209
<< obsm1 >>
rect 1104 2128 131100 132240
<< metal2 >>
rect 33046 133606 33102 134406
rect 99102 133606 99158 134406
rect 3238 0 3294 800
rect 9218 0 9274 800
rect 15198 0 15254 800
rect 21178 0 21234 800
rect 27158 0 27214 800
rect 33138 0 33194 800
rect 39118 0 39174 800
rect 45098 0 45154 800
rect 51078 0 51134 800
rect 57058 0 57114 800
rect 63038 0 63094 800
rect 69018 0 69074 800
rect 74998 0 75054 800
rect 80978 0 81034 800
rect 86958 0 87014 800
rect 92938 0 92994 800
rect 98918 0 98974 800
rect 104898 0 104954 800
rect 110878 0 110934 800
rect 116858 0 116914 800
rect 122838 0 122894 800
rect 128818 0 128874 800
<< obsm2 >>
rect 1492 133550 32990 133606
rect 33158 133550 99046 133606
rect 99214 133550 130436 133606
rect 1492 856 130436 133550
rect 1492 734 3182 856
rect 3350 734 9162 856
rect 9330 734 15142 856
rect 15310 734 21122 856
rect 21290 734 27102 856
rect 27270 734 33082 856
rect 33250 734 39062 856
rect 39230 734 45042 856
rect 45210 734 51022 856
rect 51190 734 57002 856
rect 57170 734 62982 856
rect 63150 734 68962 856
rect 69130 734 74942 856
rect 75110 734 80922 856
rect 81090 734 86902 856
rect 87070 734 92882 856
rect 93050 734 98862 856
rect 99030 734 104842 856
rect 105010 734 110822 856
rect 110990 734 116802 856
rect 116970 734 122782 856
rect 122950 734 128762 856
rect 128930 734 130436 856
<< metal3 >>
rect 0 128936 800 129056
rect 0 120096 800 120216
rect 0 111256 800 111376
rect 0 102416 800 102536
rect 0 93576 800 93696
rect 0 84736 800 84856
rect 0 75896 800 76016
rect 0 67056 800 67176
rect 0 58216 800 58336
rect 0 49376 800 49496
rect 0 40536 800 40656
rect 0 31696 800 31816
rect 0 22856 800 22976
rect 0 14016 800 14136
rect 0 5176 800 5296
<< obsm3 >>
rect 800 129136 127775 132225
rect 880 128856 127775 129136
rect 800 120296 127775 128856
rect 880 120016 127775 120296
rect 800 111456 127775 120016
rect 880 111176 127775 111456
rect 800 102616 127775 111176
rect 880 102336 127775 102616
rect 800 93776 127775 102336
rect 880 93496 127775 93776
rect 800 84936 127775 93496
rect 880 84656 127775 84936
rect 800 76096 127775 84656
rect 880 75816 127775 76096
rect 800 67256 127775 75816
rect 880 66976 127775 67256
rect 800 58416 127775 66976
rect 880 58136 127775 58416
rect 800 49576 127775 58136
rect 880 49296 127775 49576
rect 800 40736 127775 49296
rect 880 40456 127775 40736
rect 800 31896 127775 40456
rect 880 31616 127775 31896
rect 800 23056 127775 31616
rect 880 22776 127775 23056
rect 800 14216 127775 22776
rect 880 13936 127775 14216
rect 800 5376 127775 13936
rect 880 5096 127775 5376
rect 800 2143 127775 5096
<< metal4 >>
rect 4208 2128 4528 132240
rect 19568 2128 19888 132240
rect 34928 2128 35248 132240
rect 50288 2128 50608 132240
rect 65648 2128 65968 132240
rect 81008 2128 81328 132240
rect 96368 2128 96688 132240
rect 111728 2128 112048 132240
rect 127088 2128 127408 132240
<< obsm4 >>
rect 2083 5475 4128 128485
rect 4608 5475 19488 128485
rect 19968 5475 34848 128485
rect 35328 5475 50208 128485
rect 50688 5475 65568 128485
rect 66048 5475 80928 128485
rect 81408 5475 96288 128485
rect 96768 5475 111648 128485
rect 112128 5475 126533 128485
<< labels >>
rlabel metal2 s 128818 0 128874 800 6 clk_i
port 1 nsew signal input
rlabel metal2 s 99102 133606 99158 134406 6 ds_n_o
port 2 nsew signal output
rlabel metal2 s 33046 133606 33102 134406 6 ds_o
port 3 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 fifo_ack_o
port 4 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 fifo_empty_o
port 5 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 fifo_full_o
port 6 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 fifo_i[0]
port 7 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 fifo_i[10]
port 8 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 fifo_i[11]
port 9 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 fifo_i[12]
port 10 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 fifo_i[13]
port 11 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 fifo_i[14]
port 12 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 fifo_i[15]
port 13 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 fifo_i[1]
port 14 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 fifo_i[2]
port 15 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 fifo_i[3]
port 16 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 fifo_i[4]
port 17 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 fifo_i[5]
port 18 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 fifo_i[6]
port 19 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 fifo_i[7]
port 20 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 fifo_i[8]
port 21 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 fifo_i[9]
port 22 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 fifo_rdy_i
port 23 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 mode_i
port 24 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 osr_i[0]
port 25 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 osr_i[1]
port 26 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 rst_n_i
port 27 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 tst_fifo_loop_i
port 28 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 tst_sinegen_en_i
port 29 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 tst_sinegen_step_i[0]
port 30 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 tst_sinegen_step_i[1]
port 31 nsew signal input
rlabel metal3 s 0 102416 800 102536 6 tst_sinegen_step_i[2]
port 32 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 tst_sinegen_step_i[3]
port 33 nsew signal input
rlabel metal3 s 0 120096 800 120216 6 tst_sinegen_step_i[4]
port 34 nsew signal input
rlabel metal3 s 0 128936 800 129056 6 tst_sinegen_step_i[5]
port 35 nsew signal input
rlabel metal4 s 4208 2128 4528 132240 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 132240 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 132240 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 132240 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 132240 6 vccd1
port 36 nsew power bidirectional
rlabel metal3 s 0 14016 800 14136 6 volume_i[0]
port 37 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 volume_i[1]
port 38 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 volume_i[2]
port 39 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 volume_i[3]
port 40 nsew signal input
rlabel metal4 s 19568 2128 19888 132240 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 132240 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 132240 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 132240 6 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 132262 134406
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35013038
string GDS_FILE /foss/designs/openlane/audiodac/runs/foo/results/signoff/audiodac.magic.gds
string GDS_START 907054
<< end >>

