VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO audiodac
  CLASS BLOCK ;
  FOREIGN audiodac ;
  ORIGIN 0.000 0.000 ;
  SIZE 667.985 BY 678.705 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END clk_i
  PIN ds_n_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 674.705 500.850 678.705 ;
    END
  END ds_n_o
  PIN ds_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 674.705 166.890 678.705 ;
    END
  END ds_o
  PIN fifo_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 4.000 ;
    END
  END fifo_ack_o
  PIN fifo_empty_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END fifo_empty_o
  PIN fifo_full_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END fifo_full_o
  PIN fifo_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END fifo_i[0]
  PIN fifo_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END fifo_i[10]
  PIN fifo_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END fifo_i[11]
  PIN fifo_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END fifo_i[12]
  PIN fifo_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END fifo_i[13]
  PIN fifo_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END fifo_i[14]
  PIN fifo_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END fifo_i[15]
  PIN fifo_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END fifo_i[1]
  PIN fifo_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END fifo_i[2]
  PIN fifo_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END fifo_i[3]
  PIN fifo_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END fifo_i[4]
  PIN fifo_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END fifo_i[5]
  PIN fifo_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END fifo_i[6]
  PIN fifo_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END fifo_i[7]
  PIN fifo_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END fifo_i[8]
  PIN fifo_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END fifo_i[9]
  PIN fifo_rdy_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END fifo_rdy_i
  PIN mode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END mode_i
  PIN osr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END osr_i[0]
  PIN osr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END osr_i[1]
  PIN rst_n_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END rst_n_i
  PIN tst_fifo_loop_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END tst_fifo_loop_i
  PIN tst_sinegen_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END tst_sinegen_en_i
  PIN tst_sinegen_step_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END tst_sinegen_step_i[0]
  PIN tst_sinegen_step_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END tst_sinegen_step_i[1]
  PIN tst_sinegen_step_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END tst_sinegen_step_i[2]
  PIN tst_sinegen_step_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END tst_sinegen_step_i[3]
  PIN tst_sinegen_step_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END tst_sinegen_step_i[4]
  PIN tst_sinegen_step_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END tst_sinegen_step_i[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 666.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 666.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 666.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 666.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 666.640 ;
    END
  END vccd1
  PIN volume_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END volume_i[0]
  PIN volume_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END volume_i[1]
  PIN volume_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END volume_i[2]
  PIN volume_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END volume_i[3]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 666.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 666.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 666.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 666.640 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 662.400 666.485 ;
      LAYER met1 ;
        RECT 5.520 10.640 662.400 666.640 ;
      LAYER met2 ;
        RECT 7.000 674.425 166.330 674.705 ;
        RECT 167.170 674.425 500.290 674.705 ;
        RECT 501.130 674.425 660.000 674.705 ;
        RECT 7.000 4.280 660.000 674.425 ;
        RECT 7.000 3.670 14.530 4.280 ;
        RECT 15.370 3.670 44.890 4.280 ;
        RECT 45.730 3.670 75.250 4.280 ;
        RECT 76.090 3.670 105.610 4.280 ;
        RECT 106.450 3.670 135.970 4.280 ;
        RECT 136.810 3.670 166.330 4.280 ;
        RECT 167.170 3.670 196.690 4.280 ;
        RECT 197.530 3.670 227.050 4.280 ;
        RECT 227.890 3.670 257.410 4.280 ;
        RECT 258.250 3.670 287.770 4.280 ;
        RECT 288.610 3.670 318.130 4.280 ;
        RECT 318.970 3.670 348.490 4.280 ;
        RECT 349.330 3.670 378.850 4.280 ;
        RECT 379.690 3.670 409.210 4.280 ;
        RECT 410.050 3.670 439.570 4.280 ;
        RECT 440.410 3.670 469.930 4.280 ;
        RECT 470.770 3.670 500.290 4.280 ;
        RECT 501.130 3.670 530.650 4.280 ;
        RECT 531.490 3.670 561.010 4.280 ;
        RECT 561.850 3.670 591.370 4.280 ;
        RECT 592.210 3.670 621.730 4.280 ;
        RECT 622.570 3.670 652.090 4.280 ;
        RECT 652.930 3.670 660.000 4.280 ;
      LAYER met3 ;
        RECT 4.000 653.840 653.595 666.565 ;
        RECT 4.400 652.440 653.595 653.840 ;
        RECT 4.000 608.960 653.595 652.440 ;
        RECT 4.400 607.560 653.595 608.960 ;
        RECT 4.000 564.080 653.595 607.560 ;
        RECT 4.400 562.680 653.595 564.080 ;
        RECT 4.000 519.200 653.595 562.680 ;
        RECT 4.400 517.800 653.595 519.200 ;
        RECT 4.000 474.320 653.595 517.800 ;
        RECT 4.400 472.920 653.595 474.320 ;
        RECT 4.000 429.440 653.595 472.920 ;
        RECT 4.400 428.040 653.595 429.440 ;
        RECT 4.000 384.560 653.595 428.040 ;
        RECT 4.400 383.160 653.595 384.560 ;
        RECT 4.000 339.680 653.595 383.160 ;
        RECT 4.400 338.280 653.595 339.680 ;
        RECT 4.000 294.800 653.595 338.280 ;
        RECT 4.400 293.400 653.595 294.800 ;
        RECT 4.000 249.920 653.595 293.400 ;
        RECT 4.400 248.520 653.595 249.920 ;
        RECT 4.000 205.040 653.595 248.520 ;
        RECT 4.400 203.640 653.595 205.040 ;
        RECT 4.000 160.160 653.595 203.640 ;
        RECT 4.400 158.760 653.595 160.160 ;
        RECT 4.000 115.280 653.595 158.760 ;
        RECT 4.400 113.880 653.595 115.280 ;
        RECT 4.000 70.400 653.595 113.880 ;
        RECT 4.400 69.000 653.595 70.400 ;
        RECT 4.000 25.520 653.595 69.000 ;
        RECT 4.400 24.120 653.595 25.520 ;
        RECT 4.000 10.715 653.595 24.120 ;
      LAYER met4 ;
        RECT 15.935 17.175 20.640 664.865 ;
        RECT 23.040 17.175 97.440 664.865 ;
        RECT 99.840 17.175 174.240 664.865 ;
        RECT 176.640 17.175 251.040 664.865 ;
        RECT 253.440 17.175 327.840 664.865 ;
        RECT 330.240 17.175 404.640 664.865 ;
        RECT 407.040 17.175 481.440 664.865 ;
        RECT 483.840 17.175 558.240 664.865 ;
        RECT 560.640 17.175 624.385 664.865 ;
  END
END audiodac
END LIBRARY

