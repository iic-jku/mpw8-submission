// This is the unpowered netlist.
module tempsense (clk,
    conversion_finished_out,
    rst_n,
    start_conv_in,
    tick_result_out,
    vdac_result_out);
 input clk;
 output conversion_finished_out;
 input rst_n;
 input start_conv_in;
 output [11:0] tick_result_out;
 output [5:0] vdac_result_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire clknet_0_clk;
 wire net30;
 wire \dac.parallel_cells[0].vdac_batch.en_pupd ;
 wire \dac.parallel_cells[0].vdac_batch.en_vref ;
 wire \dac.parallel_cells[0].vdac_batch.npu_pd ;
 wire \dac.parallel_cells[0].vdac_batch.vout_analog ;
 wire \dac.parallel_cells[1].vdac_batch.en_pupd ;
 wire \dac.parallel_cells[1].vdac_batch.en_vref ;
 wire \dac.parallel_cells[1].vdac_batch.npu_pd ;
 wire \dac.parallel_cells[2].vdac_batch.en_pupd ;
 wire \dac.parallel_cells[2].vdac_batch.en_vref ;
 wire \dac.parallel_cells[2].vdac_batch.npu_pd ;
 wire \dac.parallel_cells[3].vdac_batch.en_pupd ;
 wire \dac.parallel_cells[3].vdac_batch.en_vref ;
 wire \dac.parallel_cells[3].vdac_batch.npu_pd ;
 wire \dac.parallel_cells[4].vdac_batch.en_pupd ;
 wire \dac.parallel_cells[4].vdac_batch.en_vref ;
 wire \dac.parallel_cells[4].vdac_batch.npu_pd ;
 wire \dac.vdac_single.en_pupd ;
 wire dcdc_trig_n_analog_w;
 wire dcdc_trigd_w;
 wire \sar.compare_end_w ;
 wire \sar.counter_r[0] ;
 wire \sar.counter_r[10] ;
 wire \sar.counter_r[11] ;
 wire \sar.counter_r[1] ;
 wire \sar.counter_r[2] ;
 wire \sar.counter_r[3] ;
 wire \sar.counter_r[4] ;
 wire \sar.counter_r[5] ;
 wire \sar.counter_r[6] ;
 wire \sar.counter_r[7] ;
 wire \sar.counter_r[9] ;
 wire \sar.current_dac_bit_r[0] ;
 wire \sar.current_dac_bit_r[1] ;
 wire \sar.current_dac_bit_r[2] ;
 wire \sar.current_dac_bit_r[3] ;
 wire \sar.current_dac_bit_r[4] ;
 wire \sar.current_dac_bit_r[5] ;
 wire \sar.dac_value_r[0] ;
 wire \sar.dac_value_r[1] ;
 wire \sar.dac_value_r[2] ;
 wire \sar.dac_value_r[3] ;
 wire \sar.dac_value_r[4] ;
 wire \sar.dac_value_r[5] ;
 wire \sar.dcdc_dat_out ;
 wire \sar.next_counter_w[0] ;
 wire \sar.next_counter_w[10] ;
 wire \sar.next_counter_w[11] ;
 wire \sar.next_counter_w[1] ;
 wire \sar.next_counter_w[2] ;
 wire \sar.next_counter_w[3] ;
 wire \sar.next_counter_w[4] ;
 wire \sar.next_counter_w[5] ;
 wire \sar.next_counter_w[6] ;
 wire \sar.next_counter_w[7] ;
 wire \sar.next_counter_w[8] ;
 wire \sar.next_counter_w[9] ;
 wire \sar.next_ticks_w[0] ;
 wire \sar.next_ticks_w[10] ;
 wire \sar.next_ticks_w[11] ;
 wire \sar.next_ticks_w[1] ;
 wire \sar.next_ticks_w[2] ;
 wire \sar.next_ticks_w[3] ;
 wire \sar.next_ticks_w[4] ;
 wire \sar.next_ticks_w[5] ;
 wire \sar.next_ticks_w[6] ;
 wire \sar.next_ticks_w[7] ;
 wire \sar.next_ticks_w[8] ;
 wire \sar.next_ticks_w[9] ;
 wire \sar.state_r[0] ;
 wire \sar.state_r[1] ;
 wire \sar.state_r[2] ;
 wire \sar.ticks_r[0] ;
 wire \sar.ticks_r[10] ;
 wire \sar.ticks_r[11] ;
 wire \sar.ticks_r[1] ;
 wire \sar.ticks_r[2] ;
 wire \sar.ticks_r[3] ;
 wire \sar.ticks_r[4] ;
 wire \sar.ticks_r[5] ;
 wire \sar.ticks_r[6] ;
 wire \sar.ticks_r[7] ;
 wire \sar.ticks_r[8] ;
 wire \sar.ticks_r[9] ;
 wire \sar.time_trigd_n_in ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sky130_fd_sc_hd__nor3b_4 _143_ (.A(\sar.state_r[2] ),
    .B(\sar.state_r[1] ),
    .C_N(\sar.state_r[0] ),
    .Y(_034_));
 sky130_fd_sc_hd__or3b_1 _144_ (.A(\sar.state_r[2] ),
    .B(\sar.state_r[0] ),
    .C_N(\sar.state_r[1] ),
    .X(_035_));
 sky130_fd_sc_hd__inv_2 _145_ (.A(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _146_ (.A(_034_),
    .B(_036_),
    .Y(\sar.dcdc_dat_out ));
 sky130_fd_sc_hd__nor3b_1 _147_ (.A(\sar.state_r[0] ),
    .B(\sar.state_r[1] ),
    .C_N(\sar.state_r[2] ),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_1 _148_ (.A(\sar.time_trigd_n_in ),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__clkbuf_4 _149_ (.A(_038_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _150_ (.A0(\sar.counter_r[0] ),
    .A1(\sar.ticks_r[0] ),
    .S(_039_),
    .X(_040_));
 sky130_fd_sc_hd__clkbuf_1 _151_ (.A(_040_),
    .X(\sar.next_ticks_w[0] ));
 sky130_fd_sc_hd__mux2_1 _152_ (.A0(\sar.counter_r[1] ),
    .A1(\sar.ticks_r[1] ),
    .S(_039_),
    .X(_041_));
 sky130_fd_sc_hd__clkbuf_1 _153_ (.A(_041_),
    .X(\sar.next_ticks_w[1] ));
 sky130_fd_sc_hd__mux2_1 _154_ (.A0(\sar.counter_r[2] ),
    .A1(\sar.ticks_r[2] ),
    .S(_039_),
    .X(_042_));
 sky130_fd_sc_hd__clkbuf_1 _155_ (.A(_042_),
    .X(\sar.next_ticks_w[2] ));
 sky130_fd_sc_hd__mux2_1 _156_ (.A0(\sar.counter_r[3] ),
    .A1(\sar.ticks_r[3] ),
    .S(_039_),
    .X(_043_));
 sky130_fd_sc_hd__clkbuf_1 _157_ (.A(_043_),
    .X(\sar.next_ticks_w[3] ));
 sky130_fd_sc_hd__mux2_1 _158_ (.A0(\sar.counter_r[4] ),
    .A1(\sar.ticks_r[4] ),
    .S(_039_),
    .X(_044_));
 sky130_fd_sc_hd__clkbuf_1 _159_ (.A(_044_),
    .X(\sar.next_ticks_w[4] ));
 sky130_fd_sc_hd__mux2_1 _160_ (.A0(\sar.counter_r[5] ),
    .A1(\sar.ticks_r[5] ),
    .S(_039_),
    .X(_045_));
 sky130_fd_sc_hd__clkbuf_1 _161_ (.A(_045_),
    .X(\sar.next_ticks_w[5] ));
 sky130_fd_sc_hd__mux2_1 _162_ (.A0(\sar.counter_r[6] ),
    .A1(\sar.ticks_r[6] ),
    .S(_039_),
    .X(_046_));
 sky130_fd_sc_hd__clkbuf_1 _163_ (.A(_046_),
    .X(\sar.next_ticks_w[6] ));
 sky130_fd_sc_hd__mux2_1 _164_ (.A0(\sar.counter_r[7] ),
    .A1(\sar.ticks_r[7] ),
    .S(_039_),
    .X(_047_));
 sky130_fd_sc_hd__clkbuf_1 _165_ (.A(_047_),
    .X(\sar.next_ticks_w[7] ));
 sky130_fd_sc_hd__mux2_1 _166_ (.A0(\sar.compare_end_w ),
    .A1(\sar.ticks_r[8] ),
    .S(_039_),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _167_ (.A(_048_),
    .X(\sar.next_ticks_w[8] ));
 sky130_fd_sc_hd__mux2_1 _168_ (.A0(\sar.counter_r[9] ),
    .A1(\sar.ticks_r[9] ),
    .S(_039_),
    .X(_049_));
 sky130_fd_sc_hd__clkbuf_1 _169_ (.A(_049_),
    .X(\sar.next_ticks_w[9] ));
 sky130_fd_sc_hd__mux2_1 _170_ (.A0(\sar.counter_r[10] ),
    .A1(\sar.ticks_r[10] ),
    .S(_038_),
    .X(_050_));
 sky130_fd_sc_hd__clkbuf_1 _171_ (.A(_050_),
    .X(\sar.next_ticks_w[10] ));
 sky130_fd_sc_hd__mux2_1 _172_ (.A0(\sar.counter_r[11] ),
    .A1(\sar.ticks_r[11] ),
    .S(_038_),
    .X(_051_));
 sky130_fd_sc_hd__clkbuf_1 _173_ (.A(_051_),
    .X(\sar.next_ticks_w[11] ));
 sky130_fd_sc_hd__and4_1 _174_ (.A(\sar.counter_r[1] ),
    .B(\sar.counter_r[0] ),
    .C(\sar.counter_r[3] ),
    .D(\sar.counter_r[2] ),
    .X(_052_));
 sky130_fd_sc_hd__clkbuf_2 _175_ (.A(_052_),
    .X(_053_));
 sky130_fd_sc_hd__and4_1 _176_ (.A(\sar.counter_r[5] ),
    .B(\sar.counter_r[4] ),
    .C(\sar.counter_r[7] ),
    .D(\sar.counter_r[6] ),
    .X(_054_));
 sky130_fd_sc_hd__and2_1 _177_ (.A(\sar.counter_r[9] ),
    .B(\sar.compare_end_w ),
    .X(_055_));
 sky130_fd_sc_hd__and4_2 _178_ (.A(\sar.counter_r[10] ),
    .B(_053_),
    .C(_054_),
    .D(_055_),
    .X(_056_));
 sky130_fd_sc_hd__nand2_4 _179_ (.A(\sar.counter_r[11] ),
    .B(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__clkbuf_4 _180_ (.A(_057_),
    .X(_058_));
 sky130_fd_sc_hd__and4bb_1 _181_ (.A_N(\sar.compare_end_w ),
    .B_N(\sar.state_r[2] ),
    .C(\sar.state_r[0] ),
    .D(\sar.state_r[1] ),
    .X(_059_));
 sky130_fd_sc_hd__or2_1 _182_ (.A(_037_),
    .B(_059_),
    .X(_060_));
 sky130_fd_sc_hd__buf_2 _183_ (.A(_060_),
    .X(_061_));
 sky130_fd_sc_hd__nand3_1 _184_ (.A(\sar.counter_r[0] ),
    .B(_058_),
    .C(_061_),
    .Y(\sar.next_counter_w[0] ));
 sky130_fd_sc_hd__o21ai_1 _185_ (.A1(\sar.counter_r[1] ),
    .A2(\sar.counter_r[0] ),
    .B1(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__a21oi_1 _186_ (.A1(\sar.counter_r[1] ),
    .A2(\sar.counter_r[0] ),
    .B1(_062_),
    .Y(\sar.next_counter_w[1] ));
 sky130_fd_sc_hd__nand3_1 _187_ (.A(\sar.counter_r[1] ),
    .B(\sar.counter_r[0] ),
    .C(\sar.counter_r[2] ),
    .Y(_063_));
 sky130_fd_sc_hd__a21o_1 _188_ (.A1(\sar.counter_r[1] ),
    .A2(\sar.counter_r[0] ),
    .B1(\sar.counter_r[2] ),
    .X(_064_));
 sky130_fd_sc_hd__and3_1 _189_ (.A(_063_),
    .B(_061_),
    .C(_064_),
    .X(_065_));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(_065_),
    .X(\sar.next_counter_w[2] ));
 sky130_fd_sc_hd__a31o_1 _191_ (.A1(\sar.counter_r[1] ),
    .A2(\sar.counter_r[0] ),
    .A3(\sar.counter_r[2] ),
    .B1(\sar.counter_r[3] ),
    .X(_066_));
 sky130_fd_sc_hd__and3b_1 _192_ (.A_N(_053_),
    .B(_061_),
    .C(_066_),
    .X(_067_));
 sky130_fd_sc_hd__clkbuf_1 _193_ (.A(_067_),
    .X(\sar.next_counter_w[3] ));
 sky130_fd_sc_hd__o21ai_1 _194_ (.A1(\sar.counter_r[4] ),
    .A2(_053_),
    .B1(_061_),
    .Y(_068_));
 sky130_fd_sc_hd__a21oi_1 _195_ (.A1(\sar.counter_r[4] ),
    .A2(_053_),
    .B1(_068_),
    .Y(\sar.next_counter_w[4] ));
 sky130_fd_sc_hd__a21o_1 _196_ (.A1(\sar.counter_r[4] ),
    .A2(_053_),
    .B1(\sar.counter_r[5] ),
    .X(_069_));
 sky130_fd_sc_hd__and3_1 _197_ (.A(\sar.counter_r[5] ),
    .B(\sar.counter_r[4] ),
    .C(_053_),
    .X(_070_));
 sky130_fd_sc_hd__clkinv_2 _198_ (.A(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__and3_1 _199_ (.A(_061_),
    .B(_069_),
    .C(_071_),
    .X(_072_));
 sky130_fd_sc_hd__clkbuf_1 _200_ (.A(_072_),
    .X(\sar.next_counter_w[5] ));
 sky130_fd_sc_hd__o21ai_1 _201_ (.A1(\sar.counter_r[6] ),
    .A2(_070_),
    .B1(_061_),
    .Y(_073_));
 sky130_fd_sc_hd__a21oi_1 _202_ (.A1(\sar.counter_r[6] ),
    .A2(_070_),
    .B1(_073_),
    .Y(\sar.next_counter_w[6] ));
 sky130_fd_sc_hd__and2_1 _203_ (.A(_053_),
    .B(_054_),
    .X(_074_));
 sky130_fd_sc_hd__a21o_1 _204_ (.A1(\sar.counter_r[6] ),
    .A2(_070_),
    .B1(\sar.counter_r[7] ),
    .X(_075_));
 sky130_fd_sc_hd__and3b_1 _205_ (.A_N(_074_),
    .B(_060_),
    .C(_075_),
    .X(_076_));
 sky130_fd_sc_hd__clkbuf_1 _206_ (.A(_076_),
    .X(\sar.next_counter_w[7] ));
 sky130_fd_sc_hd__o21ai_1 _207_ (.A1(\sar.compare_end_w ),
    .A2(_074_),
    .B1(_061_),
    .Y(_077_));
 sky130_fd_sc_hd__a21oi_1 _208_ (.A1(\sar.compare_end_w ),
    .A2(_074_),
    .B1(_077_),
    .Y(\sar.next_counter_w[8] ));
 sky130_fd_sc_hd__a31o_1 _209_ (.A1(\sar.compare_end_w ),
    .A2(_053_),
    .A3(_054_),
    .B1(\sar.counter_r[9] ),
    .X(_078_));
 sky130_fd_sc_hd__nand2_1 _210_ (.A(_061_),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__a21oi_1 _211_ (.A1(_074_),
    .A2(_055_),
    .B1(_079_),
    .Y(\sar.next_counter_w[9] ));
 sky130_fd_sc_hd__a31o_1 _212_ (.A1(_053_),
    .A2(_054_),
    .A3(_055_),
    .B1(\sar.counter_r[10] ),
    .X(_080_));
 sky130_fd_sc_hd__and3b_1 _213_ (.A_N(_056_),
    .B(_060_),
    .C(_080_),
    .X(_081_));
 sky130_fd_sc_hd__clkbuf_1 _214_ (.A(_081_),
    .X(\sar.next_counter_w[10] ));
 sky130_fd_sc_hd__or2_1 _215_ (.A(\sar.counter_r[11] ),
    .B(_056_),
    .X(_082_));
 sky130_fd_sc_hd__and3_1 _216_ (.A(_058_),
    .B(_061_),
    .C(_082_),
    .X(_083_));
 sky130_fd_sc_hd__clkbuf_1 _217_ (.A(_083_),
    .X(\sar.next_counter_w[11] ));
 sky130_fd_sc_hd__or2_1 _218_ (.A(\sar.current_dac_bit_r[4] ),
    .B(\sar.dac_value_r[4] ),
    .X(_084_));
 sky130_fd_sc_hd__or2_2 _219_ (.A(_034_),
    .B(_084_),
    .X(_085_));
 sky130_fd_sc_hd__inv_2 _220_ (.A(_085_),
    .Y(\dac.parallel_cells[4].vdac_batch.npu_pd ));
 sky130_fd_sc_hd__or2_1 _221_ (.A(\sar.current_dac_bit_r[3] ),
    .B(\sar.dac_value_r[3] ),
    .X(_086_));
 sky130_fd_sc_hd__or2_1 _222_ (.A(_034_),
    .B(_086_),
    .X(_087_));
 sky130_fd_sc_hd__clkinv_2 _223_ (.A(_087_),
    .Y(\dac.parallel_cells[3].vdac_batch.npu_pd ));
 sky130_fd_sc_hd__or2_1 _224_ (.A(\sar.current_dac_bit_r[2] ),
    .B(\sar.dac_value_r[2] ),
    .X(_088_));
 sky130_fd_sc_hd__or2_1 _225_ (.A(_034_),
    .B(_088_),
    .X(_089_));
 sky130_fd_sc_hd__inv_2 _226_ (.A(_089_),
    .Y(\dac.parallel_cells[2].vdac_batch.npu_pd ));
 sky130_fd_sc_hd__or2_1 _227_ (.A(\sar.current_dac_bit_r[1] ),
    .B(\sar.dac_value_r[1] ),
    .X(_090_));
 sky130_fd_sc_hd__or2_1 _228_ (.A(_034_),
    .B(_090_),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _229_ (.A(_091_),
    .Y(\dac.parallel_cells[1].vdac_batch.npu_pd ));
 sky130_fd_sc_hd__or3_1 _230_ (.A(\sar.current_dac_bit_r[0] ),
    .B(\sar.dac_value_r[0] ),
    .C(_034_),
    .X(_092_));
 sky130_fd_sc_hd__inv_2 _231_ (.A(_092_),
    .Y(\dac.parallel_cells[0].vdac_batch.npu_pd ));
 sky130_fd_sc_hd__nor3_4 _232_ (.A(\sar.state_r[2] ),
    .B(\sar.state_r[0] ),
    .C(\sar.state_r[1] ),
    .Y(_093_));
 sky130_fd_sc_hd__or2_1 _233_ (.A(\sar.current_dac_bit_r[5] ),
    .B(\sar.dac_value_r[5] ),
    .X(_094_));
 sky130_fd_sc_hd__or2_1 _234_ (.A(_034_),
    .B(_094_),
    .X(_095_));
 sky130_fd_sc_hd__clkbuf_4 _235_ (.A(_095_),
    .X(_096_));
 sky130_fd_sc_hd__xor2_2 _236_ (.A(_085_),
    .B(_096_),
    .X(_097_));
 sky130_fd_sc_hd__nor2_4 _237_ (.A(_093_),
    .B(_097_),
    .Y(\dac.parallel_cells[4].vdac_batch.en_pupd ));
 sky130_fd_sc_hd__or3_1 _238_ (.A(\sar.state_r[2] ),
    .B(\sar.state_r[0] ),
    .C(\sar.state_r[1] ),
    .X(_098_));
 sky130_fd_sc_hd__buf_2 _239_ (.A(_098_),
    .X(_099_));
 sky130_fd_sc_hd__and2_1 _240_ (.A(_099_),
    .B(_097_),
    .X(_100_));
 sky130_fd_sc_hd__clkbuf_4 _241_ (.A(_100_),
    .X(\dac.parallel_cells[4].vdac_batch.en_vref ));
 sky130_fd_sc_hd__xor2_1 _242_ (.A(_087_),
    .B(_096_),
    .X(_101_));
 sky130_fd_sc_hd__nor2_2 _243_ (.A(_093_),
    .B(_101_),
    .Y(\dac.parallel_cells[3].vdac_batch.en_pupd ));
 sky130_fd_sc_hd__and2_1 _244_ (.A(_099_),
    .B(_101_),
    .X(_102_));
 sky130_fd_sc_hd__clkbuf_2 _245_ (.A(_102_),
    .X(\dac.parallel_cells[3].vdac_batch.en_vref ));
 sky130_fd_sc_hd__xor2_1 _246_ (.A(_089_),
    .B(_096_),
    .X(_103_));
 sky130_fd_sc_hd__nor2_1 _247_ (.A(_093_),
    .B(_103_),
    .Y(\dac.parallel_cells[2].vdac_batch.en_pupd ));
 sky130_fd_sc_hd__and2_1 _248_ (.A(_099_),
    .B(_103_),
    .X(_104_));
 sky130_fd_sc_hd__clkbuf_1 _249_ (.A(_104_),
    .X(\dac.parallel_cells[2].vdac_batch.en_vref ));
 sky130_fd_sc_hd__xor2_1 _250_ (.A(_091_),
    .B(_096_),
    .X(_105_));
 sky130_fd_sc_hd__nor2_1 _251_ (.A(_093_),
    .B(_105_),
    .Y(\dac.parallel_cells[1].vdac_batch.en_pupd ));
 sky130_fd_sc_hd__and2_1 _252_ (.A(_099_),
    .B(_105_),
    .X(_106_));
 sky130_fd_sc_hd__clkbuf_1 _253_ (.A(_106_),
    .X(\dac.parallel_cells[1].vdac_batch.en_vref ));
 sky130_fd_sc_hd__xor2_1 _254_ (.A(_092_),
    .B(_096_),
    .X(_107_));
 sky130_fd_sc_hd__nor2_1 _255_ (.A(_093_),
    .B(_107_),
    .Y(\dac.parallel_cells[0].vdac_batch.en_pupd ));
 sky130_fd_sc_hd__and2_1 _256_ (.A(_099_),
    .B(_107_),
    .X(_108_));
 sky130_fd_sc_hd__clkbuf_1 _257_ (.A(_108_),
    .X(\dac.parallel_cells[0].vdac_batch.en_vref ));
 sky130_fd_sc_hd__nor2_1 _258_ (.A(_093_),
    .B(_096_),
    .Y(\dac.vdac_single.en_pupd ));
 sky130_fd_sc_hd__mux2_1 _259_ (.A0(\sar.next_ticks_w[0] ),
    .A1(net4),
    .S(_058_),
    .X(_109_));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(_109_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _261_ (.A0(\sar.next_ticks_w[1] ),
    .A1(net7),
    .S(_058_),
    .X(_110_));
 sky130_fd_sc_hd__clkbuf_1 _262_ (.A(_110_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _263_ (.A0(\sar.next_ticks_w[2] ),
    .A1(net8),
    .S(_058_),
    .X(_111_));
 sky130_fd_sc_hd__clkbuf_1 _264_ (.A(_111_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _265_ (.A0(\sar.next_ticks_w[3] ),
    .A1(net9),
    .S(_058_),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_1 _266_ (.A(_112_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _267_ (.A0(\sar.next_ticks_w[4] ),
    .A1(net10),
    .S(_058_),
    .X(_113_));
 sky130_fd_sc_hd__clkbuf_1 _268_ (.A(_113_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(\sar.next_ticks_w[5] ),
    .A1(net11),
    .S(_058_),
    .X(_114_));
 sky130_fd_sc_hd__clkbuf_1 _270_ (.A(_114_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _271_ (.A0(\sar.next_ticks_w[6] ),
    .A1(net12),
    .S(_057_),
    .X(_115_));
 sky130_fd_sc_hd__clkbuf_1 _272_ (.A(_115_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _273_ (.A0(\sar.next_ticks_w[7] ),
    .A1(net13),
    .S(_057_),
    .X(_116_));
 sky130_fd_sc_hd__clkbuf_1 _274_ (.A(_116_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _275_ (.A0(\sar.next_ticks_w[8] ),
    .A1(net14),
    .S(_057_),
    .X(_117_));
 sky130_fd_sc_hd__clkbuf_1 _276_ (.A(_117_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _277_ (.A0(\sar.next_ticks_w[9] ),
    .A1(net15),
    .S(_057_),
    .X(_118_));
 sky130_fd_sc_hd__clkbuf_1 _278_ (.A(_118_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _279_ (.A0(\sar.next_ticks_w[10] ),
    .A1(net5),
    .S(_057_),
    .X(_119_));
 sky130_fd_sc_hd__clkbuf_1 _280_ (.A(_119_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _281_ (.A0(\sar.next_ticks_w[11] ),
    .A1(net6),
    .S(_057_),
    .X(_120_));
 sky130_fd_sc_hd__clkbuf_1 _282_ (.A(_120_),
    .X(_009_));
 sky130_fd_sc_hd__or2_1 _283_ (.A(\sar.time_trigd_n_in ),
    .B(\sar.dac_value_r[0] ),
    .X(_121_));
 sky130_fd_sc_hd__clkinv_2 _284_ (.A(\sar.compare_end_w ),
    .Y(_122_));
 sky130_fd_sc_hd__or4_1 _285_ (.A(\sar.current_dac_bit_r[3] ),
    .B(\sar.current_dac_bit_r[2] ),
    .C(\sar.current_dac_bit_r[5] ),
    .D(\sar.current_dac_bit_r[4] ),
    .X(_123_));
 sky130_fd_sc_hd__or4b_4 _286_ (.A(_122_),
    .B(_123_),
    .C(\sar.current_dac_bit_r[1] ),
    .D_N(\sar.current_dac_bit_r[0] ),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(_121_),
    .A1(net16),
    .S(_124_),
    .X(_125_));
 sky130_fd_sc_hd__clkbuf_1 _288_ (.A(_125_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(\sar.dac_value_r[1] ),
    .A1(net17),
    .S(_124_),
    .X(_126_));
 sky130_fd_sc_hd__clkbuf_1 _290_ (.A(_126_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(\sar.dac_value_r[2] ),
    .A1(net18),
    .S(_124_),
    .X(_127_));
 sky130_fd_sc_hd__clkbuf_1 _292_ (.A(_127_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(\sar.dac_value_r[3] ),
    .A1(net19),
    .S(_124_),
    .X(_128_));
 sky130_fd_sc_hd__clkbuf_1 _294_ (.A(_128_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(\sar.dac_value_r[4] ),
    .A1(net20),
    .S(_124_),
    .X(_129_));
 sky130_fd_sc_hd__clkbuf_1 _296_ (.A(_129_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _297_ (.A0(\sar.dac_value_r[5] ),
    .A1(net21),
    .S(_124_),
    .X(_130_));
 sky130_fd_sc_hd__clkbuf_1 _298_ (.A(_130_),
    .X(_015_));
 sky130_fd_sc_hd__inv_2 _299_ (.A(net3),
    .Y(_131_));
 sky130_fd_sc_hd__a22oi_1 _300_ (.A1(_131_),
    .A2(_058_),
    .B1(_093_),
    .B2(net2),
    .Y(_016_));
 sky130_fd_sc_hd__and3b_1 _301_ (.A_N(\sar.state_r[2] ),
    .B(\sar.state_r[0] ),
    .C(\sar.state_r[1] ),
    .X(_132_));
 sky130_fd_sc_hd__and3_1 _302_ (.A(\sar.compare_end_w ),
    .B(\sar.time_trigd_n_in ),
    .C(_132_),
    .X(_133_));
 sky130_fd_sc_hd__clkbuf_2 _303_ (.A(_133_),
    .X(_134_));
 sky130_fd_sc_hd__a21oi_1 _304_ (.A1(\sar.current_dac_bit_r[0] ),
    .A2(_134_),
    .B1(\sar.dac_value_r[0] ),
    .Y(_135_));
 sky130_fd_sc_hd__nor2_1 _305_ (.A(_093_),
    .B(_135_),
    .Y(_017_));
 sky130_fd_sc_hd__o211a_1 _306_ (.A1(\sar.dac_value_r[1] ),
    .A2(_134_),
    .B1(_099_),
    .C1(_090_),
    .X(_018_));
 sky130_fd_sc_hd__o211a_1 _307_ (.A1(\sar.dac_value_r[2] ),
    .A2(_134_),
    .B1(_099_),
    .C1(_088_),
    .X(_019_));
 sky130_fd_sc_hd__o211a_1 _308_ (.A1(\sar.dac_value_r[3] ),
    .A2(_134_),
    .B1(_099_),
    .C1(_086_),
    .X(_020_));
 sky130_fd_sc_hd__o211a_1 _309_ (.A1(\sar.dac_value_r[4] ),
    .A2(_134_),
    .B1(_099_),
    .C1(_084_),
    .X(_021_));
 sky130_fd_sc_hd__o211a_1 _310_ (.A1(\sar.dac_value_r[5] ),
    .A2(_134_),
    .B1(_094_),
    .C1(_099_),
    .X(_022_));
 sky130_fd_sc_hd__a21oi_2 _311_ (.A1(\sar.counter_r[11] ),
    .A2(_056_),
    .B1(_122_),
    .Y(_136_));
 sky130_fd_sc_hd__a22o_1 _312_ (.A1(_122_),
    .A2(\sar.current_dac_bit_r[0] ),
    .B1(_136_),
    .B2(\sar.current_dac_bit_r[1] ),
    .X(_023_));
 sky130_fd_sc_hd__a22o_1 _313_ (.A1(_122_),
    .A2(\sar.current_dac_bit_r[1] ),
    .B1(\sar.current_dac_bit_r[2] ),
    .B2(_136_),
    .X(_024_));
 sky130_fd_sc_hd__a22o_1 _314_ (.A1(_122_),
    .A2(\sar.current_dac_bit_r[2] ),
    .B1(_136_),
    .B2(\sar.current_dac_bit_r[3] ),
    .X(_025_));
 sky130_fd_sc_hd__a22o_1 _315_ (.A1(_122_),
    .A2(\sar.current_dac_bit_r[3] ),
    .B1(\sar.current_dac_bit_r[4] ),
    .B2(_136_),
    .X(_026_));
 sky130_fd_sc_hd__a22o_1 _316_ (.A1(_122_),
    .A2(\sar.current_dac_bit_r[4] ),
    .B1(_136_),
    .B2(\sar.current_dac_bit_r[5] ),
    .X(_027_));
 sky130_fd_sc_hd__o21ba_1 _317_ (.A1(\sar.compare_end_w ),
    .A2(\sar.current_dac_bit_r[5] ),
    .B1_N(_136_),
    .X(_028_));
 sky130_fd_sc_hd__or3_1 _318_ (.A(\sar.current_dac_bit_r[1] ),
    .B(\sar.current_dac_bit_r[0] ),
    .C(_123_),
    .X(_137_));
 sky130_fd_sc_hd__or2_1 _319_ (.A(_035_),
    .B(_137_),
    .X(_138_));
 sky130_fd_sc_hd__or2_1 _320_ (.A(net2),
    .B(_098_),
    .X(_139_));
 sky130_fd_sc_hd__nor2_1 _321_ (.A(\sar.state_r[2] ),
    .B(_034_),
    .Y(_140_));
 sky130_fd_sc_hd__a31o_1 _322_ (.A1(_138_),
    .A2(_139_),
    .A3(_140_),
    .B1(_059_),
    .X(_029_));
 sky130_fd_sc_hd__a211o_1 _323_ (.A1(_036_),
    .A2(_137_),
    .B1(_059_),
    .C1(_034_),
    .X(_030_));
 sky130_fd_sc_hd__a21bo_1 _324_ (.A1(_037_),
    .A2(_058_),
    .B1_N(_138_),
    .X(_031_));
 sky130_fd_sc_hd__dfrtp_1 _325_ (.CLK(clknet_3_5__leaf_clk),
    .D(_032_),
    .RESET_B(net24),
    .Q(net4));
 sky130_fd_sc_hd__dfrtp_1 _326_ (.CLK(clknet_3_5__leaf_clk),
    .D(_033_),
    .RESET_B(net24),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _327_ (.CLK(clknet_3_5__leaf_clk),
    .D(_000_),
    .RESET_B(net24),
    .Q(net8));
 sky130_fd_sc_hd__dfrtp_1 _328_ (.CLK(clknet_3_5__leaf_clk),
    .D(_001_),
    .RESET_B(net24),
    .Q(net9));
 sky130_fd_sc_hd__dfrtp_1 _329_ (.CLK(clknet_3_5__leaf_clk),
    .D(_002_),
    .RESET_B(net24),
    .Q(net10));
 sky130_fd_sc_hd__dfrtp_1 _330_ (.CLK(clknet_3_7__leaf_clk),
    .D(_003_),
    .RESET_B(net26),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_1 _331_ (.CLK(clknet_3_7__leaf_clk),
    .D(_004_),
    .RESET_B(net26),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _332_ (.CLK(clknet_3_6__leaf_clk),
    .D(_005_),
    .RESET_B(net26),
    .Q(net13));
 sky130_fd_sc_hd__dfrtp_1 _333_ (.CLK(clknet_3_7__leaf_clk),
    .D(_006_),
    .RESET_B(net26),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _334_ (.CLK(clknet_3_6__leaf_clk),
    .D(_007_),
    .RESET_B(net26),
    .Q(net15));
 sky130_fd_sc_hd__dfrtp_1 _335_ (.CLK(clknet_3_7__leaf_clk),
    .D(_008_),
    .RESET_B(net26),
    .Q(net5));
 sky130_fd_sc_hd__dfrtp_1 _336_ (.CLK(clknet_3_6__leaf_clk),
    .D(_009_),
    .RESET_B(net28),
    .Q(net6));
 sky130_fd_sc_hd__dfrtp_1 _337_ (.CLK(clknet_3_0__leaf_clk),
    .D(_010_),
    .RESET_B(net28),
    .Q(net16));
 sky130_fd_sc_hd__dfrtp_1 _338_ (.CLK(clknet_3_0__leaf_clk),
    .D(_011_),
    .RESET_B(net28),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _339_ (.CLK(clknet_3_0__leaf_clk),
    .D(_012_),
    .RESET_B(net28),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _340_ (.CLK(clknet_3_2__leaf_clk),
    .D(_013_),
    .RESET_B(net22),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _341_ (.CLK(clknet_3_2__leaf_clk),
    .D(_014_),
    .RESET_B(net22),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _342_ (.CLK(clknet_3_2__leaf_clk),
    .D(_015_),
    .RESET_B(net22),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _343_ (.CLK(clknet_3_4__leaf_clk),
    .D(_016_),
    .RESET_B(net25),
    .Q(net3));
 sky130_fd_sc_hd__dfstp_1 _344_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sar.next_counter_w[0] ),
    .SET_B(net25),
    .Q(\sar.counter_r[0] ));
 sky130_fd_sc_hd__dfrtp_2 _345_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sar.next_counter_w[1] ),
    .RESET_B(net25),
    .Q(\sar.counter_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _346_ (.CLK(clknet_3_5__leaf_clk),
    .D(\sar.next_counter_w[2] ),
    .RESET_B(net24),
    .Q(\sar.counter_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _347_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sar.next_counter_w[3] ),
    .RESET_B(net24),
    .Q(\sar.counter_r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _348_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sar.next_counter_w[4] ),
    .RESET_B(net25),
    .Q(\sar.counter_r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _349_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sar.next_counter_w[5] ),
    .RESET_B(net25),
    .Q(\sar.counter_r[5] ));
 sky130_fd_sc_hd__dfrtp_1 _350_ (.CLK(clknet_3_7__leaf_clk),
    .D(\sar.next_counter_w[6] ),
    .RESET_B(net26),
    .Q(\sar.counter_r[6] ));
 sky130_fd_sc_hd__dfrtp_1 _351_ (.CLK(clknet_3_7__leaf_clk),
    .D(\sar.next_counter_w[7] ),
    .RESET_B(net26),
    .Q(\sar.counter_r[7] ));
 sky130_fd_sc_hd__dfrtp_4 _352_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sar.next_counter_w[8] ),
    .RESET_B(net27),
    .Q(\sar.compare_end_w ));
 sky130_fd_sc_hd__dfrtp_1 _353_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sar.next_counter_w[9] ),
    .RESET_B(net27),
    .Q(\sar.counter_r[9] ));
 sky130_fd_sc_hd__dfrtp_1 _354_ (.CLK(clknet_3_3__leaf_clk),
    .D(\sar.next_counter_w[10] ),
    .RESET_B(net27),
    .Q(\sar.counter_r[10] ));
 sky130_fd_sc_hd__dfrtp_2 _355_ (.CLK(clknet_3_3__leaf_clk),
    .D(\sar.next_counter_w[11] ),
    .RESET_B(net27),
    .Q(\sar.counter_r[11] ));
 sky130_fd_sc_hd__dfrtp_1 _356_ (.CLK(clknet_3_5__leaf_clk),
    .D(\sar.next_ticks_w[0] ),
    .RESET_B(net24),
    .Q(\sar.ticks_r[0] ));
 sky130_fd_sc_hd__dfrtp_1 _357_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sar.next_ticks_w[1] ),
    .RESET_B(net24),
    .Q(\sar.ticks_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _358_ (.CLK(clknet_3_5__leaf_clk),
    .D(\sar.next_ticks_w[2] ),
    .RESET_B(net24),
    .Q(\sar.ticks_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _359_ (.CLK(clknet_3_5__leaf_clk),
    .D(\sar.next_ticks_w[3] ),
    .RESET_B(net25),
    .Q(\sar.ticks_r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _360_ (.CLK(clknet_3_5__leaf_clk),
    .D(\sar.next_ticks_w[4] ),
    .RESET_B(net25),
    .Q(\sar.ticks_r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _361_ (.CLK(clknet_3_7__leaf_clk),
    .D(\sar.next_ticks_w[5] ),
    .RESET_B(net26),
    .Q(\sar.ticks_r[5] ));
 sky130_fd_sc_hd__dfrtp_1 _362_ (.CLK(clknet_3_7__leaf_clk),
    .D(\sar.next_ticks_w[6] ),
    .RESET_B(net26),
    .Q(\sar.ticks_r[6] ));
 sky130_fd_sc_hd__dfrtp_1 _363_ (.CLK(clknet_3_7__leaf_clk),
    .D(\sar.next_ticks_w[7] ),
    .RESET_B(net28),
    .Q(\sar.ticks_r[7] ));
 sky130_fd_sc_hd__dfrtp_1 _364_ (.CLK(clknet_3_7__leaf_clk),
    .D(\sar.next_ticks_w[8] ),
    .RESET_B(net27),
    .Q(\sar.ticks_r[8] ));
 sky130_fd_sc_hd__dfrtp_1 _365_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sar.next_ticks_w[9] ),
    .RESET_B(net27),
    .Q(\sar.ticks_r[9] ));
 sky130_fd_sc_hd__dfrtp_1 _366_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sar.next_ticks_w[10] ),
    .RESET_B(net27),
    .Q(\sar.ticks_r[10] ));
 sky130_fd_sc_hd__dfrtp_1 _367_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sar.next_ticks_w[11] ),
    .RESET_B(net27),
    .Q(\sar.ticks_r[11] ));
 sky130_fd_sc_hd__dfrtp_1 _368_ (.CLK(clknet_3_0__leaf_clk),
    .D(_017_),
    .RESET_B(net23),
    .Q(\sar.dac_value_r[0] ));
 sky130_fd_sc_hd__dfrtp_1 _369_ (.CLK(clknet_3_0__leaf_clk),
    .D(_018_),
    .RESET_B(net22),
    .Q(\sar.dac_value_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _370_ (.CLK(clknet_3_2__leaf_clk),
    .D(_019_),
    .RESET_B(net22),
    .Q(\sar.dac_value_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _371_ (.CLK(clknet_3_2__leaf_clk),
    .D(_020_),
    .RESET_B(net22),
    .Q(\sar.dac_value_r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _372_ (.CLK(clknet_3_2__leaf_clk),
    .D(_021_),
    .RESET_B(net22),
    .Q(\sar.dac_value_r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _373_ (.CLK(clknet_3_2__leaf_clk),
    .D(_022_),
    .RESET_B(net22),
    .Q(\sar.dac_value_r[5] ));
 sky130_fd_sc_hd__dfrtp_1 _374_ (.CLK(clknet_3_3__leaf_clk),
    .D(_023_),
    .RESET_B(net23),
    .Q(\sar.current_dac_bit_r[0] ));
 sky130_fd_sc_hd__dfrtp_1 _375_ (.CLK(clknet_3_1__leaf_clk),
    .D(_024_),
    .RESET_B(net23),
    .Q(\sar.current_dac_bit_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _376_ (.CLK(clknet_3_3__leaf_clk),
    .D(_025_),
    .RESET_B(net22),
    .Q(\sar.current_dac_bit_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _377_ (.CLK(clknet_3_3__leaf_clk),
    .D(_026_),
    .RESET_B(net22),
    .Q(\sar.current_dac_bit_r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _378_ (.CLK(clknet_3_2__leaf_clk),
    .D(_027_),
    .RESET_B(net23),
    .Q(\sar.current_dac_bit_r[4] ));
 sky130_fd_sc_hd__dfstp_1 _379_ (.CLK(clknet_3_3__leaf_clk),
    .D(_028_),
    .SET_B(net23),
    .Q(\sar.current_dac_bit_r[5] ));
 sky130_fd_sc_hd__dfrtp_4 _380_ (.CLK(clknet_3_1__leaf_clk),
    .D(_029_),
    .RESET_B(net25),
    .Q(\sar.state_r[0] ));
 sky130_fd_sc_hd__dfrtp_4 _381_ (.CLK(clknet_3_1__leaf_clk),
    .D(_030_),
    .RESET_B(net27),
    .Q(\sar.state_r[1] ));
 sky130_fd_sc_hd__dfrtp_4 _382_ (.CLK(clknet_3_4__leaf_clk),
    .D(_031_),
    .RESET_B(net25),
    .Q(\sar.state_r[2] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__conb_1 \dac.vdac_single.einvp_batch[0].pupd_30  (.HI(net30));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[0].vdac_batch.einvp_batch[0].pupd  (.A(\dac.parallel_cells[0].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[0].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[0].vdac_batch.einvp_batch[0].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[0].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[1].vdac_batch.einvp_batch[0].pupd  (.A(\dac.parallel_cells[1].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[1].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[1].vdac_batch.einvp_batch[0].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[1].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[1].vdac_batch.einvp_batch[1].pupd  (.A(\dac.parallel_cells[1].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[1].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[1].vdac_batch.einvp_batch[1].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[1].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[2].vdac_batch.einvp_batch[0].pupd  (.A(\dac.parallel_cells[2].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[2].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[2].vdac_batch.einvp_batch[0].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[2].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[2].vdac_batch.einvp_batch[1].pupd  (.A(\dac.parallel_cells[2].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[2].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[2].vdac_batch.einvp_batch[1].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[2].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[2].vdac_batch.einvp_batch[2].pupd  (.A(\dac.parallel_cells[2].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[2].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[2].vdac_batch.einvp_batch[2].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[2].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[2].vdac_batch.einvp_batch[3].pupd  (.A(\dac.parallel_cells[2].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[2].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[2].vdac_batch.einvp_batch[3].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[2].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[0].pupd  (.A(\dac.parallel_cells[3].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[0].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[1].pupd  (.A(\dac.parallel_cells[3].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[1].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[2].pupd  (.A(\dac.parallel_cells[3].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[2].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[3].pupd  (.A(\dac.parallel_cells[3].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[3].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[4].pupd  (.A(\dac.parallel_cells[3].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[4].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[5].pupd  (.A(\dac.parallel_cells[3].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[5].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[6].pupd  (.A(\dac.parallel_cells[3].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[6].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[7].pupd  (.A(\dac.parallel_cells[3].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[3].vdac_batch.einvp_batch[7].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[3].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[0].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[0].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[10].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[10].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[11].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[11].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[12].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[12].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[13].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[13].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[14].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[14].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[15].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[15].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[1].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[1].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[2].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[2].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[3].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[3].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[4].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[4].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[5].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[5].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[6].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[6].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[7].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[7].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[8].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[8].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[9].pupd  (.A(\dac.parallel_cells[4].vdac_batch.npu_pd ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.parallel_cells[4].vdac_batch.einvp_batch[9].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(\dac.parallel_cells[4].vdac_batch.en_vref ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.vdac_single.einvp_batch[0].pupd  (.A(net30),
    .TE(\dac.vdac_single.en_pupd ),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 \dac.vdac_single.einvp_batch[0].vref  (.A(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .TE(net29),
    .Z(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__einvp_1 dcdc (.A(\sar.dcdc_dat_out ),
    .TE(\dac.parallel_cells[0].vdac_batch.vout_analog ),
    .Z(dcdc_trig_n_analog_w));
 sky130_fd_sc_hd__clkinv_4 inv1 (.A(dcdc_trig_n_analog_w),
    .Y(dcdc_trigd_w));
 sky130_fd_sc_hd__clkinv_4 inv2 (.A(dcdc_trigd_w),
    .Y(\sar.time_trigd_n_in ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(start_conv_in),
    .X(net2));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(conversion_finished_out));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(tick_result_out[0]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(tick_result_out[10]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(tick_result_out[11]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(tick_result_out[1]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(tick_result_out[2]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(tick_result_out[3]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(tick_result_out[4]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(tick_result_out[5]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(tick_result_out[6]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(tick_result_out[7]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(tick_result_out[8]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(tick_result_out[9]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(vdac_result_out[0]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(vdac_result_out[1]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(vdac_result_out[2]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(vdac_result_out[3]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(vdac_result_out[4]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(vdac_result_out[5]));
 sky130_fd_sc_hd__buf_4 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net28),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net28),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_4 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_4 fanout28 (.A(net1),
    .X(net28));
 sky130_fd_sc_hd__conb_1 \dac.vdac_single.einvp_batch[0].vref_29  (.LO(net29));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__168__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__164__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__160__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__154__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__152__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__150__S (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__324__A2 (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__300__A2 (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__269__S (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__267__S (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__S (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__263__S (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__S (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__S (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__A (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__B (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__305__A (.DIODE(_093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__300__B1 (.DIODE(_093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__A (.DIODE(_093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__255__A (.DIODE(_093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A (.DIODE(_093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__247__A (.DIODE(_093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A (.DIODE(_093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__A (.DIODE(_093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__310__C1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__309__B1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__308__B1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__307__B1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__306__B1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__256__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__297__S (.DIODE(_124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__S (.DIODE(_124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__293__S (.DIODE(_124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__S (.DIODE(_124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__289__S (.DIODE(_124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__287__S (.DIODE(_124_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[9].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[6].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[5].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[4].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[3].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[1].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[11].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[0].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[8].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[7].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[2].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[15].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[14].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[13].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[12].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[4].vdac_batch.einvp_batch[10].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[3].vdac_batch.einvp_batch[5].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[3].vdac_batch.einvp_batch[6].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[3].vdac_batch.einvp_batch[2].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[3].vdac_batch.einvp_batch[0].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[3].vdac_batch.einvp_batch[7].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[3].vdac_batch.einvp_batch[4].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[3].vdac_batch.einvp_batch[3].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[3].vdac_batch.einvp_batch[1].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[0].vdac_batch.einvp_batch[0].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 ANTENNA_dcdc_TE (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[2].vdac_batch.einvp_batch[1].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[2].vdac_batch.einvp_batch[0].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[2].vdac_batch.einvp_batch[2].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[2].vdac_batch.einvp_batch[3].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.vdac_single.einvp_batch[0].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[1].vdac_batch.einvp_batch[0].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_dac.parallel_cells[1].vdac_batch.einvp_batch[1].vref_A  (.DIODE(\dac.parallel_cells[0].vdac_batch.vout_analog ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(start_conv_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__336__RESET_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__363__RESET_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__337__RESET_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__338__RESET_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__339__RESET_B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(net28));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_298 ();
endmodule

