* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for adc_top abstract view
.subckt adc_top VDD VSS clk_vcm config_1_in[0] config_1_in[10] config_1_in[11] config_1_in[12]
+ config_1_in[13] config_1_in[14] config_1_in[15] config_1_in[1] config_1_in[2] config_1_in[3]
+ config_1_in[4] config_1_in[5] config_1_in[6] config_1_in[7] config_1_in[8] config_1_in[9]
+ config_2_in[0] config_2_in[10] config_2_in[11] config_2_in[12] config_2_in[13] config_2_in[14]
+ config_2_in[15] config_2_in[1] config_2_in[2] config_2_in[3] config_2_in[4] config_2_in[5]
+ config_2_in[6] config_2_in[7] config_2_in[8] config_2_in[9] conversion_finished_out
+ dummypin[0] dummypin[10] dummypin[11] dummypin[12] dummypin[13] dummypin[14] dummypin[15]
+ dummypin[1] dummypin[2] dummypin[3] dummypin[4] dummypin[5] dummypin[6] dummypin[7]
+ dummypin[8] dummypin[9] inn_analog inp_analog result_out[0] result_out[10] result_out[11]
+ result_out[12] result_out[13] result_out[14] result_out[15] result_out[1] result_out[2]
+ result_out[3] result_out[4] result_out[5] result_out[6] result_out[7] result_out[8]
+ result_out[9] rst_n start_conversion_in
.ends

* Black-box entry subcircuit for config_reg_mux abstract view
.subckt config_reg_mux loopback_i loopback_o mux0_i[0] mux0_i[1] mux0_i[2] mux0_i[3]
+ mux0_i[4] mux0_i[5] mux1_i[0] mux1_i[1] mux1_i[2] mux1_i[3] mux1_i[4] mux1_i[5]
+ mux2_i[0] mux2_i[1] mux2_i[2] mux2_i[3] mux2_i[4] mux2_i[5] mux3_i[0] mux3_i[1]
+ mux3_i[2] mux3_i[3] mux3_i[4] mux3_i[5] mux4_i[0] mux4_i[1] mux4_i[2] mux4_i[3]
+ mux4_i[4] mux4_i[5] mux5_i[0] mux5_i[1] mux5_i[2] mux5_i[3] mux5_i[4] mux5_i[5]
+ mux6_i[0] mux6_i[1] mux6_i[2] mux6_i[3] mux6_i[4] mux6_i[5] mux7_i[0] mux7_i[1]
+ mux7_i[2] mux7_i[3] mux7_i[4] mux7_i[5] mux_adr_i[0] mux_adr_i[1] mux_adr_i[2] mux_o[0]
+ mux_o[1] mux_o[2] mux_o[3] mux_o[4] mux_o[5] reg0_o[0] reg0_o[10] reg0_o[11] reg0_o[12]
+ reg0_o[13] reg0_o[14] reg0_o[15] reg0_o[1] reg0_o[2] reg0_o[3] reg0_o[4] reg0_o[5]
+ reg0_o[6] reg0_o[7] reg0_o[8] reg0_o[9] reg1_o[0] reg1_o[10] reg1_o[11] reg1_o[12]
+ reg1_o[13] reg1_o[14] reg1_o[15] reg1_o[1] reg1_o[2] reg1_o[3] reg1_o[4] reg1_o[5]
+ reg1_o[6] reg1_o[7] reg1_o[8] reg1_o[9] reg2_o[0] reg2_o[10] reg2_o[11] reg2_o[12]
+ reg2_o[13] reg2_o[14] reg2_o[15] reg2_o[1] reg2_o[2] reg2_o[3] reg2_o[4] reg2_o[5]
+ reg2_o[6] reg2_o[7] reg2_o[8] reg2_o[9] reg3_o[0] reg3_o[10] reg3_o[11] reg3_o[12]
+ reg3_o[13] reg3_o[14] reg3_o[15] reg3_o[1] reg3_o[2] reg3_o[3] reg3_o[4] reg3_o[5]
+ reg3_o[6] reg3_o[7] reg3_o[8] reg3_o[9] reg_adr_i[0] reg_adr_i[1] reg_dat_i[0] reg_dat_i[10]
+ reg_dat_i[11] reg_dat_i[12] reg_dat_i[13] reg_dat_i[14] reg_dat_i[15] reg_dat_i[1]
+ reg_dat_i[2] reg_dat_i[3] reg_dat_i[4] reg_dat_i[5] reg_dat_i[6] reg_dat_i[7] reg_dat_i[8]
+ reg_dat_i[9] reg_wr_i rst_n_i temp0_dac_i[0] temp0_dac_i[1] temp0_dac_i[2] temp0_dac_i[3]
+ temp0_dac_i[4] temp0_dac_i[5] temp0_ticks_i[0] temp0_ticks_i[10] temp0_ticks_i[11]
+ temp0_ticks_i[1] temp0_ticks_i[2] temp0_ticks_i[3] temp0_ticks_i[4] temp0_ticks_i[5]
+ temp0_ticks_i[6] temp0_ticks_i[7] temp0_ticks_i[8] temp0_ticks_i[9] temp1_dac_i[0]
+ temp1_dac_i[1] temp1_dac_i[2] temp1_dac_i[3] temp1_dac_i[4] temp1_dac_i[5] temp1_ticks_i[0]
+ temp1_ticks_i[10] temp1_ticks_i[11] temp1_ticks_i[1] temp1_ticks_i[2] temp1_ticks_i[3]
+ temp1_ticks_i[4] temp1_ticks_i[5] temp1_ticks_i[6] temp1_ticks_i[7] temp1_ticks_i[8]
+ temp1_ticks_i[9] temp2_dac_i[0] temp2_dac_i[1] temp2_dac_i[2] temp2_dac_i[3] temp2_dac_i[4]
+ temp2_dac_i[5] temp2_ticks_i[0] temp2_ticks_i[10] temp2_ticks_i[11] temp2_ticks_i[1]
+ temp2_ticks_i[2] temp2_ticks_i[3] temp2_ticks_i[4] temp2_ticks_i[5] temp2_ticks_i[6]
+ temp2_ticks_i[7] temp2_ticks_i[8] temp2_ticks_i[9] temp3_dac_i[0] temp3_dac_i[1]
+ temp3_dac_i[2] temp3_dac_i[3] temp3_dac_i[4] temp3_dac_i[5] temp3_ticks_i[0] temp3_ticks_i[10]
+ temp3_ticks_i[11] temp3_ticks_i[1] temp3_ticks_i[2] temp3_ticks_i[3] temp3_ticks_i[4]
+ temp3_ticks_i[5] temp3_ticks_i[6] temp3_ticks_i[7] temp3_ticks_i[8] temp3_ticks_i[9]
+ temp_dac_o[0] temp_dac_o[1] temp_dac_o[2] temp_dac_o[3] temp_dac_o[4] temp_dac_o[5]
+ temp_sel_i[0] temp_sel_i[1] temp_ticks_o[0] temp_ticks_o[10] temp_ticks_o[11] temp_ticks_o[1]
+ temp_ticks_o[2] temp_ticks_o[3] temp_ticks_o[4] temp_ticks_o[5] temp_ticks_o[6]
+ temp_ticks_o[7] temp_ticks_o[8] temp_ticks_o[9] vccd1 vssd1
.ends

* Black-box entry subcircuit for tempsense abstract view
.subckt tempsense clk conversion_finished_out rst_n start_conv_in tick_result_out[0]
+ tick_result_out[10] tick_result_out[11] tick_result_out[1] tick_result_out[2] tick_result_out[3]
+ tick_result_out[4] tick_result_out[5] tick_result_out[6] tick_result_out[7] tick_result_out[8]
+ tick_result_out[9] vccd1 vdac_result_out[0] vdac_result_out[1] vdac_result_out[2]
+ vdac_result_out[3] vdac_result_out[4] vdac_result_out[5] vssd1
.ends

* Black-box entry subcircuit for audiodac abstract view
.subckt audiodac clk_i ds_n_o ds_o fifo_ack_o fifo_empty_o fifo_full_o fifo_i[0] fifo_i[10]
+ fifo_i[11] fifo_i[12] fifo_i[13] fifo_i[14] fifo_i[15] fifo_i[1] fifo_i[2] fifo_i[3]
+ fifo_i[4] fifo_i[5] fifo_i[6] fifo_i[7] fifo_i[8] fifo_i[9] fifo_rdy_i mode_i osr_i[0]
+ osr_i[1] rst_n_i tst_fifo_loop_i tst_sinegen_en_i tst_sinegen_step_i[0] tst_sinegen_step_i[1]
+ tst_sinegen_step_i[2] tst_sinegen_step_i[3] tst_sinegen_step_i[4] tst_sinegen_step_i[5]
+ vccd1 volume_i[0] volume_i[1] volume_i[2] volume_i[3] vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xadc0 vccd2 vssd2 io_in[6] la_data_out[32] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[40] la_data_out[41] la_data_out[48] la_data_out[58] la_data_out[59]
+ la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[49]
+ la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[126] adc0/dummypin[0]
+ adc0/dummypin[10] adc0/dummypin[11] adc0/dummypin[12] adc0/dummypin[13] adc0/dummypin[14]
+ adc0/dummypin[15] adc0/dummypin[1] adc0/dummypin[2] adc0/dummypin[3] adc0/dummypin[4]
+ adc0/dummypin[5] adc0/dummypin[6] adc0/dummypin[7] adc0/dummypin[8] adc0/dummypin[9]
+ analog_io[24] analog_io[23] la_data_out[110] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[111] la_data_out[112]
+ la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117]
+ la_data_out[118] la_data_out[119] io_in[5] io_in[29] adc_top
Xcfg_reg0 la_data_in[127] la_data_out[127] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[126] la_data_out[15] la_data_out[64] la_data_out[65]
+ la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[110] la_data_out[111] la_data_out[112]
+ la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117]
+ la_data_out[118] la_data_out[119] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[13] la_data_out[14]
+ io_in[23] io_in[24] io_in[25] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[1] la_data_out[2] la_data_out[3] la_data_out[4]
+ la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] la_data_out[16]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[30]
+ la_data_out[31] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[32] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[40]
+ la_data_out[41] la_data_out[48] la_data_out[58] la_data_out[59] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[49] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] io_in[27] io_in[28] io_in[7] io_in[17] io_in[18]
+ io_in[19] io_in[20] io_in[21] io_in[22] io_in[8] io_in[9] io_in[10] io_in[11] io_in[12]
+ io_in[13] io_in[14] io_in[15] io_in[16] io_in[26] io_in[5] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[88]
+ la_data_out[98] la_data_out[99] la_data_out[89] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] temp1_dac_w\[0\] temp1_dac_w\[1\] temp1_dac_w\[2\] temp1_dac_w\[3\]
+ temp1_dac_w\[4\] temp1_dac_w\[5\] temp1_tick_w\[0\] temp1_tick_w\[10\] temp1_tick_w\[11\]
+ temp1_tick_w\[1\] temp1_tick_w\[2\] temp1_tick_w\[3\] temp1_tick_w\[4\] temp1_tick_w\[5\]
+ temp1_tick_w\[6\] temp1_tick_w\[7\] temp1_tick_w\[8\] temp1_tick_w\[9\] temp2_dac_w\[0\]
+ temp2_dac_w\[1\] temp2_dac_w\[2\] temp2_dac_w\[3\] temp2_dac_w\[4\] temp2_dac_w\[5\]
+ temp2_tick_w\[0\] temp2_tick_w\[10\] temp2_tick_w\[11\] temp2_tick_w\[1\] temp2_tick_w\[2\]
+ temp2_tick_w\[3\] temp2_tick_w\[4\] temp2_tick_w\[5\] temp2_tick_w\[6\] temp2_tick_w\[7\]
+ temp2_tick_w\[8\] temp2_tick_w\[9\] temp3_dac_w\[0\] temp3_dac_w\[1\] temp3_dac_w\[2\]
+ temp3_dac_w\[3\] temp3_dac_w\[4\] temp3_dac_w\[5\] temp3_tick_w\[0\] temp3_tick_w\[10\]
+ temp3_tick_w\[11\] temp3_tick_w\[1\] temp3_tick_w\[2\] temp3_tick_w\[3\] temp3_tick_w\[4\]
+ temp3_tick_w\[5\] temp3_tick_w\[6\] temp3_tick_w\[7\] temp3_tick_w\[8\] temp3_tick_w\[9\]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[7] la_data_out[8] la_data_out[76] la_data_out[86] la_data_out[87]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] vccd1 vssd1 config_reg_mux
Xtemp0 io_in[6] la_data_out[100] io_in[5] io_in[29] la_data_out[88] la_data_out[98]
+ la_data_out[99] la_data_out[89] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ vccd1 la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] vssd1 tempsense
Xtemp1 io_in[6] la_data_out[101] io_in[5] io_in[29] temp1_tick_w\[0\] temp1_tick_w\[10\]
+ temp1_tick_w\[11\] temp1_tick_w\[1\] temp1_tick_w\[2\] temp1_tick_w\[3\] temp1_tick_w\[4\]
+ temp1_tick_w\[5\] temp1_tick_w\[6\] temp1_tick_w\[7\] temp1_tick_w\[8\] temp1_tick_w\[9\]
+ vccd1 temp1_dac_w\[0\] temp1_dac_w\[1\] temp1_dac_w\[2\] temp1_dac_w\[3\] temp1_dac_w\[4\]
+ temp1_dac_w\[5\] vssd1 tempsense
Xtemp2 io_in[6] la_data_out[102] io_in[5] io_in[29] temp2_tick_w\[0\] temp2_tick_w\[10\]
+ temp2_tick_w\[11\] temp2_tick_w\[1\] temp2_tick_w\[2\] temp2_tick_w\[3\] temp2_tick_w\[4\]
+ temp2_tick_w\[5\] temp2_tick_w\[6\] temp2_tick_w\[7\] temp2_tick_w\[8\] temp2_tick_w\[9\]
+ vccd1 temp2_dac_w\[0\] temp2_dac_w\[1\] temp2_dac_w\[2\] temp2_dac_w\[3\] temp2_dac_w\[4\]
+ temp2_dac_w\[5\] vssd1 tempsense
Xtemp3 io_in[6] la_data_out[103] io_in[5] io_in[29] temp3_tick_w\[0\] temp3_tick_w\[10\]
+ temp3_tick_w\[11\] temp3_tick_w\[1\] temp3_tick_w\[2\] temp3_tick_w\[3\] temp3_tick_w\[4\]
+ temp3_tick_w\[5\] temp3_tick_w\[6\] temp3_tick_w\[7\] temp3_tick_w\[8\] temp3_tick_w\[9\]
+ vccd1 temp3_dac_w\[0\] temp3_dac_w\[1\] temp3_dac_w\[2\] temp3_dac_w\[3\] temp3_dac_w\[4\]
+ temp3_dac_w\[5\] vssd1 tempsense
Xadac0 io_in[6] la_data_out[105] la_data_out[104] la_data_out[106] la_data_out[108]
+ la_data_out[107] io_in[7] io_in[17] io_in[18] io_in[19] io_in[20] io_in[21] io_in[22]
+ io_in[8] io_in[9] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16]
+ io_in[29] la_data_out[0] la_data_out[5] la_data_out[6] io_in[5] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] vccd1 la_data_out[1] la_data_out[2] la_data_out[3]
+ la_data_out[4] vssd1 audiodac
.ends

