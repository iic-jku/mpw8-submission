VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tempsense
  CLASS BLOCK ;
  FOREIGN tempsense ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END clk
  PIN conversion_finished_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END conversion_finished_out
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END rst_n
  PIN start_conv_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END start_conv_in
  PIN tick_result_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 6.840 150.000 7.440 ;
    END
  END tick_result_out[0]
  PIN tick_result_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 129.240 150.000 129.840 ;
    END
  END tick_result_out[10]
  PIN tick_result_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 141.480 150.000 142.080 ;
    END
  END tick_result_out[11]
  PIN tick_result_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 19.080 150.000 19.680 ;
    END
  END tick_result_out[1]
  PIN tick_result_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 31.320 150.000 31.920 ;
    END
  END tick_result_out[2]
  PIN tick_result_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 43.560 150.000 44.160 ;
    END
  END tick_result_out[3]
  PIN tick_result_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 55.800 150.000 56.400 ;
    END
  END tick_result_out[4]
  PIN tick_result_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.040 150.000 68.640 ;
    END
  END tick_result_out[5]
  PIN tick_result_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 80.280 150.000 80.880 ;
    END
  END tick_result_out[6]
  PIN tick_result_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 92.520 150.000 93.120 ;
    END
  END tick_result_out[7]
  PIN tick_result_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 104.760 150.000 105.360 ;
    END
  END tick_result_out[8]
  PIN tick_result_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 146.000 117.000 150.000 117.600 ;
    END
  END tick_result_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.720 10.640 18.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.720 10.640 42.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 10.640 66.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.720 10.640 90.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 112.720 10.640 114.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.720 10.640 138.320 138.960 ;
    END
  END vccd1
  PIN vdac_result_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END vdac_result_out[0]
  PIN vdac_result_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END vdac_result_out[1]
  PIN vdac_result_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END vdac_result_out[2]
  PIN vdac_result_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END vdac_result_out[3]
  PIN vdac_result_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END vdac_result_out[4]
  PIN vdac_result_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END vdac_result_out[5]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.720 10.640 30.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 52.720 10.640 54.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.720 10.640 78.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.720 10.640 102.320 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.720 10.640 126.320 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 144.440 138.960 ;
      LAYER met2 ;
        RECT 5.610 4.280 142.510 141.965 ;
        RECT 5.610 4.000 18.670 4.280 ;
        RECT 19.510 4.000 55.930 4.280 ;
        RECT 56.770 4.000 93.190 4.280 ;
        RECT 94.030 4.000 130.450 4.280 ;
        RECT 131.290 4.000 142.510 4.280 ;
      LAYER met3 ;
        RECT 3.990 141.080 145.600 141.945 ;
        RECT 3.990 135.680 146.000 141.080 ;
        RECT 4.400 134.280 146.000 135.680 ;
        RECT 3.990 130.240 146.000 134.280 ;
        RECT 3.990 128.840 145.600 130.240 ;
        RECT 3.990 118.000 146.000 128.840 ;
        RECT 3.990 116.600 145.600 118.000 ;
        RECT 3.990 111.200 146.000 116.600 ;
        RECT 4.400 109.800 146.000 111.200 ;
        RECT 3.990 105.760 146.000 109.800 ;
        RECT 3.990 104.360 145.600 105.760 ;
        RECT 3.990 93.520 146.000 104.360 ;
        RECT 3.990 92.120 145.600 93.520 ;
        RECT 3.990 86.720 146.000 92.120 ;
        RECT 4.400 85.320 146.000 86.720 ;
        RECT 3.990 81.280 146.000 85.320 ;
        RECT 3.990 79.880 145.600 81.280 ;
        RECT 3.990 69.040 146.000 79.880 ;
        RECT 3.990 67.640 145.600 69.040 ;
        RECT 3.990 62.240 146.000 67.640 ;
        RECT 4.400 60.840 146.000 62.240 ;
        RECT 3.990 56.800 146.000 60.840 ;
        RECT 3.990 55.400 145.600 56.800 ;
        RECT 3.990 44.560 146.000 55.400 ;
        RECT 3.990 43.160 145.600 44.560 ;
        RECT 3.990 37.760 146.000 43.160 ;
        RECT 4.400 36.360 146.000 37.760 ;
        RECT 3.990 32.320 146.000 36.360 ;
        RECT 3.990 30.920 145.600 32.320 ;
        RECT 3.990 20.080 146.000 30.920 ;
        RECT 3.990 18.680 145.600 20.080 ;
        RECT 3.990 13.280 146.000 18.680 ;
        RECT 4.400 11.880 146.000 13.280 ;
        RECT 3.990 7.840 146.000 11.880 ;
        RECT 3.990 6.975 145.600 7.840 ;
  END
END tempsense
END LIBRARY

