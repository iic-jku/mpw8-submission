magic
tech sky130A
magscale 1 2
timestamp 1670619538
<< obsli1 >>
rect 1104 2159 132480 133297
<< obsm1 >>
rect 1104 2128 132480 133328
<< metal2 >>
rect 33322 134941 33378 135741
rect 100114 134941 100170 135741
rect 2962 0 3018 800
rect 9034 0 9090 800
rect 15106 0 15162 800
rect 21178 0 21234 800
rect 27250 0 27306 800
rect 33322 0 33378 800
rect 39394 0 39450 800
rect 45466 0 45522 800
rect 51538 0 51594 800
rect 57610 0 57666 800
rect 63682 0 63738 800
rect 69754 0 69810 800
rect 75826 0 75882 800
rect 81898 0 81954 800
rect 87970 0 88026 800
rect 94042 0 94098 800
rect 100114 0 100170 800
rect 106186 0 106242 800
rect 112258 0 112314 800
rect 118330 0 118386 800
rect 124402 0 124458 800
rect 130474 0 130530 800
<< obsm2 >>
rect 1400 134885 33266 134941
rect 33434 134885 100058 134941
rect 100226 134885 132000 134941
rect 1400 856 132000 134885
rect 1400 734 2906 856
rect 3074 734 8978 856
rect 9146 734 15050 856
rect 15218 734 21122 856
rect 21290 734 27194 856
rect 27362 734 33266 856
rect 33434 734 39338 856
rect 39506 734 45410 856
rect 45578 734 51482 856
rect 51650 734 57554 856
rect 57722 734 63626 856
rect 63794 734 69698 856
rect 69866 734 75770 856
rect 75938 734 81842 856
rect 82010 734 87914 856
rect 88082 734 93986 856
rect 94154 734 100058 856
rect 100226 734 106130 856
rect 106298 734 112202 856
rect 112370 734 118274 856
rect 118442 734 124346 856
rect 124514 734 130418 856
rect 130586 734 132000 856
<< metal3 >>
rect 0 130568 800 130688
rect 0 121592 800 121712
rect 0 112616 800 112736
rect 0 103640 800 103760
rect 0 94664 800 94784
rect 0 85688 800 85808
rect 0 76712 800 76832
rect 0 67736 800 67856
rect 0 58760 800 58880
rect 0 49784 800 49904
rect 0 40808 800 40928
rect 0 31832 800 31952
rect 0 22856 800 22976
rect 0 13880 800 14000
rect 0 4904 800 5024
<< obsm3 >>
rect 800 130768 130719 133313
rect 880 130488 130719 130768
rect 800 121792 130719 130488
rect 880 121512 130719 121792
rect 800 112816 130719 121512
rect 880 112536 130719 112816
rect 800 103840 130719 112536
rect 880 103560 130719 103840
rect 800 94864 130719 103560
rect 880 94584 130719 94864
rect 800 85888 130719 94584
rect 880 85608 130719 85888
rect 800 76912 130719 85608
rect 880 76632 130719 76912
rect 800 67936 130719 76632
rect 880 67656 130719 67936
rect 800 58960 130719 67656
rect 880 58680 130719 58960
rect 800 49984 130719 58680
rect 880 49704 130719 49984
rect 800 41008 130719 49704
rect 880 40728 130719 41008
rect 800 32032 130719 40728
rect 880 31752 130719 32032
rect 800 23056 130719 31752
rect 880 22776 130719 23056
rect 800 14080 130719 22776
rect 880 13800 130719 14080
rect 800 5104 130719 13800
rect 880 4824 130719 5104
rect 800 2143 130719 4824
<< metal4 >>
rect 4208 2128 4528 133328
rect 19568 2128 19888 133328
rect 34928 2128 35248 133328
rect 50288 2128 50608 133328
rect 65648 2128 65968 133328
rect 81008 2128 81328 133328
rect 96368 2128 96688 133328
rect 111728 2128 112048 133328
rect 127088 2128 127408 133328
<< obsm4 >>
rect 3187 3435 4128 132973
rect 4608 3435 19488 132973
rect 19968 3435 34848 132973
rect 35328 3435 50208 132973
rect 50688 3435 65568 132973
rect 66048 3435 80928 132973
rect 81408 3435 96288 132973
rect 96768 3435 111648 132973
rect 112128 3435 124877 132973
<< labels >>
rlabel metal2 s 130474 0 130530 800 6 clk_i
port 1 nsew signal input
rlabel metal2 s 100114 134941 100170 135741 6 ds_n_o
port 2 nsew signal output
rlabel metal2 s 33322 134941 33378 135741 6 ds_o
port 3 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 fifo_ack_o
port 4 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 fifo_empty_o
port 5 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 fifo_full_o
port 6 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 fifo_i[0]
port 7 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 fifo_i[10]
port 8 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 fifo_i[11]
port 9 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 fifo_i[12]
port 10 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 fifo_i[13]
port 11 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 fifo_i[14]
port 12 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 fifo_i[15]
port 13 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 fifo_i[1]
port 14 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 fifo_i[2]
port 15 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 fifo_i[3]
port 16 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 fifo_i[4]
port 17 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 fifo_i[5]
port 18 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 fifo_i[6]
port 19 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 fifo_i[7]
port 20 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 fifo_i[8]
port 21 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 fifo_i[9]
port 22 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 fifo_rdy_i
port 23 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 mode_i
port 24 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 osr_i[0]
port 25 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 osr_i[1]
port 26 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 rst_n_i
port 27 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 tst_fifo_loop_i
port 28 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 tst_sinegen_en_i
port 29 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 tst_sinegen_step_i[0]
port 30 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 tst_sinegen_step_i[1]
port 31 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 tst_sinegen_step_i[2]
port 32 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 tst_sinegen_step_i[3]
port 33 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 tst_sinegen_step_i[4]
port 34 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 tst_sinegen_step_i[5]
port 35 nsew signal input
rlabel metal4 s 4208 2128 4528 133328 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 133328 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 133328 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 133328 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 133328 6 vccd1
port 36 nsew power bidirectional
rlabel metal3 s 0 13880 800 14000 6 volume_i[0]
port 37 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 volume_i[1]
port 38 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 volume_i[2]
port 39 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 volume_i[3]
port 40 nsew signal input
rlabel metal4 s 19568 2128 19888 133328 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 133328 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 133328 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 133328 6 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 133597 135741
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 37097844
string GDS_FILE /home/harald/mpw8-submission/openlane/audiodac/runs/22_12_09_21_48/results/signoff/audiodac.magic.gds
string GDS_START 1037184
<< end >>

