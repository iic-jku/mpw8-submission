VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO config_reg_mux
  CLASS BLOCK ;
  FOREIGN config_reg_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN loopback_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END loopback_i
  PIN loopback_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END loopback_o
  PIN mux0_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 9.290 296.000 9.570 300.000 ;
    END
  END mux0_i[0]
  PIN mux0_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 15.270 296.000 15.550 300.000 ;
    END
  END mux0_i[1]
  PIN mux0_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.250 296.000 21.530 300.000 ;
    END
  END mux0_i[2]
  PIN mux0_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 27.230 296.000 27.510 300.000 ;
    END
  END mux0_i[3]
  PIN mux0_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 33.210 296.000 33.490 300.000 ;
    END
  END mux0_i[4]
  PIN mux0_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.190 296.000 39.470 300.000 ;
    END
  END mux0_i[5]
  PIN mux1_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 296.000 45.450 300.000 ;
    END
  END mux1_i[0]
  PIN mux1_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.150 296.000 51.430 300.000 ;
    END
  END mux1_i[1]
  PIN mux1_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 57.130 296.000 57.410 300.000 ;
    END
  END mux1_i[2]
  PIN mux1_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 63.110 296.000 63.390 300.000 ;
    END
  END mux1_i[3]
  PIN mux1_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 69.090 296.000 69.370 300.000 ;
    END
  END mux1_i[4]
  PIN mux1_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 75.070 296.000 75.350 300.000 ;
    END
  END mux1_i[5]
  PIN mux2_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.050 296.000 81.330 300.000 ;
    END
  END mux2_i[0]
  PIN mux2_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 296.000 87.310 300.000 ;
    END
  END mux2_i[1]
  PIN mux2_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 296.000 93.290 300.000 ;
    END
  END mux2_i[2]
  PIN mux2_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 98.990 296.000 99.270 300.000 ;
    END
  END mux2_i[3]
  PIN mux2_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 104.970 296.000 105.250 300.000 ;
    END
  END mux2_i[4]
  PIN mux2_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 110.950 296.000 111.230 300.000 ;
    END
  END mux2_i[5]
  PIN mux3_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.930 296.000 117.210 300.000 ;
    END
  END mux3_i[0]
  PIN mux3_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 122.910 296.000 123.190 300.000 ;
    END
  END mux3_i[1]
  PIN mux3_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 296.000 129.170 300.000 ;
    END
  END mux3_i[2]
  PIN mux3_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 134.870 296.000 135.150 300.000 ;
    END
  END mux3_i[3]
  PIN mux3_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 140.850 296.000 141.130 300.000 ;
    END
  END mux3_i[4]
  PIN mux3_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 146.830 296.000 147.110 300.000 ;
    END
  END mux3_i[5]
  PIN mux4_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 152.810 296.000 153.090 300.000 ;
    END
  END mux4_i[0]
  PIN mux4_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 158.790 296.000 159.070 300.000 ;
    END
  END mux4_i[1]
  PIN mux4_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.770 296.000 165.050 300.000 ;
    END
  END mux4_i[2]
  PIN mux4_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 296.000 171.030 300.000 ;
    END
  END mux4_i[3]
  PIN mux4_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 176.730 296.000 177.010 300.000 ;
    END
  END mux4_i[4]
  PIN mux4_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 182.710 296.000 182.990 300.000 ;
    END
  END mux4_i[5]
  PIN mux5_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 188.690 296.000 188.970 300.000 ;
    END
  END mux5_i[0]
  PIN mux5_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 194.670 296.000 194.950 300.000 ;
    END
  END mux5_i[1]
  PIN mux5_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 200.650 296.000 200.930 300.000 ;
    END
  END mux5_i[2]
  PIN mux5_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 206.630 296.000 206.910 300.000 ;
    END
  END mux5_i[3]
  PIN mux5_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 296.000 212.890 300.000 ;
    END
  END mux5_i[4]
  PIN mux5_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 218.590 296.000 218.870 300.000 ;
    END
  END mux5_i[5]
  PIN mux6_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 224.570 296.000 224.850 300.000 ;
    END
  END mux6_i[0]
  PIN mux6_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 230.550 296.000 230.830 300.000 ;
    END
  END mux6_i[1]
  PIN mux6_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 236.530 296.000 236.810 300.000 ;
    END
  END mux6_i[2]
  PIN mux6_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 242.510 296.000 242.790 300.000 ;
    END
  END mux6_i[3]
  PIN mux6_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 248.490 296.000 248.770 300.000 ;
    END
  END mux6_i[4]
  PIN mux6_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 296.000 254.750 300.000 ;
    END
  END mux6_i[5]
  PIN mux7_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 260.450 296.000 260.730 300.000 ;
    END
  END mux7_i[0]
  PIN mux7_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 266.430 296.000 266.710 300.000 ;
    END
  END mux7_i[1]
  PIN mux7_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 272.410 296.000 272.690 300.000 ;
    END
  END mux7_i[2]
  PIN mux7_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 278.390 296.000 278.670 300.000 ;
    END
  END mux7_i[3]
  PIN mux7_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 284.370 296.000 284.650 300.000 ;
    END
  END mux7_i[4]
  PIN mux7_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 290.350 296.000 290.630 300.000 ;
    END
  END mux7_i[5]
  PIN mux_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END mux_adr_i[0]
  PIN mux_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END mux_adr_i[1]
  PIN mux_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END mux_adr_i[2]
  PIN mux_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END mux_o[0]
  PIN mux_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END mux_o[1]
  PIN mux_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END mux_o[2]
  PIN mux_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END mux_o[3]
  PIN mux_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END mux_o[4]
  PIN mux_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END mux_o[5]
  PIN reg0_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END reg0_o[0]
  PIN reg0_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END reg0_o[10]
  PIN reg0_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END reg0_o[11]
  PIN reg0_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END reg0_o[12]
  PIN reg0_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END reg0_o[13]
  PIN reg0_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END reg0_o[14]
  PIN reg0_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END reg0_o[15]
  PIN reg0_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END reg0_o[1]
  PIN reg0_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END reg0_o[2]
  PIN reg0_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END reg0_o[3]
  PIN reg0_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END reg0_o[4]
  PIN reg0_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END reg0_o[5]
  PIN reg0_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END reg0_o[6]
  PIN reg0_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END reg0_o[7]
  PIN reg0_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END reg0_o[8]
  PIN reg0_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END reg0_o[9]
  PIN reg1_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END reg1_o[0]
  PIN reg1_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END reg1_o[10]
  PIN reg1_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END reg1_o[11]
  PIN reg1_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END reg1_o[12]
  PIN reg1_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END reg1_o[13]
  PIN reg1_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END reg1_o[14]
  PIN reg1_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END reg1_o[15]
  PIN reg1_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END reg1_o[1]
  PIN reg1_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END reg1_o[2]
  PIN reg1_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END reg1_o[3]
  PIN reg1_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END reg1_o[4]
  PIN reg1_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END reg1_o[5]
  PIN reg1_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END reg1_o[6]
  PIN reg1_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END reg1_o[7]
  PIN reg1_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END reg1_o[8]
  PIN reg1_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END reg1_o[9]
  PIN reg2_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END reg2_o[0]
  PIN reg2_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END reg2_o[10]
  PIN reg2_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END reg2_o[11]
  PIN reg2_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END reg2_o[12]
  PIN reg2_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END reg2_o[13]
  PIN reg2_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END reg2_o[14]
  PIN reg2_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END reg2_o[15]
  PIN reg2_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END reg2_o[1]
  PIN reg2_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END reg2_o[2]
  PIN reg2_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END reg2_o[3]
  PIN reg2_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END reg2_o[4]
  PIN reg2_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END reg2_o[5]
  PIN reg2_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END reg2_o[6]
  PIN reg2_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END reg2_o[7]
  PIN reg2_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END reg2_o[8]
  PIN reg2_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END reg2_o[9]
  PIN reg3_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END reg3_o[0]
  PIN reg3_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END reg3_o[10]
  PIN reg3_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END reg3_o[11]
  PIN reg3_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END reg3_o[12]
  PIN reg3_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END reg3_o[13]
  PIN reg3_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END reg3_o[14]
  PIN reg3_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END reg3_o[15]
  PIN reg3_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END reg3_o[1]
  PIN reg3_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END reg3_o[2]
  PIN reg3_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END reg3_o[3]
  PIN reg3_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END reg3_o[4]
  PIN reg3_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END reg3_o[5]
  PIN reg3_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END reg3_o[6]
  PIN reg3_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END reg3_o[7]
  PIN reg3_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END reg3_o[8]
  PIN reg3_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END reg3_o[9]
  PIN reg_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END reg_adr_i[0]
  PIN reg_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END reg_adr_i[1]
  PIN reg_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END reg_dat_i[0]
  PIN reg_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END reg_dat_i[10]
  PIN reg_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END reg_dat_i[11]
  PIN reg_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END reg_dat_i[12]
  PIN reg_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END reg_dat_i[13]
  PIN reg_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END reg_dat_i[14]
  PIN reg_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END reg_dat_i[15]
  PIN reg_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END reg_dat_i[1]
  PIN reg_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END reg_dat_i[2]
  PIN reg_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END reg_dat_i[3]
  PIN reg_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END reg_dat_i[4]
  PIN reg_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END reg_dat_i[5]
  PIN reg_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END reg_dat_i[6]
  PIN reg_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END reg_dat_i[7]
  PIN reg_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END reg_dat_i[8]
  PIN reg_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END reg_dat_i[9]
  PIN reg_wr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END reg_wr_i
  PIN rst_n_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END rst_n_i
  PIN temp0_dac_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.120 300.000 4.720 ;
    END
  END temp0_dac_i[0]
  PIN temp0_dac_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.200 300.000 8.800 ;
    END
  END temp0_dac_i[1]
  PIN temp0_dac_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 12.280 300.000 12.880 ;
    END
  END temp0_dac_i[2]
  PIN temp0_dac_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.360 300.000 16.960 ;
    END
  END temp0_dac_i[3]
  PIN temp0_dac_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.440 300.000 21.040 ;
    END
  END temp0_dac_i[4]
  PIN temp0_dac_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 24.520 300.000 25.120 ;
    END
  END temp0_dac_i[5]
  PIN temp0_ticks_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.040 300.000 102.640 ;
    END
  END temp0_ticks_i[0]
  PIN temp0_ticks_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.840 300.000 143.440 ;
    END
  END temp0_ticks_i[10]
  PIN temp0_ticks_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.920 300.000 147.520 ;
    END
  END temp0_ticks_i[11]
  PIN temp0_ticks_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 106.120 300.000 106.720 ;
    END
  END temp0_ticks_i[1]
  PIN temp0_ticks_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.200 300.000 110.800 ;
    END
  END temp0_ticks_i[2]
  PIN temp0_ticks_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.280 300.000 114.880 ;
    END
  END temp0_ticks_i[3]
  PIN temp0_ticks_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.360 300.000 118.960 ;
    END
  END temp0_ticks_i[4]
  PIN temp0_ticks_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.440 300.000 123.040 ;
    END
  END temp0_ticks_i[5]
  PIN temp0_ticks_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 126.520 300.000 127.120 ;
    END
  END temp0_ticks_i[6]
  PIN temp0_ticks_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.600 300.000 131.200 ;
    END
  END temp0_ticks_i[7]
  PIN temp0_ticks_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 134.680 300.000 135.280 ;
    END
  END temp0_ticks_i[8]
  PIN temp0_ticks_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.760 300.000 139.360 ;
    END
  END temp0_ticks_i[9]
  PIN temp1_dac_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 28.600 300.000 29.200 ;
    END
  END temp1_dac_i[0]
  PIN temp1_dac_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.680 300.000 33.280 ;
    END
  END temp1_dac_i[1]
  PIN temp1_dac_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.760 300.000 37.360 ;
    END
  END temp1_dac_i[2]
  PIN temp1_dac_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.840 300.000 41.440 ;
    END
  END temp1_dac_i[3]
  PIN temp1_dac_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.920 300.000 45.520 ;
    END
  END temp1_dac_i[4]
  PIN temp1_dac_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.000 300.000 49.600 ;
    END
  END temp1_dac_i[5]
  PIN temp1_ticks_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 151.000 300.000 151.600 ;
    END
  END temp1_ticks_i[0]
  PIN temp1_ticks_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 191.800 300.000 192.400 ;
    END
  END temp1_ticks_i[10]
  PIN temp1_ticks_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.880 300.000 196.480 ;
    END
  END temp1_ticks_i[11]
  PIN temp1_ticks_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 155.080 300.000 155.680 ;
    END
  END temp1_ticks_i[1]
  PIN temp1_ticks_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.160 300.000 159.760 ;
    END
  END temp1_ticks_i[2]
  PIN temp1_ticks_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.240 300.000 163.840 ;
    END
  END temp1_ticks_i[3]
  PIN temp1_ticks_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.320 300.000 167.920 ;
    END
  END temp1_ticks_i[4]
  PIN temp1_ticks_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.400 300.000 172.000 ;
    END
  END temp1_ticks_i[5]
  PIN temp1_ticks_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 175.480 300.000 176.080 ;
    END
  END temp1_ticks_i[6]
  PIN temp1_ticks_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.560 300.000 180.160 ;
    END
  END temp1_ticks_i[7]
  PIN temp1_ticks_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 183.640 300.000 184.240 ;
    END
  END temp1_ticks_i[8]
  PIN temp1_ticks_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.720 300.000 188.320 ;
    END
  END temp1_ticks_i[9]
  PIN temp2_dac_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 53.080 300.000 53.680 ;
    END
  END temp2_dac_i[0]
  PIN temp2_dac_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.160 300.000 57.760 ;
    END
  END temp2_dac_i[1]
  PIN temp2_dac_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 61.240 300.000 61.840 ;
    END
  END temp2_dac_i[2]
  PIN temp2_dac_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.320 300.000 65.920 ;
    END
  END temp2_dac_i[3]
  PIN temp2_dac_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 69.400 300.000 70.000 ;
    END
  END temp2_dac_i[4]
  PIN temp2_dac_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.480 300.000 74.080 ;
    END
  END temp2_dac_i[5]
  PIN temp2_ticks_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 199.960 300.000 200.560 ;
    END
  END temp2_ticks_i[0]
  PIN temp2_ticks_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.760 300.000 241.360 ;
    END
  END temp2_ticks_i[10]
  PIN temp2_ticks_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.840 300.000 245.440 ;
    END
  END temp2_ticks_i[11]
  PIN temp2_ticks_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 204.040 300.000 204.640 ;
    END
  END temp2_ticks_i[1]
  PIN temp2_ticks_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.120 300.000 208.720 ;
    END
  END temp2_ticks_i[2]
  PIN temp2_ticks_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 212.200 300.000 212.800 ;
    END
  END temp2_ticks_i[3]
  PIN temp2_ticks_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.280 300.000 216.880 ;
    END
  END temp2_ticks_i[4]
  PIN temp2_ticks_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.360 300.000 220.960 ;
    END
  END temp2_ticks_i[5]
  PIN temp2_ticks_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.440 300.000 225.040 ;
    END
  END temp2_ticks_i[6]
  PIN temp2_ticks_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.520 300.000 229.120 ;
    END
  END temp2_ticks_i[7]
  PIN temp2_ticks_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.600 300.000 233.200 ;
    END
  END temp2_ticks_i[8]
  PIN temp2_ticks_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.680 300.000 237.280 ;
    END
  END temp2_ticks_i[9]
  PIN temp3_dac_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 77.560 300.000 78.160 ;
    END
  END temp3_dac_i[0]
  PIN temp3_dac_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.640 300.000 82.240 ;
    END
  END temp3_dac_i[1]
  PIN temp3_dac_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 85.720 300.000 86.320 ;
    END
  END temp3_dac_i[2]
  PIN temp3_dac_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.800 300.000 90.400 ;
    END
  END temp3_dac_i[3]
  PIN temp3_dac_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 93.880 300.000 94.480 ;
    END
  END temp3_dac_i[4]
  PIN temp3_dac_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.960 300.000 98.560 ;
    END
  END temp3_dac_i[5]
  PIN temp3_ticks_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.920 300.000 249.520 ;
    END
  END temp3_ticks_i[0]
  PIN temp3_ticks_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.720 300.000 290.320 ;
    END
  END temp3_ticks_i[10]
  PIN temp3_ticks_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 293.800 300.000 294.400 ;
    END
  END temp3_ticks_i[11]
  PIN temp3_ticks_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 253.000 300.000 253.600 ;
    END
  END temp3_ticks_i[1]
  PIN temp3_ticks_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 257.080 300.000 257.680 ;
    END
  END temp3_ticks_i[2]
  PIN temp3_ticks_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.160 300.000 261.760 ;
    END
  END temp3_ticks_i[3]
  PIN temp3_ticks_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 265.240 300.000 265.840 ;
    END
  END temp3_ticks_i[4]
  PIN temp3_ticks_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 269.320 300.000 269.920 ;
    END
  END temp3_ticks_i[5]
  PIN temp3_ticks_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.400 300.000 274.000 ;
    END
  END temp3_ticks_i[6]
  PIN temp3_ticks_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.480 300.000 278.080 ;
    END
  END temp3_ticks_i[7]
  PIN temp3_ticks_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.560 300.000 282.160 ;
    END
  END temp3_ticks_i[8]
  PIN temp3_ticks_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 285.640 300.000 286.240 ;
    END
  END temp3_ticks_i[9]
  PIN temp_dac_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END temp_dac_o[0]
  PIN temp_dac_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END temp_dac_o[1]
  PIN temp_dac_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END temp_dac_o[2]
  PIN temp_dac_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END temp_dac_o[3]
  PIN temp_dac_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END temp_dac_o[4]
  PIN temp_dac_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END temp_dac_o[5]
  PIN temp_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END temp_sel_i[0]
  PIN temp_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END temp_sel_i[1]
  PIN temp_ticks_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END temp_ticks_o[0]
  PIN temp_ticks_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END temp_ticks_o[10]
  PIN temp_ticks_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END temp_ticks_o[11]
  PIN temp_ticks_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END temp_ticks_o[1]
  PIN temp_ticks_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END temp_ticks_o[2]
  PIN temp_ticks_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END temp_ticks_o[3]
  PIN temp_ticks_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END temp_ticks_o[4]
  PIN temp_ticks_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END temp_ticks_o[5]
  PIN temp_ticks_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END temp_ticks_o[6]
  PIN temp_ticks_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END temp_ticks_o[7]
  PIN temp_ticks_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END temp_ticks_o[8]
  PIN temp_ticks_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END temp_ticks_o[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 4.670 9.900 299.850 289.300 ;
      LAYER met2 ;
        RECT 4.690 295.720 9.010 296.000 ;
        RECT 9.850 295.720 14.990 296.000 ;
        RECT 15.830 295.720 20.970 296.000 ;
        RECT 21.810 295.720 26.950 296.000 ;
        RECT 27.790 295.720 32.930 296.000 ;
        RECT 33.770 295.720 38.910 296.000 ;
        RECT 39.750 295.720 44.890 296.000 ;
        RECT 45.730 295.720 50.870 296.000 ;
        RECT 51.710 295.720 56.850 296.000 ;
        RECT 57.690 295.720 62.830 296.000 ;
        RECT 63.670 295.720 68.810 296.000 ;
        RECT 69.650 295.720 74.790 296.000 ;
        RECT 75.630 295.720 80.770 296.000 ;
        RECT 81.610 295.720 86.750 296.000 ;
        RECT 87.590 295.720 92.730 296.000 ;
        RECT 93.570 295.720 98.710 296.000 ;
        RECT 99.550 295.720 104.690 296.000 ;
        RECT 105.530 295.720 110.670 296.000 ;
        RECT 111.510 295.720 116.650 296.000 ;
        RECT 117.490 295.720 122.630 296.000 ;
        RECT 123.470 295.720 128.610 296.000 ;
        RECT 129.450 295.720 134.590 296.000 ;
        RECT 135.430 295.720 140.570 296.000 ;
        RECT 141.410 295.720 146.550 296.000 ;
        RECT 147.390 295.720 152.530 296.000 ;
        RECT 153.370 295.720 158.510 296.000 ;
        RECT 159.350 295.720 164.490 296.000 ;
        RECT 165.330 295.720 170.470 296.000 ;
        RECT 171.310 295.720 176.450 296.000 ;
        RECT 177.290 295.720 182.430 296.000 ;
        RECT 183.270 295.720 188.410 296.000 ;
        RECT 189.250 295.720 194.390 296.000 ;
        RECT 195.230 295.720 200.370 296.000 ;
        RECT 201.210 295.720 206.350 296.000 ;
        RECT 207.190 295.720 212.330 296.000 ;
        RECT 213.170 295.720 218.310 296.000 ;
        RECT 219.150 295.720 224.290 296.000 ;
        RECT 225.130 295.720 230.270 296.000 ;
        RECT 231.110 295.720 236.250 296.000 ;
        RECT 237.090 295.720 242.230 296.000 ;
        RECT 243.070 295.720 248.210 296.000 ;
        RECT 249.050 295.720 254.190 296.000 ;
        RECT 255.030 295.720 260.170 296.000 ;
        RECT 261.010 295.720 266.150 296.000 ;
        RECT 266.990 295.720 272.130 296.000 ;
        RECT 272.970 295.720 278.110 296.000 ;
        RECT 278.950 295.720 284.090 296.000 ;
        RECT 284.930 295.720 290.070 296.000 ;
        RECT 290.910 295.720 299.820 296.000 ;
        RECT 4.690 4.280 299.820 295.720 ;
        RECT 4.690 3.670 11.310 4.280 ;
        RECT 12.150 3.670 16.830 4.280 ;
        RECT 17.670 3.670 22.350 4.280 ;
        RECT 23.190 3.670 27.870 4.280 ;
        RECT 28.710 3.670 33.390 4.280 ;
        RECT 34.230 3.670 38.910 4.280 ;
        RECT 39.750 3.670 44.430 4.280 ;
        RECT 45.270 3.670 49.950 4.280 ;
        RECT 50.790 3.670 55.470 4.280 ;
        RECT 56.310 3.670 60.990 4.280 ;
        RECT 61.830 3.670 66.510 4.280 ;
        RECT 67.350 3.670 72.030 4.280 ;
        RECT 72.870 3.670 77.550 4.280 ;
        RECT 78.390 3.670 83.070 4.280 ;
        RECT 83.910 3.670 88.590 4.280 ;
        RECT 89.430 3.670 94.110 4.280 ;
        RECT 94.950 3.670 99.630 4.280 ;
        RECT 100.470 3.670 105.150 4.280 ;
        RECT 105.990 3.670 110.670 4.280 ;
        RECT 111.510 3.670 116.190 4.280 ;
        RECT 117.030 3.670 121.710 4.280 ;
        RECT 122.550 3.670 127.230 4.280 ;
        RECT 128.070 3.670 132.750 4.280 ;
        RECT 133.590 3.670 138.270 4.280 ;
        RECT 139.110 3.670 143.790 4.280 ;
        RECT 144.630 3.670 149.310 4.280 ;
        RECT 150.150 3.670 154.830 4.280 ;
        RECT 155.670 3.670 160.350 4.280 ;
        RECT 161.190 3.670 165.870 4.280 ;
        RECT 166.710 3.670 171.390 4.280 ;
        RECT 172.230 3.670 176.910 4.280 ;
        RECT 177.750 3.670 182.430 4.280 ;
        RECT 183.270 3.670 187.950 4.280 ;
        RECT 188.790 3.670 193.470 4.280 ;
        RECT 194.310 3.670 198.990 4.280 ;
        RECT 199.830 3.670 204.510 4.280 ;
        RECT 205.350 3.670 210.030 4.280 ;
        RECT 210.870 3.670 215.550 4.280 ;
        RECT 216.390 3.670 221.070 4.280 ;
        RECT 221.910 3.670 226.590 4.280 ;
        RECT 227.430 3.670 232.110 4.280 ;
        RECT 232.950 3.670 237.630 4.280 ;
        RECT 238.470 3.670 243.150 4.280 ;
        RECT 243.990 3.670 248.670 4.280 ;
        RECT 249.510 3.670 254.190 4.280 ;
        RECT 255.030 3.670 259.710 4.280 ;
        RECT 260.550 3.670 265.230 4.280 ;
        RECT 266.070 3.670 270.750 4.280 ;
        RECT 271.590 3.670 276.270 4.280 ;
        RECT 277.110 3.670 281.790 4.280 ;
        RECT 282.630 3.670 287.310 4.280 ;
        RECT 288.150 3.670 299.820 4.280 ;
      LAYER met3 ;
        RECT 3.990 293.400 295.600 294.265 ;
        RECT 3.990 290.720 296.000 293.400 ;
        RECT 3.990 289.320 295.600 290.720 ;
        RECT 3.990 286.640 296.000 289.320 ;
        RECT 3.990 285.240 295.600 286.640 ;
        RECT 3.990 282.560 296.000 285.240 ;
        RECT 3.990 281.160 295.600 282.560 ;
        RECT 3.990 278.480 296.000 281.160 ;
        RECT 4.400 277.080 295.600 278.480 ;
        RECT 3.990 274.400 296.000 277.080 ;
        RECT 4.400 273.000 295.600 274.400 ;
        RECT 3.990 270.320 296.000 273.000 ;
        RECT 4.400 268.920 295.600 270.320 ;
        RECT 3.990 266.240 296.000 268.920 ;
        RECT 4.400 264.840 295.600 266.240 ;
        RECT 3.990 262.160 296.000 264.840 ;
        RECT 4.400 260.760 295.600 262.160 ;
        RECT 3.990 258.080 296.000 260.760 ;
        RECT 4.400 256.680 295.600 258.080 ;
        RECT 3.990 254.000 296.000 256.680 ;
        RECT 4.400 252.600 295.600 254.000 ;
        RECT 3.990 249.920 296.000 252.600 ;
        RECT 4.400 248.520 295.600 249.920 ;
        RECT 3.990 245.840 296.000 248.520 ;
        RECT 4.400 244.440 295.600 245.840 ;
        RECT 3.990 241.760 296.000 244.440 ;
        RECT 4.400 240.360 295.600 241.760 ;
        RECT 3.990 237.680 296.000 240.360 ;
        RECT 4.400 236.280 295.600 237.680 ;
        RECT 3.990 233.600 296.000 236.280 ;
        RECT 4.400 232.200 295.600 233.600 ;
        RECT 3.990 229.520 296.000 232.200 ;
        RECT 4.400 228.120 295.600 229.520 ;
        RECT 3.990 225.440 296.000 228.120 ;
        RECT 4.400 224.040 295.600 225.440 ;
        RECT 3.990 221.360 296.000 224.040 ;
        RECT 4.400 219.960 295.600 221.360 ;
        RECT 3.990 217.280 296.000 219.960 ;
        RECT 4.400 215.880 295.600 217.280 ;
        RECT 3.990 213.200 296.000 215.880 ;
        RECT 4.400 211.800 295.600 213.200 ;
        RECT 3.990 209.120 296.000 211.800 ;
        RECT 4.400 207.720 295.600 209.120 ;
        RECT 3.990 205.040 296.000 207.720 ;
        RECT 4.400 203.640 295.600 205.040 ;
        RECT 3.990 200.960 296.000 203.640 ;
        RECT 4.400 199.560 295.600 200.960 ;
        RECT 3.990 196.880 296.000 199.560 ;
        RECT 4.400 195.480 295.600 196.880 ;
        RECT 3.990 192.800 296.000 195.480 ;
        RECT 4.400 191.400 295.600 192.800 ;
        RECT 3.990 188.720 296.000 191.400 ;
        RECT 4.400 187.320 295.600 188.720 ;
        RECT 3.990 184.640 296.000 187.320 ;
        RECT 4.400 183.240 295.600 184.640 ;
        RECT 3.990 180.560 296.000 183.240 ;
        RECT 4.400 179.160 295.600 180.560 ;
        RECT 3.990 176.480 296.000 179.160 ;
        RECT 4.400 175.080 295.600 176.480 ;
        RECT 3.990 172.400 296.000 175.080 ;
        RECT 4.400 171.000 295.600 172.400 ;
        RECT 3.990 168.320 296.000 171.000 ;
        RECT 4.400 166.920 295.600 168.320 ;
        RECT 3.990 164.240 296.000 166.920 ;
        RECT 4.400 162.840 295.600 164.240 ;
        RECT 3.990 160.160 296.000 162.840 ;
        RECT 4.400 158.760 295.600 160.160 ;
        RECT 3.990 156.080 296.000 158.760 ;
        RECT 4.400 154.680 295.600 156.080 ;
        RECT 3.990 152.000 296.000 154.680 ;
        RECT 4.400 150.600 295.600 152.000 ;
        RECT 3.990 147.920 296.000 150.600 ;
        RECT 4.400 146.520 295.600 147.920 ;
        RECT 3.990 143.840 296.000 146.520 ;
        RECT 4.400 142.440 295.600 143.840 ;
        RECT 3.990 139.760 296.000 142.440 ;
        RECT 4.400 138.360 295.600 139.760 ;
        RECT 3.990 135.680 296.000 138.360 ;
        RECT 4.400 134.280 295.600 135.680 ;
        RECT 3.990 131.600 296.000 134.280 ;
        RECT 4.400 130.200 295.600 131.600 ;
        RECT 3.990 127.520 296.000 130.200 ;
        RECT 4.400 126.120 295.600 127.520 ;
        RECT 3.990 123.440 296.000 126.120 ;
        RECT 4.400 122.040 295.600 123.440 ;
        RECT 3.990 119.360 296.000 122.040 ;
        RECT 4.400 117.960 295.600 119.360 ;
        RECT 3.990 115.280 296.000 117.960 ;
        RECT 4.400 113.880 295.600 115.280 ;
        RECT 3.990 111.200 296.000 113.880 ;
        RECT 4.400 109.800 295.600 111.200 ;
        RECT 3.990 107.120 296.000 109.800 ;
        RECT 4.400 105.720 295.600 107.120 ;
        RECT 3.990 103.040 296.000 105.720 ;
        RECT 4.400 101.640 295.600 103.040 ;
        RECT 3.990 98.960 296.000 101.640 ;
        RECT 4.400 97.560 295.600 98.960 ;
        RECT 3.990 94.880 296.000 97.560 ;
        RECT 4.400 93.480 295.600 94.880 ;
        RECT 3.990 90.800 296.000 93.480 ;
        RECT 4.400 89.400 295.600 90.800 ;
        RECT 3.990 86.720 296.000 89.400 ;
        RECT 4.400 85.320 295.600 86.720 ;
        RECT 3.990 82.640 296.000 85.320 ;
        RECT 4.400 81.240 295.600 82.640 ;
        RECT 3.990 78.560 296.000 81.240 ;
        RECT 4.400 77.160 295.600 78.560 ;
        RECT 3.990 74.480 296.000 77.160 ;
        RECT 4.400 73.080 295.600 74.480 ;
        RECT 3.990 70.400 296.000 73.080 ;
        RECT 4.400 69.000 295.600 70.400 ;
        RECT 3.990 66.320 296.000 69.000 ;
        RECT 4.400 64.920 295.600 66.320 ;
        RECT 3.990 62.240 296.000 64.920 ;
        RECT 4.400 60.840 295.600 62.240 ;
        RECT 3.990 58.160 296.000 60.840 ;
        RECT 4.400 56.760 295.600 58.160 ;
        RECT 3.990 54.080 296.000 56.760 ;
        RECT 4.400 52.680 295.600 54.080 ;
        RECT 3.990 50.000 296.000 52.680 ;
        RECT 4.400 48.600 295.600 50.000 ;
        RECT 3.990 45.920 296.000 48.600 ;
        RECT 4.400 44.520 295.600 45.920 ;
        RECT 3.990 41.840 296.000 44.520 ;
        RECT 4.400 40.440 295.600 41.840 ;
        RECT 3.990 37.760 296.000 40.440 ;
        RECT 4.400 36.360 295.600 37.760 ;
        RECT 3.990 33.680 296.000 36.360 ;
        RECT 4.400 32.280 295.600 33.680 ;
        RECT 3.990 29.600 296.000 32.280 ;
        RECT 4.400 28.200 295.600 29.600 ;
        RECT 3.990 25.520 296.000 28.200 ;
        RECT 4.400 24.120 295.600 25.520 ;
        RECT 3.990 21.440 296.000 24.120 ;
        RECT 4.400 20.040 295.600 21.440 ;
        RECT 3.990 17.360 296.000 20.040 ;
        RECT 3.990 15.960 295.600 17.360 ;
        RECT 3.990 13.280 296.000 15.960 ;
        RECT 3.990 11.880 295.600 13.280 ;
        RECT 3.990 9.200 296.000 11.880 ;
        RECT 3.990 7.800 295.600 9.200 ;
        RECT 3.990 5.120 296.000 7.800 ;
        RECT 3.990 4.255 295.600 5.120 ;
      LAYER met4 ;
        RECT 282.735 19.215 284.905 200.425 ;
  END
END config_reg_mux
END LIBRARY

