magic
tech sky130A
magscale 1 2
timestamp 1671811341
<< viali >>
rect 28365 27557 28399 27591
rect 1777 27421 1811 27455
rect 28181 27421 28215 27455
rect 1593 27285 1627 27319
rect 28365 26469 28399 26503
rect 28181 26333 28215 26367
rect 28181 23681 28215 23715
rect 28365 23477 28399 23511
rect 23581 22729 23615 22763
rect 23673 22661 23707 22695
rect 1777 22593 1811 22627
rect 25881 22593 25915 22627
rect 23489 22525 23523 22559
rect 1593 22389 1627 22423
rect 24041 22389 24075 22423
rect 25697 22389 25731 22423
rect 22648 22185 22682 22219
rect 24133 22185 24167 22219
rect 25592 22185 25626 22219
rect 22385 22049 22419 22083
rect 27077 22049 27111 22083
rect 27813 22049 27847 22083
rect 27905 22049 27939 22083
rect 20085 21981 20119 22015
rect 25329 21981 25363 22015
rect 20269 21845 20303 21879
rect 27353 21845 27387 21879
rect 27721 21845 27755 21879
rect 3617 21641 3651 21675
rect 23949 21641 23983 21675
rect 25973 21641 26007 21675
rect 26341 21641 26375 21675
rect 26433 21641 26467 21675
rect 19441 21573 19475 21607
rect 23397 21573 23431 21607
rect 19165 21505 19199 21539
rect 24133 21505 24167 21539
rect 27261 21505 27295 21539
rect 28181 21505 28215 21539
rect 1869 21437 1903 21471
rect 2145 21437 2179 21471
rect 23673 21437 23707 21471
rect 26617 21437 26651 21471
rect 20913 21301 20947 21335
rect 21925 21301 21959 21335
rect 27077 21301 27111 21335
rect 28365 21301 28399 21335
rect 3525 21097 3559 21131
rect 19993 21097 20027 21131
rect 22201 21097 22235 21131
rect 28089 21097 28123 21131
rect 1777 20961 1811 20995
rect 4353 20961 4387 20995
rect 4537 20961 4571 20995
rect 20453 20961 20487 20995
rect 20637 20961 20671 20995
rect 26617 20961 26651 20995
rect 16865 20893 16899 20927
rect 22017 20893 22051 20927
rect 26341 20893 26375 20927
rect 2053 20825 2087 20859
rect 4261 20825 4295 20859
rect 26065 20825 26099 20859
rect 3893 20757 3927 20791
rect 4905 20757 4939 20791
rect 17049 20757 17083 20791
rect 20361 20757 20395 20791
rect 2329 20553 2363 20587
rect 3249 20553 3283 20587
rect 21925 20553 21959 20587
rect 22385 20553 22419 20587
rect 27077 20553 27111 20587
rect 27537 20553 27571 20587
rect 18245 20485 18279 20519
rect 2513 20417 2547 20451
rect 3157 20417 3191 20451
rect 18521 20417 18555 20451
rect 22293 20417 22327 20451
rect 26709 20417 26743 20451
rect 27445 20417 27479 20451
rect 3433 20349 3467 20383
rect 22477 20349 22511 20383
rect 22937 20349 22971 20383
rect 27629 20349 27663 20383
rect 2789 20281 2823 20315
rect 3801 20213 3835 20247
rect 16773 20213 16807 20247
rect 26525 20213 26559 20247
rect 2421 20009 2455 20043
rect 16865 20009 16899 20043
rect 22017 20009 22051 20043
rect 27905 20009 27939 20043
rect 17325 19873 17359 19907
rect 17417 19873 17451 19907
rect 26157 19873 26191 19907
rect 26433 19873 26467 19907
rect 2605 19805 2639 19839
rect 21741 19805 21775 19839
rect 17233 19669 17267 19703
rect 19533 19465 19567 19499
rect 17785 19329 17819 19363
rect 23305 19329 23339 19363
rect 18061 19261 18095 19295
rect 23581 19261 23615 19295
rect 25053 19125 25087 19159
rect 6745 18921 6779 18955
rect 18245 18921 18279 18955
rect 23949 18921 23983 18955
rect 24501 18853 24535 18887
rect 21281 18785 21315 18819
rect 24961 18785 24995 18819
rect 25053 18785 25087 18819
rect 4997 18717 5031 18751
rect 18429 18717 18463 18751
rect 21097 18717 21131 18751
rect 24133 18717 24167 18751
rect 28181 18717 28215 18751
rect 5273 18649 5307 18683
rect 24869 18649 24903 18683
rect 20913 18581 20947 18615
rect 28365 18581 28399 18615
rect 2973 18377 3007 18411
rect 21557 18377 21591 18411
rect 24317 18377 24351 18411
rect 27077 18377 27111 18411
rect 7665 18309 7699 18343
rect 2237 18241 2271 18275
rect 19809 18241 19843 18275
rect 26709 18241 26743 18275
rect 27445 18241 27479 18275
rect 27537 18241 27571 18275
rect 4445 18173 4479 18207
rect 4721 18173 4755 18207
rect 7389 18173 7423 18207
rect 20085 18173 20119 18207
rect 27629 18173 27663 18207
rect 2421 18037 2455 18071
rect 5089 18037 5123 18071
rect 9137 18037 9171 18071
rect 26525 18037 26559 18071
rect 4077 17833 4111 17867
rect 5273 17833 5307 17867
rect 24685 17833 24719 17867
rect 28089 17833 28123 17867
rect 18153 17765 18187 17799
rect 20361 17765 20395 17799
rect 20913 17765 20947 17799
rect 2973 17697 3007 17731
rect 3249 17697 3283 17731
rect 21373 17697 21407 17731
rect 26617 17697 26651 17731
rect 4353 17629 4387 17663
rect 4442 17629 4476 17663
rect 4537 17629 4571 17663
rect 4721 17629 4755 17663
rect 5529 17629 5563 17663
rect 5641 17629 5675 17663
rect 5733 17629 5767 17663
rect 5917 17629 5951 17663
rect 6653 17629 6687 17663
rect 7665 17629 7699 17663
rect 8033 17629 8067 17663
rect 16497 17629 16531 17663
rect 17509 17629 17543 17663
rect 18245 17629 18279 17663
rect 19809 17629 19843 17663
rect 19993 17629 20027 17663
rect 21097 17629 21131 17663
rect 21189 17629 21223 17663
rect 21281 17629 21315 17663
rect 24501 17629 24535 17663
rect 26341 17629 26375 17663
rect 6469 17561 6503 17595
rect 7757 17561 7791 17595
rect 7849 17561 7883 17595
rect 20085 17561 20119 17595
rect 1501 17493 1535 17527
rect 6285 17493 6319 17527
rect 7481 17493 7515 17527
rect 16313 17493 16347 17527
rect 20177 17493 20211 17527
rect 1593 17289 1627 17323
rect 2237 17289 2271 17323
rect 18613 17289 18647 17323
rect 19533 17289 19567 17323
rect 21005 17289 21039 17323
rect 2697 17221 2731 17255
rect 5089 17221 5123 17255
rect 5273 17221 5307 17255
rect 7849 17221 7883 17255
rect 12817 17221 12851 17255
rect 17325 17221 17359 17255
rect 20453 17221 20487 17255
rect 20637 17221 20671 17255
rect 23765 17221 23799 17255
rect 1777 17153 1811 17187
rect 2605 17153 2639 17187
rect 14933 17153 14967 17187
rect 15945 17153 15979 17187
rect 16129 17153 16163 17187
rect 17141 17153 17175 17187
rect 18245 17153 18279 17187
rect 19809 17153 19843 17187
rect 19901 17153 19935 17187
rect 19993 17153 20027 17187
rect 20361 17153 20395 17187
rect 20913 17153 20947 17187
rect 21097 17153 21131 17187
rect 23489 17153 23523 17187
rect 2881 17085 2915 17119
rect 3341 17085 3375 17119
rect 7573 17085 7607 17119
rect 14565 17085 14599 17119
rect 15577 17085 15611 17119
rect 19717 17085 19751 17119
rect 23213 17085 23247 17119
rect 6009 17017 6043 17051
rect 15669 17017 15703 17051
rect 20637 17017 20671 17051
rect 5457 16949 5491 16983
rect 9321 16949 9355 16983
rect 10333 16949 10367 16983
rect 11621 16949 11655 16983
rect 13139 16949 13173 16983
rect 17509 16949 17543 16983
rect 18613 16949 18647 16983
rect 18797 16949 18831 16983
rect 25237 16949 25271 16983
rect 14197 16745 14231 16779
rect 17509 16745 17543 16779
rect 17693 16745 17727 16779
rect 24133 16745 24167 16779
rect 24501 16745 24535 16779
rect 10517 16609 10551 16643
rect 15209 16609 15243 16643
rect 15485 16609 15519 16643
rect 16957 16609 16991 16643
rect 21741 16609 21775 16643
rect 25053 16609 25087 16643
rect 7573 16541 7607 16575
rect 7941 16541 7975 16575
rect 9689 16541 9723 16575
rect 10057 16541 10091 16575
rect 14381 16541 14415 16575
rect 14657 16541 14691 16575
rect 14841 16541 14875 16575
rect 19349 16541 19383 16575
rect 28181 16541 28215 16575
rect 7665 16473 7699 16507
rect 7757 16473 7791 16507
rect 9873 16473 9907 16507
rect 9965 16473 9999 16507
rect 10793 16473 10827 16507
rect 17677 16473 17711 16507
rect 17877 16473 17911 16507
rect 18705 16473 18739 16507
rect 22017 16473 22051 16507
rect 24961 16473 24995 16507
rect 7389 16405 7423 16439
rect 10241 16405 10275 16439
rect 12265 16405 12299 16439
rect 18429 16405 18463 16439
rect 19533 16405 19567 16439
rect 23489 16405 23523 16439
rect 24869 16405 24903 16439
rect 28365 16405 28399 16439
rect 22109 16201 22143 16235
rect 25237 16201 25271 16235
rect 27537 16201 27571 16235
rect 4629 16133 4663 16167
rect 7941 16133 7975 16167
rect 9137 16133 9171 16167
rect 15393 16133 15427 16167
rect 3985 16065 4019 16099
rect 4077 16065 4111 16099
rect 4169 16065 4203 16099
rect 4353 16065 4387 16099
rect 4813 16065 4847 16099
rect 7733 16065 7767 16099
rect 7841 16065 7875 16099
rect 8125 16065 8159 16099
rect 9413 16065 9447 16099
rect 10057 16065 10091 16099
rect 15209 16065 15243 16099
rect 21925 16065 21959 16099
rect 25053 16065 25087 16099
rect 26525 16065 26559 16099
rect 27629 16065 27663 16099
rect 9229 15997 9263 16031
rect 10425 15997 10459 16031
rect 11621 15997 11655 16031
rect 11897 15997 11931 16031
rect 13369 15997 13403 16031
rect 27721 15997 27755 16031
rect 9597 15929 9631 15963
rect 10517 15929 10551 15963
rect 10977 15929 11011 15963
rect 27169 15929 27203 15963
rect 3709 15861 3743 15895
rect 4997 15861 5031 15895
rect 5273 15861 5307 15895
rect 7573 15861 7607 15895
rect 9137 15861 9171 15895
rect 10609 15861 10643 15895
rect 18061 15861 18095 15895
rect 26709 15861 26743 15895
rect 1777 15657 1811 15691
rect 3267 15657 3301 15691
rect 9137 15657 9171 15691
rect 11713 15657 11747 15691
rect 20361 15657 20395 15691
rect 20545 15657 20579 15691
rect 28365 15657 28399 15691
rect 19349 15589 19383 15623
rect 19993 15589 20027 15623
rect 24501 15589 24535 15623
rect 3525 15521 3559 15555
rect 5273 15521 5307 15555
rect 22569 15521 22603 15555
rect 26893 15521 26927 15555
rect 7021 15453 7055 15487
rect 7389 15453 7423 15487
rect 19533 15453 19567 15487
rect 19717 15453 19751 15487
rect 26249 15453 26283 15487
rect 26617 15453 26651 15487
rect 9413 15385 9447 15419
rect 10425 15385 10459 15419
rect 20821 15385 20855 15419
rect 25973 15385 26007 15419
rect 8677 15317 8711 15351
rect 12541 15317 12575 15351
rect 20361 15317 20395 15351
rect 18797 15113 18831 15147
rect 20729 15113 20763 15147
rect 21925 15113 21959 15147
rect 25053 15113 25087 15147
rect 25513 15113 25547 15147
rect 5641 15045 5675 15079
rect 7849 15045 7883 15079
rect 11897 15045 11931 15079
rect 18613 15045 18647 15079
rect 19165 15045 19199 15079
rect 22293 15045 22327 15079
rect 3157 14977 3191 15011
rect 5825 14977 5859 15011
rect 6837 14977 6871 15011
rect 7021 14977 7055 15011
rect 7573 14977 7607 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 12173 14977 12207 15011
rect 12449 14977 12483 15011
rect 18889 14977 18923 15011
rect 19349 14977 19383 15011
rect 19441 14977 19475 15011
rect 22109 14977 22143 15011
rect 22385 14977 22419 15011
rect 25145 14977 25179 15011
rect 3433 14909 3467 14943
rect 9321 14909 9355 14943
rect 12541 14909 12575 14943
rect 19165 14909 19199 14943
rect 24869 14909 24903 14943
rect 11621 14841 11655 14875
rect 17141 14841 17175 14875
rect 4905 14773 4939 14807
rect 6009 14773 6043 14807
rect 7205 14773 7239 14807
rect 12449 14773 12483 14807
rect 12817 14773 12851 14807
rect 18613 14773 18647 14807
rect 24409 14773 24443 14807
rect 3893 14569 3927 14603
rect 18337 14569 18371 14603
rect 21557 14569 21591 14603
rect 14933 14433 14967 14467
rect 17417 14433 17451 14467
rect 4149 14365 4183 14399
rect 4274 14359 4308 14393
rect 4374 14362 4408 14396
rect 4537 14365 4571 14399
rect 5181 14365 5215 14399
rect 6469 14365 6503 14399
rect 17233 14365 17267 14399
rect 18153 14365 18187 14399
rect 21741 14365 21775 14399
rect 21833 14365 21867 14399
rect 5365 14297 5399 14331
rect 6653 14297 6687 14331
rect 6837 14297 6871 14331
rect 15209 14297 15243 14331
rect 16957 14297 16991 14331
rect 17969 14297 18003 14331
rect 22109 14297 22143 14331
rect 4813 14229 4847 14263
rect 5549 14229 5583 14263
rect 21925 14229 21959 14263
rect 17417 14025 17451 14059
rect 21458 14025 21492 14059
rect 24225 14025 24259 14059
rect 6561 13957 6595 13991
rect 18429 13957 18463 13991
rect 21557 13957 21591 13991
rect 21925 13957 21959 13991
rect 22753 13957 22787 13991
rect 24961 13957 24995 13991
rect 12725 13889 12759 13923
rect 13093 13889 13127 13923
rect 13553 13889 13587 13923
rect 14105 13889 14139 13923
rect 15301 13889 15335 13923
rect 15393 13889 15427 13923
rect 15577 13889 15611 13923
rect 15669 13889 15703 13923
rect 17325 13889 17359 13923
rect 17509 13889 17543 13923
rect 20177 13889 20211 13923
rect 21281 13889 21315 13923
rect 21373 13889 21407 13923
rect 22201 13889 22235 13923
rect 24593 13889 24627 13923
rect 27261 13889 27295 13923
rect 28181 13889 28215 13923
rect 13921 13821 13955 13855
rect 18153 13821 18187 13855
rect 21925 13821 21959 13855
rect 22477 13821 22511 13855
rect 6745 13753 6779 13787
rect 15117 13753 15151 13787
rect 12541 13685 12575 13719
rect 22109 13685 22143 13719
rect 27077 13685 27111 13719
rect 28365 13685 28399 13719
rect 10793 13481 10827 13515
rect 11161 13481 11195 13515
rect 13737 13481 13771 13515
rect 14657 13481 14691 13515
rect 14841 13481 14875 13515
rect 15393 13481 15427 13515
rect 20545 13481 20579 13515
rect 22109 13481 22143 13515
rect 17417 13413 17451 13447
rect 13737 13345 13771 13379
rect 14289 13345 14323 13379
rect 16865 13345 16899 13379
rect 26893 13345 26927 13379
rect 2421 13277 2455 13311
rect 8677 13277 8711 13311
rect 9045 13277 9079 13311
rect 11161 13277 11195 13311
rect 11253 13277 11287 13311
rect 13369 13277 13403 13311
rect 14197 13277 14231 13311
rect 14381 13277 14415 13311
rect 15485 13277 15519 13311
rect 16681 13277 16715 13311
rect 20821 13277 20855 13311
rect 22845 13277 22879 13311
rect 24961 13277 24995 13311
rect 26617 13277 26651 13311
rect 4721 13209 4755 13243
rect 4905 13209 4939 13243
rect 9321 13209 9355 13243
rect 15025 13209 15059 13243
rect 15761 13209 15795 13243
rect 15945 13209 15979 13243
rect 17417 13209 17451 13243
rect 2237 13141 2271 13175
rect 5089 13141 5123 13175
rect 11529 13141 11563 13175
rect 13001 13141 13035 13175
rect 14825 13141 14859 13175
rect 16129 13141 16163 13175
rect 16957 13141 16991 13175
rect 23029 13141 23063 13175
rect 25145 13141 25179 13175
rect 28365 13141 28399 13175
rect 9597 12937 9631 12971
rect 10057 12937 10091 12971
rect 16773 12937 16807 12971
rect 20571 12937 20605 12971
rect 27261 12937 27295 12971
rect 27721 12937 27755 12971
rect 1777 12869 1811 12903
rect 5733 12869 5767 12903
rect 8309 12869 8343 12903
rect 10793 12869 10827 12903
rect 20361 12869 20395 12903
rect 21373 12869 21407 12903
rect 22077 12869 22111 12903
rect 22293 12869 22327 12903
rect 25881 12869 25915 12903
rect 27629 12869 27663 12903
rect 4077 12801 4111 12835
rect 4166 12804 4200 12838
rect 4282 12801 4316 12835
rect 4445 12801 4479 12835
rect 5549 12801 5583 12835
rect 5917 12801 5951 12835
rect 6837 12801 6871 12835
rect 7297 12801 7331 12835
rect 8493 12801 8527 12835
rect 9505 12801 9539 12835
rect 9689 12801 9723 12835
rect 9965 12801 9999 12835
rect 10251 12801 10285 12835
rect 10977 12801 11011 12835
rect 12265 12801 12299 12835
rect 14197 12801 14231 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 21189 12801 21223 12835
rect 21465 12801 21499 12835
rect 26157 12801 26191 12835
rect 1501 12733 1535 12767
rect 6745 12733 6779 12767
rect 15945 12733 15979 12767
rect 27813 12733 27847 12767
rect 10241 12665 10275 12699
rect 21005 12665 21039 12699
rect 21925 12665 21959 12699
rect 3249 12597 3283 12631
rect 3801 12597 3835 12631
rect 4813 12597 4847 12631
rect 6469 12597 6503 12631
rect 7389 12597 7423 12631
rect 8677 12597 8711 12631
rect 10609 12597 10643 12631
rect 12357 12597 12391 12631
rect 13829 12597 13863 12631
rect 16957 12597 16991 12631
rect 20545 12597 20579 12631
rect 20729 12597 20763 12631
rect 22109 12597 22143 12631
rect 24409 12597 24443 12631
rect 26709 12597 26743 12631
rect 1593 12393 1627 12427
rect 2237 12393 2271 12427
rect 15485 12393 15519 12427
rect 15669 12393 15703 12427
rect 25421 12393 25455 12427
rect 12357 12325 12391 12359
rect 2881 12257 2915 12291
rect 7021 12257 7055 12291
rect 7665 12257 7699 12291
rect 11621 12257 11655 12291
rect 12081 12257 12115 12291
rect 12725 12257 12759 12291
rect 13093 12257 13127 12291
rect 17601 12257 17635 12291
rect 17693 12257 17727 12291
rect 19993 12257 20027 12291
rect 21741 12257 21775 12291
rect 24777 12257 24811 12291
rect 24961 12257 24995 12291
rect 1777 12189 1811 12223
rect 2697 12189 2731 12223
rect 6193 12189 6227 12223
rect 6377 12189 6411 12223
rect 6653 12189 6687 12223
rect 7297 12189 7331 12223
rect 11713 12189 11747 12223
rect 13001 12189 13035 12223
rect 13185 12189 13219 12223
rect 16037 12189 16071 12223
rect 17509 12189 17543 12223
rect 25053 12189 25087 12223
rect 2605 12121 2639 12155
rect 6285 12121 6319 12155
rect 9873 12121 9907 12155
rect 15669 12121 15703 12155
rect 20269 12121 20303 12155
rect 3433 12053 3467 12087
rect 3893 12053 3927 12087
rect 5917 12053 5951 12087
rect 7021 12053 7055 12087
rect 7665 12053 7699 12087
rect 12357 12053 12391 12087
rect 13553 12053 13587 12087
rect 17325 12053 17359 12087
rect 24133 12053 24167 12087
rect 4537 11849 4571 11883
rect 17417 11849 17451 11883
rect 20545 11849 20579 11883
rect 3985 11781 4019 11815
rect 6837 11713 6871 11747
rect 7021 11713 7055 11747
rect 7297 11713 7331 11747
rect 12909 11713 12943 11747
rect 13093 11713 13127 11747
rect 13369 11713 13403 11747
rect 17785 11713 17819 11747
rect 20729 11713 20763 11747
rect 23489 11713 23523 11747
rect 27261 11713 27295 11747
rect 28181 11713 28215 11747
rect 4261 11645 4295 11679
rect 6653 11645 6687 11679
rect 7849 11645 7883 11679
rect 12725 11645 12759 11679
rect 17877 11645 17911 11679
rect 18061 11577 18095 11611
rect 2513 11509 2547 11543
rect 7481 11509 7515 11543
rect 13553 11509 13587 11543
rect 13921 11509 13955 11543
rect 18429 11509 18463 11543
rect 23673 11509 23707 11543
rect 27077 11509 27111 11543
rect 28365 11509 28399 11543
rect 7941 11305 7975 11339
rect 11345 11305 11379 11339
rect 13001 11305 13035 11339
rect 13737 11305 13771 11339
rect 7297 11169 7331 11203
rect 7573 11169 7607 11203
rect 9597 11169 9631 11203
rect 9873 11169 9907 11203
rect 13369 11169 13403 11203
rect 13737 11169 13771 11203
rect 22385 11169 22419 11203
rect 26801 11169 26835 11203
rect 4261 11101 4295 11135
rect 4629 11101 4663 11135
rect 6929 11101 6963 11135
rect 7941 11101 7975 11135
rect 8217 11101 8251 11135
rect 9505 11101 9539 11135
rect 10149 11101 10183 11135
rect 16037 11101 16071 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17233 11101 17267 11135
rect 17601 11101 17635 11135
rect 17785 11101 17819 11135
rect 24133 11101 24167 11135
rect 26525 11101 26559 11135
rect 6561 11033 6595 11067
rect 23857 11033 23891 11067
rect 4629 10965 4663 10999
rect 6929 10965 6963 10999
rect 10241 10965 10275 10999
rect 15393 10965 15427 10999
rect 17969 10965 18003 10999
rect 28273 10965 28307 10999
rect 4629 10761 4663 10795
rect 5273 10761 5307 10795
rect 9137 10761 9171 10795
rect 13185 10761 13219 10795
rect 23489 10761 23523 10795
rect 23949 10761 23983 10795
rect 27261 10761 27295 10795
rect 27629 10761 27663 10795
rect 27721 10761 27755 10795
rect 19257 10693 19291 10727
rect 20729 10693 20763 10727
rect 21005 10693 21039 10727
rect 4629 10625 4663 10659
rect 5273 10625 5307 10659
rect 5641 10625 5675 10659
rect 7849 10625 7883 10659
rect 9873 10625 9907 10659
rect 10425 10625 10459 10659
rect 11069 10625 11103 10659
rect 11253 10625 11287 10659
rect 11897 10625 11931 10659
rect 12817 10625 12851 10659
rect 13185 10625 13219 10659
rect 13461 10625 13495 10659
rect 15485 10625 15519 10659
rect 15669 10625 15703 10659
rect 16313 10625 16347 10659
rect 20453 10625 20487 10659
rect 20545 10625 20579 10659
rect 21281 10625 21315 10659
rect 23581 10625 23615 10659
rect 4261 10557 4295 10591
rect 4905 10557 4939 10591
rect 10793 10557 10827 10591
rect 11161 10557 11195 10591
rect 16221 10557 16255 10591
rect 17509 10557 17543 10591
rect 19533 10557 19567 10591
rect 21005 10557 21039 10591
rect 21189 10557 21223 10591
rect 22937 10557 22971 10591
rect 23397 10557 23431 10591
rect 27813 10557 27847 10591
rect 5641 10489 5675 10523
rect 12081 10489 12115 10523
rect 15669 10489 15703 10523
rect 10425 10421 10459 10455
rect 15945 10421 15979 10455
rect 16313 10421 16347 10455
rect 20729 10421 20763 10455
rect 26709 10421 26743 10455
rect 12541 10217 12575 10251
rect 13185 10217 13219 10251
rect 13829 10217 13863 10251
rect 14933 10217 14967 10251
rect 21833 10217 21867 10251
rect 4629 10149 4663 10183
rect 5273 10149 5307 10183
rect 9505 10149 9539 10183
rect 10149 10149 10183 10183
rect 4905 10081 4939 10115
rect 5917 10081 5951 10115
rect 6193 10081 6227 10115
rect 12173 10081 12207 10115
rect 15761 10081 15795 10115
rect 17785 10081 17819 10115
rect 20361 10081 20395 10115
rect 4261 10013 4295 10047
rect 5825 10013 5859 10047
rect 6653 10013 6687 10047
rect 6837 10013 6871 10047
rect 9137 10013 9171 10047
rect 9781 10013 9815 10047
rect 10425 10013 10459 10047
rect 12817 10013 12851 10047
rect 13185 10013 13219 10047
rect 13461 10013 13495 10047
rect 13829 10013 13863 10047
rect 15117 10013 15151 10047
rect 20085 10013 20119 10047
rect 6469 9945 6503 9979
rect 16037 9945 16071 9979
rect 4629 9877 4663 9911
rect 5273 9877 5307 9911
rect 7205 9877 7239 9911
rect 9505 9877 9539 9911
rect 10149 9877 10183 9911
rect 4629 9673 4663 9707
rect 5273 9673 5307 9707
rect 9137 9673 9171 9707
rect 12817 9673 12851 9707
rect 13461 9673 13495 9707
rect 11989 9605 12023 9639
rect 12265 9605 12299 9639
rect 17601 9605 17635 9639
rect 4629 9537 4663 9571
rect 5273 9537 5307 9571
rect 8309 9537 8343 9571
rect 8493 9537 8527 9571
rect 9781 9537 9815 9571
rect 10149 9537 10183 9571
rect 10701 9537 10735 9571
rect 11805 9537 11839 9571
rect 16957 9537 16991 9571
rect 17233 9537 17267 9571
rect 17785 9537 17819 9571
rect 24685 9537 24719 9571
rect 27261 9537 27295 9571
rect 28181 9537 28215 9571
rect 4261 9469 4295 9503
rect 4905 9469 4939 9503
rect 8401 9469 8435 9503
rect 8769 9469 8803 9503
rect 9505 9469 9539 9503
rect 10517 9469 10551 9503
rect 11161 9469 11195 9503
rect 11621 9469 11655 9503
rect 12817 9469 12851 9503
rect 13185 9469 13219 9503
rect 16773 9469 16807 9503
rect 17049 9469 17083 9503
rect 17141 9469 17175 9503
rect 9137 9401 9171 9435
rect 17969 9401 18003 9435
rect 9781 9333 9815 9367
rect 10885 9333 10919 9367
rect 24869 9333 24903 9367
rect 27077 9333 27111 9367
rect 28365 9333 28399 9367
rect 12265 9129 12299 9163
rect 12725 9129 12759 9163
rect 13001 9129 13035 9163
rect 13369 9129 13403 9163
rect 14197 9129 14231 9163
rect 4629 9061 4663 9095
rect 4261 8993 4295 9027
rect 9413 8993 9447 9027
rect 13369 8993 13403 9027
rect 14197 8993 14231 9027
rect 14841 8993 14875 9027
rect 25973 8993 26007 9027
rect 26801 8993 26835 9027
rect 7113 8925 7147 8959
rect 11805 8925 11839 8959
rect 13737 8925 13771 8959
rect 14565 8925 14599 8959
rect 21557 8925 21591 8959
rect 26249 8925 26283 8959
rect 26525 8925 26559 8959
rect 8125 8857 8159 8891
rect 11989 8857 12023 8891
rect 21833 8857 21867 8891
rect 4629 8789 4663 8823
rect 23305 8789 23339 8823
rect 24501 8789 24535 8823
rect 28273 8789 28307 8823
rect 2973 8585 3007 8619
rect 13093 8585 13127 8619
rect 13737 8585 13771 8619
rect 14381 8585 14415 8619
rect 15025 8585 15059 8619
rect 17969 8585 18003 8619
rect 21373 8585 21407 8619
rect 22477 8585 22511 8619
rect 24777 8585 24811 8619
rect 25237 8585 25271 8619
rect 27261 8585 27295 8619
rect 27629 8585 27663 8619
rect 27721 8585 27755 8619
rect 18245 8517 18279 8551
rect 21189 8517 21223 8551
rect 2329 8449 2363 8483
rect 3065 8449 3099 8483
rect 7205 8449 7239 8483
rect 7941 8449 7975 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 8861 8449 8895 8483
rect 12725 8449 12759 8483
rect 13369 8449 13403 8483
rect 14013 8449 14047 8483
rect 14657 8449 14691 8483
rect 20821 8449 20855 8483
rect 21925 8449 21959 8483
rect 22109 8449 22143 8483
rect 22661 8449 22695 8483
rect 24869 8449 24903 8483
rect 3157 8381 3191 8415
rect 3617 8381 3651 8415
rect 7665 8381 7699 8415
rect 9321 8381 9355 8415
rect 12449 8381 12483 8415
rect 13093 8381 13127 8415
rect 24225 8381 24259 8415
rect 24685 8381 24719 8415
rect 26709 8381 26743 8415
rect 27813 8381 27847 8415
rect 2605 8313 2639 8347
rect 13737 8313 13771 8347
rect 14381 8313 14415 8347
rect 15025 8313 15059 8347
rect 15301 8313 15335 8347
rect 2145 8245 2179 8279
rect 7113 8245 7147 8279
rect 9045 8245 9079 8279
rect 19533 8245 19567 8279
rect 21189 8245 21223 8279
rect 7021 8041 7055 8075
rect 7665 8041 7699 8075
rect 8585 8041 8619 8075
rect 12633 8041 12667 8075
rect 13001 8041 13035 8075
rect 13369 8041 13403 8075
rect 20453 8041 20487 8075
rect 23397 8041 23431 8075
rect 14197 7973 14231 8007
rect 14841 7973 14875 8007
rect 1685 7905 1719 7939
rect 1961 7905 1995 7939
rect 6653 7905 6687 7939
rect 7297 7905 7331 7939
rect 13369 7905 13403 7939
rect 13737 7905 13771 7939
rect 14565 7905 14599 7939
rect 7021 7837 7055 7871
rect 7665 7837 7699 7871
rect 9505 7837 9539 7871
rect 20821 7837 20855 7871
rect 23213 7837 23247 7871
rect 9873 7769 9907 7803
rect 22845 7769 22879 7803
rect 23121 7769 23155 7803
rect 3433 7701 3467 7735
rect 3893 7701 3927 7735
rect 14197 7701 14231 7735
rect 22293 7701 22327 7735
rect 23029 7701 23063 7735
rect 1593 7497 1627 7531
rect 6101 7497 6135 7531
rect 7021 7497 7055 7531
rect 7665 7497 7699 7531
rect 9873 7497 9907 7531
rect 10333 7497 10367 7531
rect 11069 7497 11103 7531
rect 13921 7497 13955 7531
rect 21925 7497 21959 7531
rect 1777 7361 1811 7395
rect 5733 7361 5767 7395
rect 6653 7361 6687 7395
rect 7297 7361 7331 7395
rect 11069 7361 11103 7395
rect 11621 7361 11655 7395
rect 22201 7361 22235 7395
rect 10701 7293 10735 7327
rect 19165 7293 19199 7327
rect 19533 7293 19567 7327
rect 22109 7293 22143 7327
rect 22293 7293 22327 7327
rect 22385 7293 22419 7327
rect 6101 7225 6135 7259
rect 7021 7225 7055 7259
rect 7665 7225 7699 7259
rect 17739 7157 17773 7191
rect 5733 6953 5767 6987
rect 6377 6953 6411 6987
rect 7021 6953 7055 6987
rect 7665 6953 7699 6987
rect 8309 6953 8343 6987
rect 9689 6953 9723 6987
rect 10425 6953 10459 6987
rect 11069 6953 11103 6987
rect 11713 6953 11747 6987
rect 12357 6953 12391 6987
rect 12633 6953 12667 6987
rect 18613 6953 18647 6987
rect 21005 6953 21039 6987
rect 5365 6817 5399 6851
rect 6009 6817 6043 6851
rect 6653 6817 6687 6851
rect 7297 6817 7331 6851
rect 7941 6817 7975 6851
rect 10057 6817 10091 6851
rect 10701 6817 10735 6851
rect 11345 6817 11379 6851
rect 11989 6817 12023 6851
rect 12357 6817 12391 6851
rect 22385 6817 22419 6851
rect 5733 6749 5767 6783
rect 6377 6749 6411 6783
rect 7021 6749 7055 6783
rect 7665 6749 7699 6783
rect 8309 6749 8343 6783
rect 10425 6749 10459 6783
rect 11069 6749 11103 6783
rect 11713 6749 11747 6783
rect 18337 6749 18371 6783
rect 18613 6749 18647 6783
rect 21649 6749 21683 6783
rect 21925 6749 21959 6783
rect 25237 6749 25271 6783
rect 27261 6749 27295 6783
rect 28181 6749 28215 6783
rect 18521 6681 18555 6715
rect 20821 6681 20855 6715
rect 21037 6681 21071 6715
rect 21465 6681 21499 6715
rect 21833 6681 21867 6715
rect 22661 6681 22695 6715
rect 18889 6613 18923 6647
rect 21189 6613 21223 6647
rect 24133 6613 24167 6647
rect 25421 6613 25455 6647
rect 27077 6613 27111 6647
rect 27629 6613 27663 6647
rect 28365 6613 28399 6647
rect 4077 6409 4111 6443
rect 5273 6409 5307 6443
rect 6101 6409 6135 6443
rect 7021 6409 7055 6443
rect 7665 6409 7699 6443
rect 8309 6409 8343 6443
rect 9045 6409 9079 6443
rect 9413 6409 9447 6443
rect 21097 6409 21131 6443
rect 22385 6409 22419 6443
rect 27261 6409 27295 6443
rect 21189 6341 21223 6375
rect 21373 6341 21407 6375
rect 26249 6341 26283 6375
rect 27629 6341 27663 6375
rect 4077 6273 4111 6307
rect 5733 6273 5767 6307
rect 6653 6273 6687 6307
rect 7297 6273 7331 6307
rect 7941 6273 7975 6307
rect 8309 6273 8343 6307
rect 9413 6273 9447 6307
rect 9781 6273 9815 6307
rect 10057 6273 10091 6307
rect 10701 6273 10735 6307
rect 11621 6273 11655 6307
rect 12265 6273 12299 6307
rect 12633 6273 12667 6307
rect 19717 6273 19751 6307
rect 19809 6273 19843 6307
rect 21097 6273 21131 6307
rect 22201 6273 22235 6307
rect 4445 6205 4479 6239
rect 4721 6205 4755 6239
rect 10425 6205 10459 6239
rect 11069 6205 11103 6239
rect 11989 6205 12023 6239
rect 12909 6205 12943 6239
rect 13277 6205 13311 6239
rect 19533 6205 19567 6239
rect 26525 6205 26559 6239
rect 27721 6205 27755 6239
rect 27813 6205 27847 6239
rect 6101 6137 6135 6171
rect 7021 6137 7055 6171
rect 7665 6137 7699 6171
rect 10425 6069 10459 6103
rect 11069 6069 11103 6103
rect 11989 6069 12023 6103
rect 12633 6069 12667 6103
rect 13277 6069 13311 6103
rect 13553 6069 13587 6103
rect 19625 6069 19659 6103
rect 24777 6069 24811 6103
rect 9321 5865 9355 5899
rect 12357 5865 12391 5899
rect 12633 5865 12667 5899
rect 24685 5865 24719 5899
rect 25697 5865 25731 5899
rect 28365 5865 28399 5899
rect 6653 5797 6687 5831
rect 7297 5797 7331 5831
rect 11713 5797 11747 5831
rect 19349 5797 19383 5831
rect 7021 5729 7055 5763
rect 7665 5729 7699 5763
rect 10057 5729 10091 5763
rect 10701 5729 10735 5763
rect 11345 5729 11379 5763
rect 11989 5729 12023 5763
rect 12357 5729 12391 5763
rect 25053 5729 25087 5763
rect 25237 5729 25271 5763
rect 26893 5729 26927 5763
rect 10425 5661 10459 5695
rect 11069 5661 11103 5695
rect 19349 5661 19383 5695
rect 19625 5661 19659 5695
rect 25329 5661 25363 5695
rect 26617 5661 26651 5695
rect 9781 5593 9815 5627
rect 6653 5525 6687 5559
rect 7297 5525 7331 5559
rect 10425 5525 10459 5559
rect 11069 5525 11103 5559
rect 11713 5525 11747 5559
rect 19533 5525 19567 5559
rect 9965 5321 9999 5355
rect 10425 5321 10459 5355
rect 10701 5321 10735 5355
rect 11713 5321 11747 5355
rect 11989 5321 12023 5355
rect 20545 5321 20579 5355
rect 10701 5185 10735 5219
rect 11069 5185 11103 5219
rect 18797 5185 18831 5219
rect 19073 5117 19107 5151
rect 23029 4981 23063 5015
rect 10609 4777 10643 4811
rect 11161 4777 11195 4811
rect 21833 4641 21867 4675
rect 22753 4641 22787 4675
rect 23765 4641 23799 4675
rect 22477 4573 22511 4607
rect 23489 4573 23523 4607
rect 26709 4573 26743 4607
rect 26985 4505 27019 4539
rect 3341 4437 3375 4471
rect 22109 4437 22143 4471
rect 22569 4437 22603 4471
rect 23121 4437 23155 4471
rect 23581 4437 23615 4471
rect 28457 4437 28491 4471
rect 2881 4233 2915 4267
rect 27721 4233 27755 4267
rect 3893 4165 3927 4199
rect 22569 4165 22603 4199
rect 20545 4097 20579 4131
rect 22017 4097 22051 4131
rect 23213 4097 23247 4131
rect 25421 4097 25455 4131
rect 27629 4097 27663 4131
rect 2973 4029 3007 4063
rect 3157 4029 3191 4063
rect 26709 4029 26743 4063
rect 27813 4029 27847 4063
rect 22201 3961 22235 3995
rect 23397 3961 23431 3995
rect 2513 3893 2547 3927
rect 3801 3893 3835 3927
rect 20453 3893 20487 3927
rect 22845 3893 22879 3927
rect 25237 3893 25271 3927
rect 27261 3893 27295 3927
rect 3433 3689 3467 3723
rect 21097 3689 21131 3723
rect 23121 3689 23155 3723
rect 27077 3689 27111 3723
rect 28365 3689 28399 3723
rect 1685 3553 1719 3587
rect 18705 3553 18739 3587
rect 19349 3553 19383 3587
rect 21373 3553 21407 3587
rect 21649 3553 21683 3587
rect 24869 3553 24903 3587
rect 3893 3485 3927 3519
rect 18521 3485 18555 3519
rect 18797 3485 18831 3519
rect 18894 3485 18928 3519
rect 27261 3485 27295 3519
rect 28181 3485 28215 3519
rect 1961 3417 1995 3451
rect 18245 3417 18279 3451
rect 18705 3417 18739 3451
rect 19625 3417 19659 3451
rect 25145 3417 25179 3451
rect 26617 3349 26651 3383
rect 2237 3145 2271 3179
rect 2973 3145 3007 3179
rect 19717 3145 19751 3179
rect 24041 3145 24075 3179
rect 25421 3145 25455 3179
rect 25789 3145 25823 3179
rect 20085 3077 20119 3111
rect 20453 3077 20487 3111
rect 22569 3077 22603 3111
rect 1777 3009 1811 3043
rect 2421 3009 2455 3043
rect 3249 3009 3283 3043
rect 22293 3009 22327 3043
rect 25881 3009 25915 3043
rect 18429 2941 18463 2975
rect 25145 2941 25179 2975
rect 25973 2941 26007 2975
rect 3709 2873 3743 2907
rect 1593 2805 1627 2839
rect 11621 2601 11655 2635
rect 18797 2601 18831 2635
rect 11805 2397 11839 2431
rect 12081 2397 12115 2431
rect 18981 2397 19015 2431
rect 19349 2397 19383 2431
rect 26249 2397 26283 2431
rect 28181 2397 28215 2431
rect 26433 2261 26467 2295
rect 28365 2261 28399 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 3350 27770
rect 3402 27718 3414 27770
rect 3466 27718 3478 27770
rect 3530 27718 3542 27770
rect 3594 27718 3606 27770
rect 3658 27718 8150 27770
rect 8202 27718 8214 27770
rect 8266 27718 8278 27770
rect 8330 27718 8342 27770
rect 8394 27718 8406 27770
rect 8458 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 17750 27770
rect 17802 27718 17814 27770
rect 17866 27718 17878 27770
rect 17930 27718 17942 27770
rect 17994 27718 18006 27770
rect 18058 27718 22550 27770
rect 22602 27718 22614 27770
rect 22666 27718 22678 27770
rect 22730 27718 22742 27770
rect 22794 27718 22806 27770
rect 22858 27718 27350 27770
rect 27402 27718 27414 27770
rect 27466 27718 27478 27770
rect 27530 27718 27542 27770
rect 27594 27718 27606 27770
rect 27658 27718 28888 27770
rect 1104 27696 28888 27718
rect 28350 27588 28356 27600
rect 28311 27560 28356 27588
rect 28350 27548 28356 27560
rect 28408 27548 28414 27600
rect 1765 27455 1823 27461
rect 1765 27421 1777 27455
rect 1811 27452 1823 27455
rect 3050 27452 3056 27464
rect 1811 27424 3056 27452
rect 1811 27421 1823 27424
rect 1765 27415 1823 27421
rect 3050 27412 3056 27424
rect 3108 27412 3114 27464
rect 27798 27412 27804 27464
rect 27856 27452 27862 27464
rect 28169 27455 28227 27461
rect 28169 27452 28181 27455
rect 27856 27424 28181 27452
rect 27856 27412 27862 27424
rect 28169 27421 28181 27424
rect 28215 27421 28227 27455
rect 28169 27415 28227 27421
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 1104 27226 28888 27248
rect 1104 27174 5750 27226
rect 5802 27174 5814 27226
rect 5866 27174 5878 27226
rect 5930 27174 5942 27226
rect 5994 27174 6006 27226
rect 6058 27174 10550 27226
rect 10602 27174 10614 27226
rect 10666 27174 10678 27226
rect 10730 27174 10742 27226
rect 10794 27174 10806 27226
rect 10858 27174 15350 27226
rect 15402 27174 15414 27226
rect 15466 27174 15478 27226
rect 15530 27174 15542 27226
rect 15594 27174 15606 27226
rect 15658 27174 20150 27226
rect 20202 27174 20214 27226
rect 20266 27174 20278 27226
rect 20330 27174 20342 27226
rect 20394 27174 20406 27226
rect 20458 27174 24950 27226
rect 25002 27174 25014 27226
rect 25066 27174 25078 27226
rect 25130 27174 25142 27226
rect 25194 27174 25206 27226
rect 25258 27174 28888 27226
rect 1104 27152 28888 27174
rect 1104 26682 28888 26704
rect 1104 26630 3350 26682
rect 3402 26630 3414 26682
rect 3466 26630 3478 26682
rect 3530 26630 3542 26682
rect 3594 26630 3606 26682
rect 3658 26630 8150 26682
rect 8202 26630 8214 26682
rect 8266 26630 8278 26682
rect 8330 26630 8342 26682
rect 8394 26630 8406 26682
rect 8458 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 17750 26682
rect 17802 26630 17814 26682
rect 17866 26630 17878 26682
rect 17930 26630 17942 26682
rect 17994 26630 18006 26682
rect 18058 26630 22550 26682
rect 22602 26630 22614 26682
rect 22666 26630 22678 26682
rect 22730 26630 22742 26682
rect 22794 26630 22806 26682
rect 22858 26630 27350 26682
rect 27402 26630 27414 26682
rect 27466 26630 27478 26682
rect 27530 26630 27542 26682
rect 27594 26630 27606 26682
rect 27658 26630 28888 26682
rect 1104 26608 28888 26630
rect 28350 26500 28356 26512
rect 28311 26472 28356 26500
rect 28350 26460 28356 26472
rect 28408 26460 28414 26512
rect 27706 26324 27712 26376
rect 27764 26364 27770 26376
rect 28169 26367 28227 26373
rect 28169 26364 28181 26367
rect 27764 26336 28181 26364
rect 27764 26324 27770 26336
rect 28169 26333 28181 26336
rect 28215 26333 28227 26367
rect 28169 26327 28227 26333
rect 1104 26138 28888 26160
rect 1104 26086 5750 26138
rect 5802 26086 5814 26138
rect 5866 26086 5878 26138
rect 5930 26086 5942 26138
rect 5994 26086 6006 26138
rect 6058 26086 10550 26138
rect 10602 26086 10614 26138
rect 10666 26086 10678 26138
rect 10730 26086 10742 26138
rect 10794 26086 10806 26138
rect 10858 26086 15350 26138
rect 15402 26086 15414 26138
rect 15466 26086 15478 26138
rect 15530 26086 15542 26138
rect 15594 26086 15606 26138
rect 15658 26086 20150 26138
rect 20202 26086 20214 26138
rect 20266 26086 20278 26138
rect 20330 26086 20342 26138
rect 20394 26086 20406 26138
rect 20458 26086 24950 26138
rect 25002 26086 25014 26138
rect 25066 26086 25078 26138
rect 25130 26086 25142 26138
rect 25194 26086 25206 26138
rect 25258 26086 28888 26138
rect 1104 26064 28888 26086
rect 1104 25594 28888 25616
rect 1104 25542 3350 25594
rect 3402 25542 3414 25594
rect 3466 25542 3478 25594
rect 3530 25542 3542 25594
rect 3594 25542 3606 25594
rect 3658 25542 8150 25594
rect 8202 25542 8214 25594
rect 8266 25542 8278 25594
rect 8330 25542 8342 25594
rect 8394 25542 8406 25594
rect 8458 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 17750 25594
rect 17802 25542 17814 25594
rect 17866 25542 17878 25594
rect 17930 25542 17942 25594
rect 17994 25542 18006 25594
rect 18058 25542 22550 25594
rect 22602 25542 22614 25594
rect 22666 25542 22678 25594
rect 22730 25542 22742 25594
rect 22794 25542 22806 25594
rect 22858 25542 27350 25594
rect 27402 25542 27414 25594
rect 27466 25542 27478 25594
rect 27530 25542 27542 25594
rect 27594 25542 27606 25594
rect 27658 25542 28888 25594
rect 1104 25520 28888 25542
rect 1104 25050 28888 25072
rect 1104 24998 5750 25050
rect 5802 24998 5814 25050
rect 5866 24998 5878 25050
rect 5930 24998 5942 25050
rect 5994 24998 6006 25050
rect 6058 24998 10550 25050
rect 10602 24998 10614 25050
rect 10666 24998 10678 25050
rect 10730 24998 10742 25050
rect 10794 24998 10806 25050
rect 10858 24998 15350 25050
rect 15402 24998 15414 25050
rect 15466 24998 15478 25050
rect 15530 24998 15542 25050
rect 15594 24998 15606 25050
rect 15658 24998 20150 25050
rect 20202 24998 20214 25050
rect 20266 24998 20278 25050
rect 20330 24998 20342 25050
rect 20394 24998 20406 25050
rect 20458 24998 24950 25050
rect 25002 24998 25014 25050
rect 25066 24998 25078 25050
rect 25130 24998 25142 25050
rect 25194 24998 25206 25050
rect 25258 24998 28888 25050
rect 1104 24976 28888 24998
rect 1104 24506 28888 24528
rect 1104 24454 3350 24506
rect 3402 24454 3414 24506
rect 3466 24454 3478 24506
rect 3530 24454 3542 24506
rect 3594 24454 3606 24506
rect 3658 24454 8150 24506
rect 8202 24454 8214 24506
rect 8266 24454 8278 24506
rect 8330 24454 8342 24506
rect 8394 24454 8406 24506
rect 8458 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 17750 24506
rect 17802 24454 17814 24506
rect 17866 24454 17878 24506
rect 17930 24454 17942 24506
rect 17994 24454 18006 24506
rect 18058 24454 22550 24506
rect 22602 24454 22614 24506
rect 22666 24454 22678 24506
rect 22730 24454 22742 24506
rect 22794 24454 22806 24506
rect 22858 24454 27350 24506
rect 27402 24454 27414 24506
rect 27466 24454 27478 24506
rect 27530 24454 27542 24506
rect 27594 24454 27606 24506
rect 27658 24454 28888 24506
rect 1104 24432 28888 24454
rect 1104 23962 28888 23984
rect 1104 23910 5750 23962
rect 5802 23910 5814 23962
rect 5866 23910 5878 23962
rect 5930 23910 5942 23962
rect 5994 23910 6006 23962
rect 6058 23910 10550 23962
rect 10602 23910 10614 23962
rect 10666 23910 10678 23962
rect 10730 23910 10742 23962
rect 10794 23910 10806 23962
rect 10858 23910 15350 23962
rect 15402 23910 15414 23962
rect 15466 23910 15478 23962
rect 15530 23910 15542 23962
rect 15594 23910 15606 23962
rect 15658 23910 20150 23962
rect 20202 23910 20214 23962
rect 20266 23910 20278 23962
rect 20330 23910 20342 23962
rect 20394 23910 20406 23962
rect 20458 23910 24950 23962
rect 25002 23910 25014 23962
rect 25066 23910 25078 23962
rect 25130 23910 25142 23962
rect 25194 23910 25206 23962
rect 25258 23910 28888 23962
rect 1104 23888 28888 23910
rect 24210 23672 24216 23724
rect 24268 23712 24274 23724
rect 28169 23715 28227 23721
rect 28169 23712 28181 23715
rect 24268 23684 28181 23712
rect 24268 23672 24274 23684
rect 28169 23681 28181 23684
rect 28215 23681 28227 23715
rect 28169 23675 28227 23681
rect 28350 23508 28356 23520
rect 28311 23480 28356 23508
rect 28350 23468 28356 23480
rect 28408 23468 28414 23520
rect 1104 23418 28888 23440
rect 1104 23366 3350 23418
rect 3402 23366 3414 23418
rect 3466 23366 3478 23418
rect 3530 23366 3542 23418
rect 3594 23366 3606 23418
rect 3658 23366 8150 23418
rect 8202 23366 8214 23418
rect 8266 23366 8278 23418
rect 8330 23366 8342 23418
rect 8394 23366 8406 23418
rect 8458 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 17750 23418
rect 17802 23366 17814 23418
rect 17866 23366 17878 23418
rect 17930 23366 17942 23418
rect 17994 23366 18006 23418
rect 18058 23366 22550 23418
rect 22602 23366 22614 23418
rect 22666 23366 22678 23418
rect 22730 23366 22742 23418
rect 22794 23366 22806 23418
rect 22858 23366 27350 23418
rect 27402 23366 27414 23418
rect 27466 23366 27478 23418
rect 27530 23366 27542 23418
rect 27594 23366 27606 23418
rect 27658 23366 28888 23418
rect 1104 23344 28888 23366
rect 1104 22874 28888 22896
rect 1104 22822 5750 22874
rect 5802 22822 5814 22874
rect 5866 22822 5878 22874
rect 5930 22822 5942 22874
rect 5994 22822 6006 22874
rect 6058 22822 10550 22874
rect 10602 22822 10614 22874
rect 10666 22822 10678 22874
rect 10730 22822 10742 22874
rect 10794 22822 10806 22874
rect 10858 22822 15350 22874
rect 15402 22822 15414 22874
rect 15466 22822 15478 22874
rect 15530 22822 15542 22874
rect 15594 22822 15606 22874
rect 15658 22822 20150 22874
rect 20202 22822 20214 22874
rect 20266 22822 20278 22874
rect 20330 22822 20342 22874
rect 20394 22822 20406 22874
rect 20458 22822 24950 22874
rect 25002 22822 25014 22874
rect 25066 22822 25078 22874
rect 25130 22822 25142 22874
rect 25194 22822 25206 22874
rect 25258 22822 28888 22874
rect 1104 22800 28888 22822
rect 23569 22763 23627 22769
rect 23569 22729 23581 22763
rect 23615 22760 23627 22763
rect 24210 22760 24216 22772
rect 23615 22732 24216 22760
rect 23615 22729 23627 22732
rect 23569 22723 23627 22729
rect 24210 22720 24216 22732
rect 24268 22720 24274 22772
rect 23474 22652 23480 22704
rect 23532 22692 23538 22704
rect 23661 22695 23719 22701
rect 23661 22692 23673 22695
rect 23532 22664 23673 22692
rect 23532 22652 23538 22664
rect 23661 22661 23673 22664
rect 23707 22661 23719 22695
rect 23661 22655 23719 22661
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 3142 22624 3148 22636
rect 1811 22596 3148 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 3142 22584 3148 22596
rect 3200 22584 3206 22636
rect 25866 22624 25872 22636
rect 25827 22596 25872 22624
rect 25866 22584 25872 22596
rect 25924 22584 25930 22636
rect 23477 22559 23535 22565
rect 23477 22525 23489 22559
rect 23523 22525 23535 22559
rect 23477 22519 23535 22525
rect 23492 22488 23520 22519
rect 26602 22488 26608 22500
rect 23492 22460 26608 22488
rect 26602 22448 26608 22460
rect 26660 22448 26666 22500
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 24029 22423 24087 22429
rect 24029 22389 24041 22423
rect 24075 22420 24087 22423
rect 24118 22420 24124 22432
rect 24075 22392 24124 22420
rect 24075 22389 24087 22392
rect 24029 22383 24087 22389
rect 24118 22380 24124 22392
rect 24176 22380 24182 22432
rect 25682 22420 25688 22432
rect 25643 22392 25688 22420
rect 25682 22380 25688 22392
rect 25740 22380 25746 22432
rect 1104 22330 28888 22352
rect 1104 22278 3350 22330
rect 3402 22278 3414 22330
rect 3466 22278 3478 22330
rect 3530 22278 3542 22330
rect 3594 22278 3606 22330
rect 3658 22278 8150 22330
rect 8202 22278 8214 22330
rect 8266 22278 8278 22330
rect 8330 22278 8342 22330
rect 8394 22278 8406 22330
rect 8458 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 17750 22330
rect 17802 22278 17814 22330
rect 17866 22278 17878 22330
rect 17930 22278 17942 22330
rect 17994 22278 18006 22330
rect 18058 22278 22550 22330
rect 22602 22278 22614 22330
rect 22666 22278 22678 22330
rect 22730 22278 22742 22330
rect 22794 22278 22806 22330
rect 22858 22278 27350 22330
rect 27402 22278 27414 22330
rect 27466 22278 27478 22330
rect 27530 22278 27542 22330
rect 27594 22278 27606 22330
rect 27658 22278 28888 22330
rect 1104 22256 28888 22278
rect 22636 22219 22694 22225
rect 22636 22185 22648 22219
rect 22682 22216 22694 22219
rect 23934 22216 23940 22228
rect 22682 22188 23940 22216
rect 22682 22185 22694 22188
rect 22636 22179 22694 22185
rect 23934 22176 23940 22188
rect 23992 22176 23998 22228
rect 24121 22219 24179 22225
rect 24121 22185 24133 22219
rect 24167 22216 24179 22219
rect 24210 22216 24216 22228
rect 24167 22188 24216 22216
rect 24167 22185 24179 22188
rect 24121 22179 24179 22185
rect 24210 22176 24216 22188
rect 24268 22176 24274 22228
rect 25580 22219 25638 22225
rect 25580 22185 25592 22219
rect 25626 22216 25638 22219
rect 25682 22216 25688 22228
rect 25626 22188 25688 22216
rect 25626 22185 25638 22188
rect 25580 22179 25638 22185
rect 25682 22176 25688 22188
rect 25740 22176 25746 22228
rect 19150 22040 19156 22092
rect 19208 22080 19214 22092
rect 22373 22083 22431 22089
rect 22373 22080 22385 22083
rect 19208 22052 22385 22080
rect 19208 22040 19214 22052
rect 22373 22049 22385 22052
rect 22419 22080 22431 22083
rect 23658 22080 23664 22092
rect 22419 22052 23664 22080
rect 22419 22049 22431 22052
rect 22373 22043 22431 22049
rect 23658 22040 23664 22052
rect 23716 22040 23722 22092
rect 27065 22083 27123 22089
rect 27065 22049 27077 22083
rect 27111 22080 27123 22083
rect 27614 22080 27620 22092
rect 27111 22052 27620 22080
rect 27111 22049 27123 22052
rect 27065 22043 27123 22049
rect 27614 22040 27620 22052
rect 27672 22040 27678 22092
rect 27798 22080 27804 22092
rect 27759 22052 27804 22080
rect 27798 22040 27804 22052
rect 27856 22040 27862 22092
rect 27893 22083 27951 22089
rect 27893 22049 27905 22083
rect 27939 22049 27951 22083
rect 27893 22043 27951 22049
rect 19978 21972 19984 22024
rect 20036 22012 20042 22024
rect 20073 22015 20131 22021
rect 20073 22012 20085 22015
rect 20036 21984 20085 22012
rect 20036 21972 20042 21984
rect 20073 21981 20085 21984
rect 20119 21981 20131 22015
rect 25314 22012 25320 22024
rect 25275 21984 25320 22012
rect 20073 21975 20131 21981
rect 25314 21972 25320 21984
rect 25372 21972 25378 22024
rect 27338 21972 27344 22024
rect 27396 22012 27402 22024
rect 27908 22012 27936 22043
rect 27396 21984 27936 22012
rect 27396 21972 27402 21984
rect 26050 21944 26056 21956
rect 23874 21916 26056 21944
rect 26050 21904 26056 21916
rect 26108 21904 26114 21956
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 20257 21879 20315 21885
rect 20257 21876 20269 21879
rect 19484 21848 20269 21876
rect 19484 21836 19490 21848
rect 20257 21845 20269 21848
rect 20303 21876 20315 21879
rect 26326 21876 26332 21888
rect 20303 21848 26332 21876
rect 20303 21845 20315 21848
rect 20257 21839 20315 21845
rect 26326 21836 26332 21848
rect 26384 21836 26390 21888
rect 27246 21836 27252 21888
rect 27304 21876 27310 21888
rect 27341 21879 27399 21885
rect 27341 21876 27353 21879
rect 27304 21848 27353 21876
rect 27304 21836 27310 21848
rect 27341 21845 27353 21848
rect 27387 21845 27399 21879
rect 27706 21876 27712 21888
rect 27667 21848 27712 21876
rect 27341 21839 27399 21845
rect 27706 21836 27712 21848
rect 27764 21836 27770 21888
rect 1104 21786 28888 21808
rect 1104 21734 5750 21786
rect 5802 21734 5814 21786
rect 5866 21734 5878 21786
rect 5930 21734 5942 21786
rect 5994 21734 6006 21786
rect 6058 21734 10550 21786
rect 10602 21734 10614 21786
rect 10666 21734 10678 21786
rect 10730 21734 10742 21786
rect 10794 21734 10806 21786
rect 10858 21734 15350 21786
rect 15402 21734 15414 21786
rect 15466 21734 15478 21786
rect 15530 21734 15542 21786
rect 15594 21734 15606 21786
rect 15658 21734 20150 21786
rect 20202 21734 20214 21786
rect 20266 21734 20278 21786
rect 20330 21734 20342 21786
rect 20394 21734 20406 21786
rect 20458 21734 24950 21786
rect 25002 21734 25014 21786
rect 25066 21734 25078 21786
rect 25130 21734 25142 21786
rect 25194 21734 25206 21786
rect 25258 21734 28888 21786
rect 1104 21712 28888 21734
rect 3050 21632 3056 21684
rect 3108 21672 3114 21684
rect 3605 21675 3663 21681
rect 3605 21672 3617 21675
rect 3108 21644 3617 21672
rect 3108 21632 3114 21644
rect 3605 21641 3617 21644
rect 3651 21641 3663 21675
rect 3605 21635 3663 21641
rect 18230 21632 18236 21684
rect 18288 21672 18294 21684
rect 23934 21672 23940 21684
rect 18288 21644 23612 21672
rect 23895 21644 23940 21672
rect 18288 21632 18294 21644
rect 2774 21564 2780 21616
rect 2832 21564 2838 21616
rect 19426 21604 19432 21616
rect 19387 21576 19432 21604
rect 19426 21564 19432 21576
rect 19484 21564 19490 21616
rect 19518 21564 19524 21616
rect 19576 21604 19582 21616
rect 23385 21607 23443 21613
rect 19576 21576 19918 21604
rect 19576 21564 19582 21576
rect 23385 21573 23397 21607
rect 23431 21604 23443 21607
rect 23474 21604 23480 21616
rect 23431 21576 23480 21604
rect 23431 21573 23443 21576
rect 23385 21567 23443 21573
rect 23474 21564 23480 21576
rect 23532 21564 23538 21616
rect 23584 21604 23612 21644
rect 23934 21632 23940 21644
rect 23992 21632 23998 21684
rect 25866 21632 25872 21684
rect 25924 21672 25930 21684
rect 25961 21675 26019 21681
rect 25961 21672 25973 21675
rect 25924 21644 25973 21672
rect 25924 21632 25930 21644
rect 25961 21641 25973 21644
rect 26007 21641 26019 21675
rect 26326 21672 26332 21684
rect 26287 21644 26332 21672
rect 25961 21635 26019 21641
rect 26326 21632 26332 21644
rect 26384 21632 26390 21684
rect 26421 21675 26479 21681
rect 26421 21641 26433 21675
rect 26467 21672 26479 21675
rect 27614 21672 27620 21684
rect 26467 21644 27620 21672
rect 26467 21641 26479 21644
rect 26421 21635 26479 21641
rect 27614 21632 27620 21644
rect 27672 21632 27678 21684
rect 27706 21604 27712 21616
rect 23584 21576 27712 21604
rect 27706 21564 27712 21576
rect 27764 21564 27770 21616
rect 19150 21536 19156 21548
rect 19111 21508 19156 21536
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 24118 21536 24124 21548
rect 1762 21428 1768 21480
rect 1820 21468 1826 21480
rect 1857 21471 1915 21477
rect 1857 21468 1869 21471
rect 1820 21440 1869 21468
rect 1820 21428 1826 21440
rect 1857 21437 1869 21440
rect 1903 21437 1915 21471
rect 2130 21468 2136 21480
rect 2091 21440 2136 21468
rect 1857 21431 1915 21437
rect 2130 21428 2136 21440
rect 2188 21428 2194 21480
rect 19518 21428 19524 21480
rect 19576 21468 19582 21480
rect 22296 21468 22324 21522
rect 24079 21508 24124 21536
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 27246 21536 27252 21548
rect 27207 21508 27252 21536
rect 27246 21496 27252 21508
rect 27304 21496 27310 21548
rect 28166 21536 28172 21548
rect 28127 21508 28172 21536
rect 28166 21496 28172 21508
rect 28224 21496 28230 21548
rect 23658 21468 23664 21480
rect 19576 21440 22324 21468
rect 23571 21440 23664 21468
rect 19576 21428 19582 21440
rect 23658 21428 23664 21440
rect 23716 21468 23722 21480
rect 26602 21468 26608 21480
rect 23716 21440 26234 21468
rect 26515 21440 26608 21468
rect 23716 21428 23722 21440
rect 26206 21400 26234 21440
rect 26602 21428 26608 21440
rect 26660 21428 26666 21480
rect 26326 21400 26332 21412
rect 26206 21372 26332 21400
rect 26326 21360 26332 21372
rect 26384 21360 26390 21412
rect 26620 21400 26648 21428
rect 27246 21400 27252 21412
rect 26620 21372 27252 21400
rect 27246 21360 27252 21372
rect 27304 21360 27310 21412
rect 20438 21292 20444 21344
rect 20496 21332 20502 21344
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20496 21304 20913 21332
rect 20496 21292 20502 21304
rect 20901 21301 20913 21304
rect 20947 21301 20959 21335
rect 20901 21295 20959 21301
rect 21913 21335 21971 21341
rect 21913 21301 21925 21335
rect 21959 21332 21971 21335
rect 22370 21332 22376 21344
rect 21959 21304 22376 21332
rect 21959 21301 21971 21304
rect 21913 21295 21971 21301
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 26602 21292 26608 21344
rect 26660 21332 26666 21344
rect 27065 21335 27123 21341
rect 27065 21332 27077 21335
rect 26660 21304 27077 21332
rect 26660 21292 26666 21304
rect 27065 21301 27077 21304
rect 27111 21301 27123 21335
rect 28350 21332 28356 21344
rect 28311 21304 28356 21332
rect 27065 21295 27123 21301
rect 28350 21292 28356 21304
rect 28408 21292 28414 21344
rect 1104 21242 28888 21264
rect 1104 21190 3350 21242
rect 3402 21190 3414 21242
rect 3466 21190 3478 21242
rect 3530 21190 3542 21242
rect 3594 21190 3606 21242
rect 3658 21190 8150 21242
rect 8202 21190 8214 21242
rect 8266 21190 8278 21242
rect 8330 21190 8342 21242
rect 8394 21190 8406 21242
rect 8458 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 17750 21242
rect 17802 21190 17814 21242
rect 17866 21190 17878 21242
rect 17930 21190 17942 21242
rect 17994 21190 18006 21242
rect 18058 21190 22550 21242
rect 22602 21190 22614 21242
rect 22666 21190 22678 21242
rect 22730 21190 22742 21242
rect 22794 21190 22806 21242
rect 22858 21190 27350 21242
rect 27402 21190 27414 21242
rect 27466 21190 27478 21242
rect 27530 21190 27542 21242
rect 27594 21190 27606 21242
rect 27658 21190 28888 21242
rect 1104 21168 28888 21190
rect 3142 21088 3148 21140
rect 3200 21128 3206 21140
rect 3513 21131 3571 21137
rect 3513 21128 3525 21131
rect 3200 21100 3525 21128
rect 3200 21088 3206 21100
rect 3513 21097 3525 21100
rect 3559 21097 3571 21131
rect 19978 21128 19984 21140
rect 19939 21100 19984 21128
rect 3513 21091 3571 21097
rect 1762 20992 1768 21004
rect 1723 20964 1768 20992
rect 1762 20952 1768 20964
rect 1820 20992 1826 21004
rect 3234 20992 3240 21004
rect 1820 20964 3240 20992
rect 1820 20952 1826 20964
rect 3234 20952 3240 20964
rect 3292 20952 3298 21004
rect 3528 20992 3556 21091
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 22189 21131 22247 21137
rect 22189 21097 22201 21131
rect 22235 21128 22247 21131
rect 23474 21128 23480 21140
rect 22235 21100 23480 21128
rect 22235 21097 22247 21100
rect 22189 21091 22247 21097
rect 23474 21088 23480 21100
rect 23532 21088 23538 21140
rect 27798 21088 27804 21140
rect 27856 21128 27862 21140
rect 28077 21131 28135 21137
rect 28077 21128 28089 21131
rect 27856 21100 28089 21128
rect 27856 21088 27862 21100
rect 28077 21097 28089 21100
rect 28123 21097 28135 21131
rect 28077 21091 28135 21097
rect 4341 20995 4399 21001
rect 4341 20992 4353 20995
rect 3528 20964 4353 20992
rect 4341 20961 4353 20964
rect 4387 20961 4399 20995
rect 4341 20955 4399 20961
rect 4525 20995 4583 21001
rect 4525 20961 4537 20995
rect 4571 20992 4583 20995
rect 4890 20992 4896 21004
rect 4571 20964 4896 20992
rect 4571 20961 4583 20964
rect 4525 20955 4583 20961
rect 4890 20952 4896 20964
rect 4948 20952 4954 21004
rect 20438 20992 20444 21004
rect 20399 20964 20444 20992
rect 20438 20952 20444 20964
rect 20496 20952 20502 21004
rect 20625 20995 20683 21001
rect 20625 20961 20637 20995
rect 20671 20992 20683 20995
rect 20714 20992 20720 21004
rect 20671 20964 20720 20992
rect 20671 20961 20683 20964
rect 20625 20955 20683 20961
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 26602 20992 26608 21004
rect 26563 20964 26608 20992
rect 26602 20952 26608 20964
rect 26660 20952 26666 21004
rect 16850 20924 16856 20936
rect 16811 20896 16856 20924
rect 16850 20884 16856 20896
rect 16908 20884 16914 20936
rect 22002 20924 22008 20936
rect 21963 20896 22008 20924
rect 22002 20884 22008 20896
rect 22060 20884 22066 20936
rect 26326 20924 26332 20936
rect 26287 20896 26332 20924
rect 26326 20884 26332 20896
rect 26384 20884 26390 20936
rect 2038 20856 2044 20868
rect 1999 20828 2044 20856
rect 2038 20816 2044 20828
rect 2096 20816 2102 20868
rect 2774 20816 2780 20868
rect 2832 20816 2838 20868
rect 4249 20859 4307 20865
rect 4249 20825 4261 20859
rect 4295 20856 4307 20859
rect 6730 20856 6736 20868
rect 4295 20828 6736 20856
rect 4295 20825 4307 20828
rect 4249 20819 4307 20825
rect 6730 20816 6736 20828
rect 6788 20816 6794 20868
rect 26050 20856 26056 20868
rect 25963 20828 26056 20856
rect 26050 20816 26056 20828
rect 26108 20856 26114 20868
rect 26108 20828 26234 20856
rect 26108 20816 26114 20828
rect 3878 20788 3884 20800
rect 3839 20760 3884 20788
rect 3878 20748 3884 20760
rect 3936 20748 3942 20800
rect 4890 20788 4896 20800
rect 4851 20760 4896 20788
rect 4890 20748 4896 20760
rect 4948 20748 4954 20800
rect 17037 20791 17095 20797
rect 17037 20757 17049 20791
rect 17083 20788 17095 20791
rect 18230 20788 18236 20800
rect 17083 20760 18236 20788
rect 17083 20757 17095 20760
rect 17037 20751 17095 20757
rect 18230 20748 18236 20760
rect 18288 20748 18294 20800
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 20349 20791 20407 20797
rect 20349 20788 20361 20791
rect 19576 20760 20361 20788
rect 19576 20748 19582 20760
rect 20349 20757 20361 20760
rect 20395 20757 20407 20791
rect 26206 20788 26234 20828
rect 26712 20828 27094 20856
rect 26712 20788 26740 20828
rect 26206 20760 26740 20788
rect 20349 20751 20407 20757
rect 1104 20698 28888 20720
rect 1104 20646 5750 20698
rect 5802 20646 5814 20698
rect 5866 20646 5878 20698
rect 5930 20646 5942 20698
rect 5994 20646 6006 20698
rect 6058 20646 10550 20698
rect 10602 20646 10614 20698
rect 10666 20646 10678 20698
rect 10730 20646 10742 20698
rect 10794 20646 10806 20698
rect 10858 20646 15350 20698
rect 15402 20646 15414 20698
rect 15466 20646 15478 20698
rect 15530 20646 15542 20698
rect 15594 20646 15606 20698
rect 15658 20646 20150 20698
rect 20202 20646 20214 20698
rect 20266 20646 20278 20698
rect 20330 20646 20342 20698
rect 20394 20646 20406 20698
rect 20458 20646 24950 20698
rect 25002 20646 25014 20698
rect 25066 20646 25078 20698
rect 25130 20646 25142 20698
rect 25194 20646 25206 20698
rect 25258 20646 28888 20698
rect 1104 20624 28888 20646
rect 2130 20544 2136 20596
rect 2188 20584 2194 20596
rect 2317 20587 2375 20593
rect 2317 20584 2329 20587
rect 2188 20556 2329 20584
rect 2188 20544 2194 20556
rect 2317 20553 2329 20556
rect 2363 20553 2375 20587
rect 2317 20547 2375 20553
rect 3050 20544 3056 20596
rect 3108 20584 3114 20596
rect 3237 20587 3295 20593
rect 3237 20584 3249 20587
rect 3108 20556 3249 20584
rect 3108 20544 3114 20556
rect 3237 20553 3249 20556
rect 3283 20553 3295 20587
rect 3237 20547 3295 20553
rect 21913 20587 21971 20593
rect 21913 20553 21925 20587
rect 21959 20584 21971 20587
rect 22002 20584 22008 20596
rect 21959 20556 22008 20584
rect 21959 20553 21971 20556
rect 21913 20547 21971 20553
rect 22002 20544 22008 20556
rect 22060 20544 22066 20596
rect 22370 20584 22376 20596
rect 22331 20556 22376 20584
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 27065 20587 27123 20593
rect 27065 20553 27077 20587
rect 27111 20553 27123 20587
rect 27065 20547 27123 20553
rect 27525 20587 27583 20593
rect 27525 20553 27537 20587
rect 27571 20584 27583 20587
rect 28166 20584 28172 20596
rect 27571 20556 28172 20584
rect 27571 20553 27583 20556
rect 27525 20547 27583 20553
rect 18230 20516 18236 20528
rect 18191 20488 18236 20516
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 2501 20451 2559 20457
rect 2501 20417 2513 20451
rect 2547 20448 2559 20451
rect 3142 20448 3148 20460
rect 2547 20420 2820 20448
rect 3103 20420 3148 20448
rect 2547 20417 2559 20420
rect 2501 20411 2559 20417
rect 2792 20321 2820 20420
rect 3142 20408 3148 20420
rect 3200 20408 3206 20460
rect 17126 20408 17132 20460
rect 17184 20408 17190 20460
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20448 18567 20451
rect 19150 20448 19156 20460
rect 18555 20420 19156 20448
rect 18555 20417 18567 20420
rect 18509 20411 18567 20417
rect 19150 20408 19156 20420
rect 19208 20448 19214 20460
rect 19794 20448 19800 20460
rect 19208 20420 19800 20448
rect 19208 20408 19214 20420
rect 19794 20408 19800 20420
rect 19852 20408 19858 20460
rect 21266 20408 21272 20460
rect 21324 20448 21330 20460
rect 22281 20451 22339 20457
rect 22281 20448 22293 20451
rect 21324 20420 22293 20448
rect 21324 20408 21330 20420
rect 22281 20417 22293 20420
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 26697 20451 26755 20457
rect 26697 20417 26709 20451
rect 26743 20448 26755 20451
rect 27080 20448 27108 20547
rect 28166 20544 28172 20556
rect 28224 20544 28230 20596
rect 26743 20420 27108 20448
rect 27433 20451 27491 20457
rect 26743 20417 26755 20420
rect 26697 20411 26755 20417
rect 27433 20417 27445 20451
rect 27479 20417 27491 20451
rect 27433 20411 27491 20417
rect 3421 20383 3479 20389
rect 3421 20349 3433 20383
rect 3467 20380 3479 20383
rect 4890 20380 4896 20392
rect 3467 20352 4896 20380
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 2777 20315 2835 20321
rect 2777 20281 2789 20315
rect 2823 20281 2835 20315
rect 2777 20275 2835 20281
rect 3804 20256 3832 20352
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 22462 20380 22468 20392
rect 22423 20352 22468 20380
rect 22462 20340 22468 20352
rect 22520 20380 22526 20392
rect 22925 20383 22983 20389
rect 22925 20380 22937 20383
rect 22520 20352 22937 20380
rect 22520 20340 22526 20352
rect 22925 20349 22937 20352
rect 22971 20380 22983 20383
rect 24302 20380 24308 20392
rect 22971 20352 24308 20380
rect 22971 20349 22983 20352
rect 22925 20343 22983 20349
rect 24302 20340 24308 20352
rect 24360 20340 24366 20392
rect 24854 20340 24860 20392
rect 24912 20380 24918 20392
rect 27448 20380 27476 20411
rect 27617 20383 27675 20389
rect 27617 20380 27629 20383
rect 24912 20352 27476 20380
rect 27540 20352 27629 20380
rect 24912 20340 24918 20352
rect 27246 20272 27252 20324
rect 27304 20312 27310 20324
rect 27540 20312 27568 20352
rect 27617 20349 27629 20352
rect 27663 20349 27675 20383
rect 27617 20343 27675 20349
rect 27304 20284 27568 20312
rect 27304 20272 27310 20284
rect 3786 20244 3792 20256
rect 3747 20216 3792 20244
rect 3786 20204 3792 20216
rect 3844 20204 3850 20256
rect 16758 20244 16764 20256
rect 16719 20216 16764 20244
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 26418 20204 26424 20256
rect 26476 20244 26482 20256
rect 26513 20247 26571 20253
rect 26513 20244 26525 20247
rect 26476 20216 26525 20244
rect 26476 20204 26482 20216
rect 26513 20213 26525 20216
rect 26559 20213 26571 20247
rect 26513 20207 26571 20213
rect 1104 20154 28888 20176
rect 1104 20102 3350 20154
rect 3402 20102 3414 20154
rect 3466 20102 3478 20154
rect 3530 20102 3542 20154
rect 3594 20102 3606 20154
rect 3658 20102 8150 20154
rect 8202 20102 8214 20154
rect 8266 20102 8278 20154
rect 8330 20102 8342 20154
rect 8394 20102 8406 20154
rect 8458 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 17750 20154
rect 17802 20102 17814 20154
rect 17866 20102 17878 20154
rect 17930 20102 17942 20154
rect 17994 20102 18006 20154
rect 18058 20102 22550 20154
rect 22602 20102 22614 20154
rect 22666 20102 22678 20154
rect 22730 20102 22742 20154
rect 22794 20102 22806 20154
rect 22858 20102 27350 20154
rect 27402 20102 27414 20154
rect 27466 20102 27478 20154
rect 27530 20102 27542 20154
rect 27594 20102 27606 20154
rect 27658 20102 28888 20154
rect 1104 20080 28888 20102
rect 2038 20000 2044 20052
rect 2096 20040 2102 20052
rect 2409 20043 2467 20049
rect 2409 20040 2421 20043
rect 2096 20012 2421 20040
rect 2096 20000 2102 20012
rect 2409 20009 2421 20012
rect 2455 20009 2467 20043
rect 16850 20040 16856 20052
rect 16811 20012 16856 20040
rect 2409 20003 2467 20009
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 22005 20043 22063 20049
rect 22005 20009 22017 20043
rect 22051 20040 22063 20043
rect 22462 20040 22468 20052
rect 22051 20012 22468 20040
rect 22051 20009 22063 20012
rect 22005 20003 22063 20009
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 27893 20043 27951 20049
rect 27893 20009 27905 20043
rect 27939 20040 27951 20043
rect 28166 20040 28172 20052
rect 27939 20012 28172 20040
rect 27939 20009 27951 20012
rect 27893 20003 27951 20009
rect 28166 20000 28172 20012
rect 28224 20000 28230 20052
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 17313 19907 17371 19913
rect 17313 19904 17325 19907
rect 16816 19876 17325 19904
rect 16816 19864 16822 19876
rect 17313 19873 17325 19876
rect 17359 19873 17371 19907
rect 17313 19867 17371 19873
rect 17402 19864 17408 19916
rect 17460 19904 17466 19916
rect 20714 19904 20720 19916
rect 17460 19876 20720 19904
rect 17460 19864 17466 19876
rect 20714 19864 20720 19876
rect 20772 19904 20778 19916
rect 20772 19876 21772 19904
rect 20772 19864 20778 19876
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19836 2651 19839
rect 3878 19836 3884 19848
rect 2639 19808 3884 19836
rect 2639 19805 2651 19808
rect 2593 19799 2651 19805
rect 3878 19796 3884 19808
rect 3936 19796 3942 19848
rect 21744 19845 21772 19876
rect 23290 19864 23296 19916
rect 23348 19904 23354 19916
rect 25314 19904 25320 19916
rect 23348 19876 25320 19904
rect 23348 19864 23354 19876
rect 25314 19864 25320 19876
rect 25372 19904 25378 19916
rect 26145 19907 26203 19913
rect 26145 19904 26157 19907
rect 25372 19876 26157 19904
rect 25372 19864 25378 19876
rect 26145 19873 26157 19876
rect 26191 19873 26203 19907
rect 26418 19904 26424 19916
rect 26379 19876 26424 19904
rect 26145 19867 26203 19873
rect 26418 19864 26424 19876
rect 26476 19864 26482 19916
rect 21729 19839 21787 19845
rect 21729 19805 21741 19839
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 26252 19740 26910 19768
rect 26252 19712 26280 19740
rect 17221 19703 17279 19709
rect 17221 19669 17233 19703
rect 17267 19700 17279 19703
rect 17494 19700 17500 19712
rect 17267 19672 17500 19700
rect 17267 19669 17279 19672
rect 17221 19663 17279 19669
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 26234 19660 26240 19712
rect 26292 19660 26298 19712
rect 26804 19700 26832 19740
rect 27706 19700 27712 19712
rect 26804 19672 27712 19700
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 1104 19610 28888 19632
rect 1104 19558 5750 19610
rect 5802 19558 5814 19610
rect 5866 19558 5878 19610
rect 5930 19558 5942 19610
rect 5994 19558 6006 19610
rect 6058 19558 10550 19610
rect 10602 19558 10614 19610
rect 10666 19558 10678 19610
rect 10730 19558 10742 19610
rect 10794 19558 10806 19610
rect 10858 19558 15350 19610
rect 15402 19558 15414 19610
rect 15466 19558 15478 19610
rect 15530 19558 15542 19610
rect 15594 19558 15606 19610
rect 15658 19558 20150 19610
rect 20202 19558 20214 19610
rect 20266 19558 20278 19610
rect 20330 19558 20342 19610
rect 20394 19558 20406 19610
rect 20458 19558 24950 19610
rect 25002 19558 25014 19610
rect 25066 19558 25078 19610
rect 25130 19558 25142 19610
rect 25194 19558 25206 19610
rect 25258 19558 28888 19610
rect 1104 19536 28888 19558
rect 19334 19496 19340 19508
rect 18432 19468 19340 19496
rect 16574 19388 16580 19440
rect 16632 19428 16638 19440
rect 17126 19428 17132 19440
rect 16632 19400 17132 19428
rect 16632 19388 16638 19400
rect 17126 19388 17132 19400
rect 17184 19428 17190 19440
rect 18432 19428 18460 19468
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 19518 19496 19524 19508
rect 19479 19468 19524 19496
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 19352 19428 19380 19456
rect 17184 19400 18538 19428
rect 19352 19400 24058 19428
rect 17184 19388 17190 19400
rect 17218 19320 17224 19372
rect 17276 19360 17282 19372
rect 17773 19363 17831 19369
rect 17773 19360 17785 19363
rect 17276 19332 17785 19360
rect 17276 19320 17282 19332
rect 17773 19329 17785 19332
rect 17819 19329 17831 19363
rect 23290 19360 23296 19372
rect 23251 19332 23296 19360
rect 17773 19323 17831 19329
rect 23290 19320 23296 19332
rect 23348 19320 23354 19372
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19292 18107 19295
rect 18138 19292 18144 19304
rect 18095 19264 18144 19292
rect 18095 19261 18107 19264
rect 18049 19255 18107 19261
rect 18138 19252 18144 19264
rect 18196 19252 18202 19304
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 24854 19292 24860 19304
rect 23615 19264 24860 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 24946 19116 24952 19168
rect 25004 19156 25010 19168
rect 25041 19159 25099 19165
rect 25041 19156 25053 19159
rect 25004 19128 25053 19156
rect 25004 19116 25010 19128
rect 25041 19125 25053 19128
rect 25087 19125 25099 19159
rect 25041 19119 25099 19125
rect 1104 19066 28888 19088
rect 1104 19014 3350 19066
rect 3402 19014 3414 19066
rect 3466 19014 3478 19066
rect 3530 19014 3542 19066
rect 3594 19014 3606 19066
rect 3658 19014 8150 19066
rect 8202 19014 8214 19066
rect 8266 19014 8278 19066
rect 8330 19014 8342 19066
rect 8394 19014 8406 19066
rect 8458 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 17750 19066
rect 17802 19014 17814 19066
rect 17866 19014 17878 19066
rect 17930 19014 17942 19066
rect 17994 19014 18006 19066
rect 18058 19014 22550 19066
rect 22602 19014 22614 19066
rect 22666 19014 22678 19066
rect 22730 19014 22742 19066
rect 22794 19014 22806 19066
rect 22858 19014 27350 19066
rect 27402 19014 27414 19066
rect 27466 19014 27478 19066
rect 27530 19014 27542 19066
rect 27594 19014 27606 19066
rect 27658 19014 28888 19066
rect 1104 18992 28888 19014
rect 6730 18952 6736 18964
rect 6691 18924 6736 18952
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 18233 18955 18291 18961
rect 18233 18952 18245 18955
rect 18196 18924 18245 18952
rect 18196 18912 18202 18924
rect 18233 18921 18245 18924
rect 18279 18921 18291 18955
rect 18233 18915 18291 18921
rect 23937 18955 23995 18961
rect 23937 18921 23949 18955
rect 23983 18952 23995 18955
rect 24854 18952 24860 18964
rect 23983 18924 24860 18952
rect 23983 18921 23995 18924
rect 23937 18915 23995 18921
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 24489 18887 24547 18893
rect 24489 18853 24501 18887
rect 24535 18853 24547 18887
rect 24489 18847 24547 18853
rect 21266 18816 21272 18828
rect 21227 18788 21272 18816
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 3234 18708 3240 18760
rect 3292 18748 3298 18760
rect 4985 18751 5043 18757
rect 4985 18748 4997 18751
rect 3292 18720 4997 18748
rect 3292 18708 3298 18720
rect 4985 18717 4997 18720
rect 5031 18717 5043 18751
rect 4985 18711 5043 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 18782 18748 18788 18760
rect 18463 18720 18788 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 24121 18751 24179 18757
rect 24121 18717 24133 18751
rect 24167 18748 24179 18751
rect 24504 18748 24532 18847
rect 24946 18816 24952 18828
rect 24907 18788 24952 18816
rect 24946 18776 24952 18788
rect 25004 18776 25010 18828
rect 25041 18819 25099 18825
rect 25041 18785 25053 18819
rect 25087 18785 25099 18819
rect 25041 18779 25099 18785
rect 24167 18720 24532 18748
rect 24167 18717 24179 18720
rect 24121 18711 24179 18717
rect 5258 18680 5264 18692
rect 5219 18652 5264 18680
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 21100 18680 21128 18711
rect 21542 18680 21548 18692
rect 5644 18652 5750 18680
rect 21100 18652 21548 18680
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 3970 18612 3976 18624
rect 2832 18584 3976 18612
rect 2832 18572 2838 18584
rect 3970 18572 3976 18584
rect 4028 18612 4034 18624
rect 5644 18612 5672 18652
rect 21542 18640 21548 18652
rect 21600 18680 21606 18692
rect 24857 18683 24915 18689
rect 24857 18680 24869 18683
rect 21600 18652 24869 18680
rect 21600 18640 21606 18652
rect 24857 18649 24869 18652
rect 24903 18649 24915 18683
rect 25056 18680 25084 18779
rect 28166 18748 28172 18760
rect 28127 18720 28172 18748
rect 28166 18708 28172 18720
rect 28224 18708 28230 18760
rect 24857 18643 24915 18649
rect 24964 18652 25084 18680
rect 8294 18612 8300 18624
rect 4028 18584 8300 18612
rect 4028 18572 4034 18584
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 20898 18612 20904 18624
rect 20859 18584 20904 18612
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 24302 18572 24308 18624
rect 24360 18612 24366 18624
rect 24964 18612 24992 18652
rect 28350 18612 28356 18624
rect 24360 18584 24992 18612
rect 28311 18584 28356 18612
rect 24360 18572 24366 18584
rect 28350 18572 28356 18584
rect 28408 18572 28414 18624
rect 1104 18522 28888 18544
rect 1104 18470 5750 18522
rect 5802 18470 5814 18522
rect 5866 18470 5878 18522
rect 5930 18470 5942 18522
rect 5994 18470 6006 18522
rect 6058 18470 10550 18522
rect 10602 18470 10614 18522
rect 10666 18470 10678 18522
rect 10730 18470 10742 18522
rect 10794 18470 10806 18522
rect 10858 18470 15350 18522
rect 15402 18470 15414 18522
rect 15466 18470 15478 18522
rect 15530 18470 15542 18522
rect 15594 18470 15606 18522
rect 15658 18470 20150 18522
rect 20202 18470 20214 18522
rect 20266 18470 20278 18522
rect 20330 18470 20342 18522
rect 20394 18470 20406 18522
rect 20458 18470 24950 18522
rect 25002 18470 25014 18522
rect 25066 18470 25078 18522
rect 25130 18470 25142 18522
rect 25194 18470 25206 18522
rect 25258 18470 28888 18522
rect 1104 18448 28888 18470
rect 2961 18411 3019 18417
rect 2961 18377 2973 18411
rect 3007 18408 3019 18411
rect 3142 18408 3148 18420
rect 3007 18380 3148 18408
rect 3007 18377 3019 18380
rect 2961 18371 3019 18377
rect 3142 18368 3148 18380
rect 3200 18408 3206 18420
rect 4062 18408 4068 18420
rect 3200 18380 4068 18408
rect 3200 18368 3206 18380
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 21358 18368 21364 18420
rect 21416 18408 21422 18420
rect 21545 18411 21603 18417
rect 21545 18408 21557 18411
rect 21416 18380 21557 18408
rect 21416 18368 21422 18380
rect 21545 18377 21557 18380
rect 21591 18377 21603 18411
rect 24302 18408 24308 18420
rect 24263 18380 24308 18408
rect 21545 18371 21603 18377
rect 24302 18368 24308 18380
rect 24360 18368 24366 18420
rect 27065 18411 27123 18417
rect 27065 18377 27077 18411
rect 27111 18377 27123 18411
rect 27065 18371 27123 18377
rect 2774 18300 2780 18352
rect 2832 18340 2838 18352
rect 2832 18312 3266 18340
rect 2832 18300 2838 18312
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 7653 18343 7711 18349
rect 7653 18340 7665 18343
rect 7432 18312 7665 18340
rect 7432 18300 7438 18312
rect 7653 18309 7665 18312
rect 7699 18309 7711 18343
rect 7653 18303 7711 18309
rect 8294 18300 8300 18352
rect 8352 18300 8358 18352
rect 19334 18300 19340 18352
rect 19392 18340 19398 18352
rect 20530 18340 20536 18352
rect 19392 18312 20536 18340
rect 19392 18300 19398 18312
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 2222 18272 2228 18284
rect 2183 18244 2228 18272
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 19794 18272 19800 18284
rect 19755 18244 19800 18272
rect 19794 18232 19800 18244
rect 19852 18232 19858 18284
rect 26697 18275 26755 18281
rect 26697 18241 26709 18275
rect 26743 18272 26755 18275
rect 27080 18272 27108 18371
rect 26743 18244 27108 18272
rect 27433 18275 27491 18281
rect 26743 18241 26755 18244
rect 26697 18235 26755 18241
rect 27433 18241 27445 18275
rect 27479 18241 27491 18275
rect 27433 18235 27491 18241
rect 27525 18275 27583 18281
rect 27525 18241 27537 18275
rect 27571 18272 27583 18275
rect 28166 18272 28172 18284
rect 27571 18244 28172 18272
rect 27571 18241 27583 18244
rect 27525 18235 27583 18241
rect 4430 18204 4436 18216
rect 4391 18176 4436 18204
rect 4430 18164 4436 18176
rect 4488 18164 4494 18216
rect 4709 18207 4767 18213
rect 4709 18173 4721 18207
rect 4755 18204 4767 18207
rect 7377 18207 7435 18213
rect 7377 18204 7389 18207
rect 4755 18176 7389 18204
rect 4755 18173 4767 18176
rect 4709 18167 4767 18173
rect 7377 18173 7389 18176
rect 7423 18173 7435 18207
rect 7377 18167 7435 18173
rect 20073 18207 20131 18213
rect 20073 18173 20085 18207
rect 20119 18204 20131 18207
rect 20622 18204 20628 18216
rect 20119 18176 20628 18204
rect 20119 18173 20131 18176
rect 20073 18167 20131 18173
rect 2409 18071 2467 18077
rect 2409 18037 2421 18071
rect 2455 18068 2467 18071
rect 2866 18068 2872 18080
rect 2455 18040 2872 18068
rect 2455 18037 2467 18040
rect 2409 18031 2467 18037
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 3234 18028 3240 18080
rect 3292 18068 3298 18080
rect 4724 18068 4752 18167
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 24854 18164 24860 18216
rect 24912 18204 24918 18216
rect 27448 18204 27476 18235
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 27617 18207 27675 18213
rect 27617 18204 27629 18207
rect 24912 18176 27476 18204
rect 27540 18176 27629 18204
rect 24912 18164 24918 18176
rect 27246 18096 27252 18148
rect 27304 18136 27310 18148
rect 27540 18136 27568 18176
rect 27617 18173 27629 18176
rect 27663 18173 27675 18207
rect 27617 18167 27675 18173
rect 27304 18108 27568 18136
rect 27304 18096 27310 18108
rect 5074 18068 5080 18080
rect 3292 18040 4752 18068
rect 5035 18040 5080 18068
rect 3292 18028 3298 18040
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 9122 18068 9128 18080
rect 9083 18040 9128 18068
rect 9122 18028 9128 18040
rect 9180 18028 9186 18080
rect 20530 18028 20536 18080
rect 20588 18068 20594 18080
rect 21174 18068 21180 18080
rect 20588 18040 21180 18068
rect 20588 18028 20594 18040
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 26513 18071 26571 18077
rect 26513 18037 26525 18071
rect 26559 18068 26571 18071
rect 26602 18068 26608 18080
rect 26559 18040 26608 18068
rect 26559 18037 26571 18040
rect 26513 18031 26571 18037
rect 26602 18028 26608 18040
rect 26660 18028 26666 18080
rect 1104 17978 28888 18000
rect 1104 17926 3350 17978
rect 3402 17926 3414 17978
rect 3466 17926 3478 17978
rect 3530 17926 3542 17978
rect 3594 17926 3606 17978
rect 3658 17926 8150 17978
rect 8202 17926 8214 17978
rect 8266 17926 8278 17978
rect 8330 17926 8342 17978
rect 8394 17926 8406 17978
rect 8458 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 17750 17978
rect 17802 17926 17814 17978
rect 17866 17926 17878 17978
rect 17930 17926 17942 17978
rect 17994 17926 18006 17978
rect 18058 17926 22550 17978
rect 22602 17926 22614 17978
rect 22666 17926 22678 17978
rect 22730 17926 22742 17978
rect 22794 17926 22806 17978
rect 22858 17926 27350 17978
rect 27402 17926 27414 17978
rect 27466 17926 27478 17978
rect 27530 17926 27542 17978
rect 27594 17926 27606 17978
rect 27658 17926 28888 17978
rect 1104 17904 28888 17926
rect 4065 17867 4123 17873
rect 4065 17833 4077 17867
rect 4111 17864 4123 17867
rect 4430 17864 4436 17876
rect 4111 17836 4436 17864
rect 4111 17833 4123 17836
rect 4065 17827 4123 17833
rect 4430 17824 4436 17836
rect 4488 17824 4494 17876
rect 5258 17864 5264 17876
rect 5219 17836 5264 17864
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 24673 17867 24731 17873
rect 24673 17833 24685 17867
rect 24719 17864 24731 17867
rect 24854 17864 24860 17876
rect 24719 17836 24860 17864
rect 24719 17833 24731 17836
rect 24673 17827 24731 17833
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 28077 17867 28135 17873
rect 28077 17833 28089 17867
rect 28123 17864 28135 17867
rect 28166 17864 28172 17876
rect 28123 17836 28172 17864
rect 28123 17833 28135 17836
rect 28077 17827 28135 17833
rect 28166 17824 28172 17836
rect 28224 17824 28230 17876
rect 4338 17756 4344 17808
rect 4396 17756 4402 17808
rect 18138 17796 18144 17808
rect 18099 17768 18144 17796
rect 18138 17756 18144 17768
rect 18196 17756 18202 17808
rect 19518 17756 19524 17808
rect 19576 17796 19582 17808
rect 19978 17796 19984 17808
rect 19576 17768 19984 17796
rect 19576 17756 19582 17768
rect 19978 17756 19984 17768
rect 20036 17796 20042 17808
rect 20349 17799 20407 17805
rect 20349 17796 20361 17799
rect 20036 17768 20361 17796
rect 20036 17756 20042 17768
rect 20349 17765 20361 17768
rect 20395 17765 20407 17799
rect 20349 17759 20407 17765
rect 20806 17756 20812 17808
rect 20864 17796 20870 17808
rect 20901 17799 20959 17805
rect 20901 17796 20913 17799
rect 20864 17768 20913 17796
rect 20864 17756 20870 17768
rect 20901 17765 20913 17768
rect 20947 17765 20959 17799
rect 20901 17759 20959 17765
rect 2866 17688 2872 17740
rect 2924 17728 2930 17740
rect 2961 17731 3019 17737
rect 2961 17728 2973 17731
rect 2924 17700 2973 17728
rect 2924 17688 2930 17700
rect 2961 17697 2973 17700
rect 3007 17697 3019 17731
rect 3234 17728 3240 17740
rect 3195 17700 3240 17728
rect 2961 17691 3019 17697
rect 3234 17688 3240 17700
rect 3292 17688 3298 17740
rect 4356 17728 4384 17756
rect 21358 17728 21364 17740
rect 4356 17700 4473 17728
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4445 17669 4473 17700
rect 5460 17700 6684 17728
rect 21319 17700 21364 17728
rect 4341 17663 4399 17669
rect 4341 17660 4353 17663
rect 4120 17632 4353 17660
rect 4120 17620 4126 17632
rect 4341 17629 4353 17632
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 4430 17663 4488 17669
rect 4430 17629 4442 17663
rect 4476 17629 4488 17663
rect 4430 17623 4488 17629
rect 4522 17620 4528 17672
rect 4580 17660 4586 17672
rect 4709 17663 4767 17669
rect 4580 17632 4625 17660
rect 4580 17620 4586 17632
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 5074 17660 5080 17672
rect 4755 17632 5080 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 5074 17620 5080 17632
rect 5132 17660 5138 17672
rect 5258 17660 5264 17672
rect 5132 17632 5264 17660
rect 5132 17620 5138 17632
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 5460 17660 5488 17700
rect 5517 17663 5575 17669
rect 5517 17660 5529 17663
rect 5460 17632 5529 17660
rect 5517 17629 5529 17632
rect 5563 17629 5575 17663
rect 5517 17623 5575 17629
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17629 5687 17663
rect 5629 17623 5687 17629
rect 2682 17592 2688 17604
rect 2530 17564 2688 17592
rect 2682 17552 2688 17564
rect 2740 17552 2746 17604
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 4338 17484 4344 17536
rect 4396 17524 4402 17536
rect 5644 17524 5672 17623
rect 5718 17620 5724 17672
rect 5776 17660 5782 17672
rect 6656 17669 6684 17700
rect 21358 17688 21364 17700
rect 21416 17688 21422 17740
rect 26602 17728 26608 17740
rect 26563 17700 26608 17728
rect 26602 17688 26608 17700
rect 26660 17688 26666 17740
rect 5905 17663 5963 17669
rect 5776 17632 5821 17660
rect 5776 17620 5782 17632
rect 5905 17629 5917 17663
rect 5951 17660 5963 17663
rect 6641 17663 6699 17669
rect 5951 17632 6316 17660
rect 5951 17629 5963 17632
rect 5905 17623 5963 17629
rect 6288 17536 6316 17632
rect 6641 17629 6653 17663
rect 6687 17660 6699 17663
rect 6730 17660 6736 17672
rect 6687 17632 6736 17660
rect 6687 17629 6699 17632
rect 6641 17623 6699 17629
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 7650 17660 7656 17672
rect 7611 17632 7656 17660
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 8018 17660 8024 17672
rect 7979 17632 8024 17660
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 16482 17660 16488 17672
rect 16443 17632 16488 17660
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 17494 17660 17500 17672
rect 17455 17632 17500 17660
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 18230 17660 18236 17672
rect 18143 17632 18236 17660
rect 18230 17620 18236 17632
rect 18288 17660 18294 17672
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 18288 17632 19809 17660
rect 18288 17620 18294 17632
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17660 20039 17663
rect 20714 17660 20720 17672
rect 20027 17632 20720 17660
rect 20027 17629 20039 17632
rect 19981 17623 20039 17629
rect 20714 17620 20720 17632
rect 20772 17660 20778 17672
rect 20898 17660 20904 17672
rect 20772 17632 20904 17660
rect 20772 17620 20778 17632
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 21177 17663 21235 17669
rect 21177 17629 21189 17663
rect 21223 17629 21235 17663
rect 21177 17623 21235 17629
rect 6457 17595 6515 17601
rect 6457 17561 6469 17595
rect 6503 17592 6515 17595
rect 7742 17592 7748 17604
rect 6503 17564 7604 17592
rect 7703 17564 7748 17592
rect 6503 17561 6515 17564
rect 6457 17555 6515 17561
rect 6270 17524 6276 17536
rect 4396 17496 5672 17524
rect 6231 17496 6276 17524
rect 4396 17484 4402 17496
rect 6270 17484 6276 17496
rect 6328 17484 6334 17536
rect 7466 17524 7472 17536
rect 7427 17496 7472 17524
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 7576 17524 7604 17564
rect 7742 17552 7748 17564
rect 7800 17552 7806 17604
rect 7837 17595 7895 17601
rect 7837 17561 7849 17595
rect 7883 17592 7895 17595
rect 8478 17592 8484 17604
rect 7883 17564 8484 17592
rect 7883 17561 7895 17564
rect 7837 17555 7895 17561
rect 7852 17524 7880 17555
rect 8478 17552 8484 17564
rect 8536 17592 8542 17604
rect 9122 17592 9128 17604
rect 8536 17564 9128 17592
rect 8536 17552 8542 17564
rect 9122 17552 9128 17564
rect 9180 17552 9186 17604
rect 20073 17595 20131 17601
rect 20073 17561 20085 17595
rect 20119 17592 20131 17595
rect 21100 17592 21128 17623
rect 20119 17564 21128 17592
rect 21192 17592 21220 17623
rect 21266 17620 21272 17672
rect 21324 17660 21330 17672
rect 21542 17660 21548 17672
rect 21324 17632 21548 17660
rect 21324 17620 21330 17632
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 24486 17660 24492 17672
rect 24447 17632 24492 17660
rect 24486 17620 24492 17632
rect 24544 17620 24550 17672
rect 26326 17660 26332 17672
rect 26287 17632 26332 17660
rect 26326 17620 26332 17632
rect 26384 17620 26390 17672
rect 27706 17620 27712 17672
rect 27764 17620 27770 17672
rect 21450 17592 21456 17604
rect 21192 17564 21456 17592
rect 20119 17561 20131 17564
rect 20073 17555 20131 17561
rect 7576 17496 7880 17524
rect 15838 17484 15844 17536
rect 15896 17524 15902 17536
rect 16301 17527 16359 17533
rect 16301 17524 16313 17527
rect 15896 17496 16313 17524
rect 15896 17484 15902 17496
rect 16301 17493 16313 17496
rect 16347 17493 16359 17527
rect 16301 17487 16359 17493
rect 19794 17484 19800 17536
rect 19852 17524 19858 17536
rect 20088 17524 20116 17555
rect 19852 17496 20116 17524
rect 20165 17527 20223 17533
rect 19852 17484 19858 17496
rect 20165 17493 20177 17527
rect 20211 17524 20223 17527
rect 20530 17524 20536 17536
rect 20211 17496 20536 17524
rect 20211 17493 20223 17496
rect 20165 17487 20223 17493
rect 20530 17484 20536 17496
rect 20588 17524 20594 17536
rect 21192 17524 21220 17564
rect 21450 17552 21456 17564
rect 21508 17552 21514 17604
rect 20588 17496 21220 17524
rect 20588 17484 20594 17496
rect 1104 17434 28888 17456
rect 1104 17382 5750 17434
rect 5802 17382 5814 17434
rect 5866 17382 5878 17434
rect 5930 17382 5942 17434
rect 5994 17382 6006 17434
rect 6058 17382 10550 17434
rect 10602 17382 10614 17434
rect 10666 17382 10678 17434
rect 10730 17382 10742 17434
rect 10794 17382 10806 17434
rect 10858 17382 15350 17434
rect 15402 17382 15414 17434
rect 15466 17382 15478 17434
rect 15530 17382 15542 17434
rect 15594 17382 15606 17434
rect 15658 17382 20150 17434
rect 20202 17382 20214 17434
rect 20266 17382 20278 17434
rect 20330 17382 20342 17434
rect 20394 17382 20406 17434
rect 20458 17382 24950 17434
rect 25002 17382 25014 17434
rect 25066 17382 25078 17434
rect 25130 17382 25142 17434
rect 25194 17382 25206 17434
rect 25258 17382 28888 17434
rect 1104 17360 28888 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 2222 17320 2228 17332
rect 2183 17292 2228 17320
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 7926 17320 7932 17332
rect 5276 17292 7932 17320
rect 2685 17255 2743 17261
rect 2685 17252 2697 17255
rect 1780 17224 2697 17252
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 1780 17193 1808 17224
rect 2685 17221 2697 17224
rect 2731 17221 2743 17255
rect 2685 17215 2743 17221
rect 4062 17212 4068 17264
rect 4120 17252 4126 17264
rect 5276 17261 5304 17292
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 18601 17323 18659 17329
rect 18601 17289 18613 17323
rect 18647 17320 18659 17323
rect 19521 17323 19579 17329
rect 19521 17320 19533 17323
rect 18647 17292 19533 17320
rect 18647 17289 18659 17292
rect 18601 17283 18659 17289
rect 19521 17289 19533 17292
rect 19567 17289 19579 17323
rect 20530 17320 20536 17332
rect 19521 17283 19579 17289
rect 19996 17292 20536 17320
rect 5077 17255 5135 17261
rect 5077 17252 5089 17255
rect 4120 17224 5089 17252
rect 4120 17212 4126 17224
rect 5077 17221 5089 17224
rect 5123 17221 5135 17255
rect 5077 17215 5135 17221
rect 5261 17255 5319 17261
rect 5261 17221 5273 17255
rect 5307 17221 5319 17255
rect 5261 17215 5319 17221
rect 7466 17212 7472 17264
rect 7524 17252 7530 17264
rect 7837 17255 7895 17261
rect 7837 17252 7849 17255
rect 7524 17224 7849 17252
rect 7524 17212 7530 17224
rect 7837 17221 7849 17224
rect 7883 17221 7895 17255
rect 7837 17215 7895 17221
rect 8570 17212 8576 17264
rect 8628 17212 8634 17264
rect 12805 17255 12863 17261
rect 12805 17252 12817 17255
rect 12406 17224 12817 17252
rect 1765 17187 1823 17193
rect 1765 17184 1777 17187
rect 1544 17156 1777 17184
rect 1544 17144 1550 17156
rect 1765 17153 1777 17156
rect 1811 17153 1823 17187
rect 2590 17184 2596 17196
rect 2551 17156 2596 17184
rect 1765 17147 1823 17153
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 3329 17119 3387 17125
rect 3329 17116 3341 17119
rect 2915 17088 3341 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 3329 17085 3341 17088
rect 3375 17116 3387 17119
rect 3786 17116 3792 17128
rect 3375 17088 3792 17116
rect 3375 17085 3387 17088
rect 3329 17079 3387 17085
rect 3786 17076 3792 17088
rect 3844 17116 3850 17128
rect 4062 17116 4068 17128
rect 3844 17088 4068 17116
rect 3844 17076 3850 17088
rect 4062 17076 4068 17088
rect 4120 17116 4126 17128
rect 7558 17116 7564 17128
rect 4120 17088 6132 17116
rect 7519 17088 7564 17116
rect 4120 17076 4126 17088
rect 5258 17008 5264 17060
rect 5316 17048 5322 17060
rect 5534 17048 5540 17060
rect 5316 17020 5540 17048
rect 5316 17008 5322 17020
rect 5534 17008 5540 17020
rect 5592 17048 5598 17060
rect 5997 17051 6055 17057
rect 5997 17048 6009 17051
rect 5592 17020 6009 17048
rect 5592 17008 5598 17020
rect 5997 17017 6009 17020
rect 6043 17017 6055 17051
rect 6104 17048 6132 17088
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 10042 17116 10048 17128
rect 7668 17088 10048 17116
rect 7668 17048 7696 17088
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 6104 17020 7696 17048
rect 5997 17011 6055 17017
rect 12406 16992 12434 17224
rect 12805 17221 12817 17224
rect 12851 17252 12863 17255
rect 15102 17252 15108 17264
rect 12851 17224 13570 17252
rect 14936 17224 15108 17252
rect 12851 17221 12863 17224
rect 12805 17215 12863 17221
rect 14936 17193 14964 17224
rect 15102 17212 15108 17224
rect 15160 17252 15166 17264
rect 17218 17252 17224 17264
rect 15160 17224 17224 17252
rect 15160 17212 15166 17224
rect 17218 17212 17224 17224
rect 17276 17212 17282 17264
rect 17313 17255 17371 17261
rect 17313 17221 17325 17255
rect 17359 17252 17371 17255
rect 17494 17252 17500 17264
rect 17359 17224 17500 17252
rect 17359 17221 17371 17224
rect 17313 17215 17371 17221
rect 17494 17212 17500 17224
rect 17552 17212 17558 17264
rect 19996 17252 20024 17292
rect 20530 17280 20536 17292
rect 20588 17280 20594 17332
rect 20993 17323 21051 17329
rect 20993 17320 21005 17323
rect 20640 17292 21005 17320
rect 19904 17224 20024 17252
rect 14921 17187 14979 17193
rect 14921 17153 14933 17187
rect 14967 17153 14979 17187
rect 14921 17147 14979 17153
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17184 16175 17187
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 16163 17156 17141 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 18230 17184 18236 17196
rect 18191 17156 18236 17184
rect 17129 17147 17187 17153
rect 14550 17116 14556 17128
rect 14511 17088 14556 17116
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 15565 17119 15623 17125
rect 15565 17085 15577 17119
rect 15611 17116 15623 17119
rect 15746 17116 15752 17128
rect 15611 17088 15752 17116
rect 15611 17085 15623 17088
rect 15565 17079 15623 17085
rect 15746 17076 15752 17088
rect 15804 17076 15810 17128
rect 15948 17116 15976 17147
rect 16942 17116 16948 17128
rect 15948 17088 16948 17116
rect 16942 17076 16948 17088
rect 17000 17076 17006 17128
rect 17144 17116 17172 17147
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 19794 17184 19800 17196
rect 19755 17156 19800 17184
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 19904 17193 19932 17224
rect 20070 17212 20076 17264
rect 20128 17252 20134 17264
rect 20640 17261 20668 17292
rect 20993 17289 21005 17292
rect 21039 17289 21051 17323
rect 24762 17320 24768 17332
rect 20993 17283 21051 17289
rect 23768 17292 24768 17320
rect 23768 17261 23796 17292
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 20441 17255 20499 17261
rect 20441 17252 20453 17255
rect 20128 17224 20453 17252
rect 20128 17212 20134 17224
rect 20441 17221 20453 17224
rect 20487 17221 20499 17255
rect 20441 17215 20499 17221
rect 20625 17255 20683 17261
rect 20625 17221 20637 17255
rect 20671 17221 20683 17255
rect 20625 17215 20683 17221
rect 23753 17255 23811 17261
rect 23753 17221 23765 17255
rect 23799 17221 23811 17255
rect 26050 17252 26056 17264
rect 24978 17238 26056 17252
rect 23753 17215 23811 17221
rect 24964 17224 26056 17238
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17184 20039 17187
rect 20162 17184 20168 17196
rect 20027 17156 20168 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 20162 17144 20168 17156
rect 20220 17144 20226 17196
rect 20349 17187 20407 17193
rect 20349 17153 20361 17187
rect 20395 17184 20407 17187
rect 20714 17184 20720 17196
rect 20395 17156 20720 17184
rect 20395 17153 20407 17156
rect 20349 17147 20407 17153
rect 18248 17116 18276 17144
rect 17144 17088 18276 17116
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 19751 17088 20024 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 15194 17008 15200 17060
rect 15252 17048 15258 17060
rect 15657 17051 15715 17057
rect 15657 17048 15669 17051
rect 15252 17020 15669 17048
rect 15252 17008 15258 17020
rect 15657 17017 15669 17020
rect 15703 17017 15715 17051
rect 19334 17048 19340 17060
rect 15657 17011 15715 17017
rect 18616 17020 19340 17048
rect 4522 16940 4528 16992
rect 4580 16980 4586 16992
rect 5445 16983 5503 16989
rect 5445 16980 5457 16983
rect 4580 16952 5457 16980
rect 4580 16940 4586 16952
rect 5445 16949 5457 16952
rect 5491 16980 5503 16983
rect 5626 16980 5632 16992
rect 5491 16952 5632 16980
rect 5491 16949 5503 16952
rect 5445 16943 5503 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 9306 16980 9312 16992
rect 9267 16952 9312 16980
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 9824 16952 10333 16980
rect 9824 16940 9830 16952
rect 10321 16949 10333 16952
rect 10367 16980 10379 16983
rect 10870 16980 10876 16992
rect 10367 16952 10876 16980
rect 10367 16949 10379 16952
rect 10321 16943 10379 16949
rect 10870 16940 10876 16952
rect 10928 16980 10934 16992
rect 11609 16983 11667 16989
rect 11609 16980 11621 16983
rect 10928 16952 11621 16980
rect 10928 16940 10934 16952
rect 11609 16949 11621 16952
rect 11655 16980 11667 16983
rect 12342 16980 12348 16992
rect 11655 16952 12348 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 12342 16940 12348 16952
rect 12400 16952 12434 16992
rect 12400 16940 12406 16952
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 13127 16983 13185 16989
rect 13127 16980 13139 16983
rect 12860 16952 13139 16980
rect 12860 16940 12866 16952
rect 13127 16949 13139 16952
rect 13173 16949 13185 16983
rect 13127 16943 13185 16949
rect 17497 16983 17555 16989
rect 17497 16949 17509 16983
rect 17543 16980 17555 16983
rect 17586 16980 17592 16992
rect 17543 16952 17592 16980
rect 17543 16949 17555 16952
rect 17497 16943 17555 16949
rect 17586 16940 17592 16952
rect 17644 16940 17650 16992
rect 18616 16989 18644 17020
rect 19334 17008 19340 17020
rect 19392 17008 19398 17060
rect 19996 17048 20024 17088
rect 20364 17048 20392 17147
rect 20714 17144 20720 17156
rect 20772 17144 20778 17196
rect 20806 17144 20812 17196
rect 20864 17184 20870 17196
rect 20901 17187 20959 17193
rect 20901 17184 20913 17187
rect 20864 17156 20913 17184
rect 20864 17144 20870 17156
rect 20901 17153 20913 17156
rect 20947 17153 20959 17187
rect 20901 17147 20959 17153
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 21048 17156 21097 17184
rect 21048 17144 21054 17156
rect 21085 17153 21097 17156
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 23290 17144 23296 17196
rect 23348 17184 23354 17196
rect 23477 17187 23535 17193
rect 23477 17184 23489 17187
rect 23348 17156 23489 17184
rect 23348 17144 23354 17156
rect 23477 17153 23489 17156
rect 23523 17153 23535 17187
rect 23477 17147 23535 17153
rect 23106 17076 23112 17128
rect 23164 17116 23170 17128
rect 23201 17119 23259 17125
rect 23201 17116 23213 17119
rect 23164 17088 23213 17116
rect 23164 17076 23170 17088
rect 23201 17085 23213 17088
rect 23247 17116 23259 17119
rect 24964 17116 24992 17224
rect 26050 17212 26056 17224
rect 26108 17212 26114 17264
rect 23247 17088 24992 17116
rect 23247 17085 23259 17088
rect 23201 17079 23259 17085
rect 20622 17048 20628 17060
rect 19996 17020 20392 17048
rect 20583 17020 20628 17048
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 18601 16983 18659 16989
rect 18601 16949 18613 16983
rect 18647 16949 18659 16983
rect 18782 16980 18788 16992
rect 18743 16952 18788 16980
rect 18601 16943 18659 16949
rect 18782 16940 18788 16952
rect 18840 16940 18846 16992
rect 19978 16940 19984 16992
rect 20036 16980 20042 16992
rect 20162 16980 20168 16992
rect 20036 16952 20168 16980
rect 20036 16940 20042 16952
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 24946 16940 24952 16992
rect 25004 16980 25010 16992
rect 25225 16983 25283 16989
rect 25225 16980 25237 16983
rect 25004 16952 25237 16980
rect 25004 16940 25010 16952
rect 25225 16949 25237 16952
rect 25271 16949 25283 16983
rect 25225 16943 25283 16949
rect 1104 16890 28888 16912
rect 1104 16838 3350 16890
rect 3402 16838 3414 16890
rect 3466 16838 3478 16890
rect 3530 16838 3542 16890
rect 3594 16838 3606 16890
rect 3658 16838 8150 16890
rect 8202 16838 8214 16890
rect 8266 16838 8278 16890
rect 8330 16838 8342 16890
rect 8394 16838 8406 16890
rect 8458 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 17750 16890
rect 17802 16838 17814 16890
rect 17866 16838 17878 16890
rect 17930 16838 17942 16890
rect 17994 16838 18006 16890
rect 18058 16838 22550 16890
rect 22602 16838 22614 16890
rect 22666 16838 22678 16890
rect 22730 16838 22742 16890
rect 22794 16838 22806 16890
rect 22858 16838 27350 16890
rect 27402 16838 27414 16890
rect 27466 16838 27478 16890
rect 27530 16838 27542 16890
rect 27594 16838 27606 16890
rect 27658 16838 28888 16890
rect 1104 16816 28888 16838
rect 14185 16779 14243 16785
rect 14185 16745 14197 16779
rect 14231 16776 14243 16779
rect 14550 16776 14556 16788
rect 14231 16748 14556 16776
rect 14231 16745 14243 16748
rect 14185 16739 14243 16745
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 17497 16779 17555 16785
rect 17497 16776 17509 16779
rect 16540 16748 17509 16776
rect 16540 16736 16546 16748
rect 17497 16745 17509 16748
rect 17543 16745 17555 16779
rect 17497 16739 17555 16745
rect 17681 16779 17739 16785
rect 17681 16745 17693 16779
rect 17727 16776 17739 16779
rect 19150 16776 19156 16788
rect 17727 16748 19156 16776
rect 17727 16745 17739 16748
rect 17681 16739 17739 16745
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 24118 16776 24124 16788
rect 24031 16748 24124 16776
rect 24118 16736 24124 16748
rect 24176 16776 24182 16788
rect 24302 16776 24308 16788
rect 24176 16748 24308 16776
rect 24176 16736 24182 16748
rect 24302 16736 24308 16748
rect 24360 16736 24366 16788
rect 24486 16776 24492 16788
rect 24447 16748 24492 16776
rect 24486 16736 24492 16748
rect 24544 16736 24550 16788
rect 24578 16668 24584 16720
rect 24636 16708 24642 16720
rect 24636 16680 25084 16708
rect 24636 16668 24642 16680
rect 8478 16640 8484 16652
rect 7576 16612 8484 16640
rect 7576 16581 7604 16612
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 12250 16640 12256 16652
rect 10551 16612 12256 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 12860 16612 14688 16640
rect 12860 16600 12866 16612
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16541 7619 16575
rect 7926 16572 7932 16584
rect 7887 16544 7932 16572
rect 7561 16535 7619 16541
rect 7926 16532 7932 16544
rect 7984 16572 7990 16584
rect 8202 16572 8208 16584
rect 7984 16544 8208 16572
rect 7984 16532 7990 16544
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 9674 16572 9680 16584
rect 8312 16544 9680 16572
rect 7653 16507 7711 16513
rect 7653 16473 7665 16507
rect 7699 16473 7711 16507
rect 7653 16467 7711 16473
rect 7745 16507 7803 16513
rect 7745 16473 7757 16507
rect 7791 16504 7803 16507
rect 8018 16504 8024 16516
rect 7791 16476 8024 16504
rect 7791 16473 7803 16476
rect 7745 16467 7803 16473
rect 7374 16436 7380 16448
rect 7335 16408 7380 16436
rect 7374 16396 7380 16408
rect 7432 16396 7438 16448
rect 7668 16436 7696 16467
rect 8018 16464 8024 16476
rect 8076 16504 8082 16516
rect 8312 16504 8340 16544
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16572 10103 16575
rect 10410 16572 10416 16584
rect 10091 16544 10416 16572
rect 10091 16541 10103 16544
rect 10045 16535 10103 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 14660 16581 14688 16612
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15197 16643 15255 16649
rect 15197 16640 15209 16643
rect 15160 16612 15209 16640
rect 15160 16600 15166 16612
rect 15197 16609 15209 16612
rect 15243 16609 15255 16643
rect 15197 16603 15255 16609
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16640 15531 16643
rect 15838 16640 15844 16652
rect 15519 16612 15844 16640
rect 15519 16609 15531 16612
rect 15473 16603 15531 16609
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 16942 16640 16948 16652
rect 16855 16612 16948 16640
rect 16942 16600 16948 16612
rect 17000 16640 17006 16652
rect 17494 16640 17500 16652
rect 17000 16612 17500 16640
rect 17000 16600 17006 16612
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 19150 16600 19156 16652
rect 19208 16640 19214 16652
rect 21729 16643 21787 16649
rect 19208 16612 19564 16640
rect 19208 16600 19214 16612
rect 14369 16575 14427 16581
rect 14369 16572 14381 16575
rect 12124 16544 14381 16572
rect 12124 16532 12130 16544
rect 14369 16541 14381 16544
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16574 14703 16575
rect 14691 16546 14725 16574
rect 14826 16572 14832 16584
rect 14691 16541 14703 16546
rect 14787 16544 14832 16572
rect 14645 16535 14703 16541
rect 8076 16476 8340 16504
rect 8076 16464 8082 16476
rect 9122 16464 9128 16516
rect 9180 16504 9186 16516
rect 9861 16507 9919 16513
rect 9861 16504 9873 16507
rect 9180 16476 9873 16504
rect 9180 16464 9186 16476
rect 9861 16473 9873 16476
rect 9907 16473 9919 16507
rect 9861 16467 9919 16473
rect 9950 16464 9956 16516
rect 10008 16504 10014 16516
rect 10781 16507 10839 16513
rect 10008 16476 10053 16504
rect 10008 16464 10014 16476
rect 10781 16473 10793 16507
rect 10827 16473 10839 16507
rect 10781 16467 10839 16473
rect 7834 16436 7840 16448
rect 7668 16408 7840 16436
rect 7834 16396 7840 16408
rect 7892 16436 7898 16448
rect 9968 16436 9996 16464
rect 7892 16408 9996 16436
rect 10229 16439 10287 16445
rect 7892 16396 7898 16408
rect 10229 16405 10241 16439
rect 10275 16436 10287 16439
rect 10796 16436 10824 16467
rect 10870 16464 10876 16516
rect 10928 16504 10934 16516
rect 14384 16504 14412 16535
rect 14826 16532 14832 16544
rect 14884 16532 14890 16584
rect 16574 16532 16580 16584
rect 16632 16532 16638 16584
rect 19337 16575 19395 16581
rect 19337 16541 19349 16575
rect 19383 16572 19395 16575
rect 19426 16572 19432 16584
rect 19383 16544 19432 16572
rect 19383 16541 19395 16544
rect 19337 16535 19395 16541
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 15194 16504 15200 16516
rect 10928 16476 11270 16504
rect 14384 16476 15200 16504
rect 10928 16464 10934 16476
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 17678 16513 17684 16516
rect 17665 16507 17684 16513
rect 17665 16473 17677 16507
rect 17665 16467 17684 16473
rect 17678 16464 17684 16467
rect 17736 16464 17742 16516
rect 17865 16507 17923 16513
rect 17865 16473 17877 16507
rect 17911 16473 17923 16507
rect 17865 16467 17923 16473
rect 10275 16408 10824 16436
rect 10275 16405 10287 16408
rect 10229 16399 10287 16405
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 12253 16439 12311 16445
rect 12253 16436 12265 16439
rect 12216 16408 12265 16436
rect 12216 16396 12222 16408
rect 12253 16405 12265 16408
rect 12299 16405 12311 16439
rect 17880 16436 17908 16467
rect 18138 16464 18144 16516
rect 18196 16504 18202 16516
rect 18690 16504 18696 16516
rect 18196 16476 18696 16504
rect 18196 16464 18202 16476
rect 18690 16464 18696 16476
rect 18748 16464 18754 16516
rect 18230 16436 18236 16448
rect 17880 16408 18236 16436
rect 12253 16399 12311 16405
rect 18230 16396 18236 16408
rect 18288 16436 18294 16448
rect 19536 16445 19564 16612
rect 21729 16609 21741 16643
rect 21775 16640 21787 16643
rect 22002 16640 22008 16652
rect 21775 16612 22008 16640
rect 21775 16609 21787 16612
rect 21729 16603 21787 16609
rect 22002 16600 22008 16612
rect 22060 16640 22066 16652
rect 23290 16640 23296 16652
rect 22060 16612 23296 16640
rect 22060 16600 22066 16612
rect 23290 16600 23296 16612
rect 23348 16640 23354 16652
rect 25056 16649 25084 16680
rect 25041 16643 25099 16649
rect 23348 16612 24992 16640
rect 23348 16600 23354 16612
rect 24854 16572 24860 16584
rect 23138 16544 24860 16572
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 24964 16572 24992 16612
rect 25041 16609 25053 16643
rect 25087 16609 25099 16643
rect 25041 16603 25099 16609
rect 26602 16572 26608 16584
rect 24964 16544 26608 16572
rect 26602 16532 26608 16544
rect 26660 16532 26666 16584
rect 28166 16572 28172 16584
rect 28127 16544 28172 16572
rect 28166 16532 28172 16544
rect 28224 16532 28230 16584
rect 22005 16507 22063 16513
rect 22005 16473 22017 16507
rect 22051 16504 22063 16507
rect 22094 16504 22100 16516
rect 22051 16476 22100 16504
rect 22051 16473 22063 16476
rect 22005 16467 22063 16473
rect 22094 16464 22100 16476
rect 22152 16464 22158 16516
rect 24946 16504 24952 16516
rect 24907 16476 24952 16504
rect 24946 16464 24952 16476
rect 25004 16464 25010 16516
rect 18417 16439 18475 16445
rect 18417 16436 18429 16439
rect 18288 16408 18429 16436
rect 18288 16396 18294 16408
rect 18417 16405 18429 16408
rect 18463 16405 18475 16439
rect 18417 16399 18475 16405
rect 19521 16439 19579 16445
rect 19521 16405 19533 16439
rect 19567 16405 19579 16439
rect 19521 16399 19579 16405
rect 22186 16396 22192 16448
rect 22244 16436 22250 16448
rect 23477 16439 23535 16445
rect 23477 16436 23489 16439
rect 22244 16408 23489 16436
rect 22244 16396 22250 16408
rect 23477 16405 23489 16408
rect 23523 16436 23535 16439
rect 24857 16439 24915 16445
rect 24857 16436 24869 16439
rect 23523 16408 24869 16436
rect 23523 16405 23535 16408
rect 23477 16399 23535 16405
rect 24857 16405 24869 16408
rect 24903 16405 24915 16439
rect 28350 16436 28356 16448
rect 28311 16408 28356 16436
rect 24857 16399 24915 16405
rect 28350 16396 28356 16408
rect 28408 16396 28414 16448
rect 1104 16346 28888 16368
rect 1104 16294 5750 16346
rect 5802 16294 5814 16346
rect 5866 16294 5878 16346
rect 5930 16294 5942 16346
rect 5994 16294 6006 16346
rect 6058 16294 10550 16346
rect 10602 16294 10614 16346
rect 10666 16294 10678 16346
rect 10730 16294 10742 16346
rect 10794 16294 10806 16346
rect 10858 16294 15350 16346
rect 15402 16294 15414 16346
rect 15466 16294 15478 16346
rect 15530 16294 15542 16346
rect 15594 16294 15606 16346
rect 15658 16294 20150 16346
rect 20202 16294 20214 16346
rect 20266 16294 20278 16346
rect 20330 16294 20342 16346
rect 20394 16294 20406 16346
rect 20458 16294 24950 16346
rect 25002 16294 25014 16346
rect 25066 16294 25078 16346
rect 25130 16294 25142 16346
rect 25194 16294 25206 16346
rect 25258 16294 28888 16346
rect 1104 16272 28888 16294
rect 7742 16192 7748 16244
rect 7800 16192 7806 16244
rect 12802 16232 12808 16244
rect 9508 16204 12808 16232
rect 4617 16167 4675 16173
rect 4617 16164 4629 16167
rect 3988 16136 4629 16164
rect 2590 16056 2596 16108
rect 2648 16096 2654 16108
rect 3988 16105 4016 16136
rect 4617 16133 4629 16136
rect 4663 16133 4675 16167
rect 7760 16164 7788 16192
rect 7929 16167 7987 16173
rect 7760 16136 7880 16164
rect 4617 16127 4675 16133
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 2648 16068 3985 16096
rect 2648 16056 2654 16068
rect 3973 16065 3985 16068
rect 4019 16065 4031 16099
rect 3973 16059 4031 16065
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 4080 15960 4108 16059
rect 4154 16056 4160 16108
rect 4212 16096 4218 16108
rect 4341 16099 4399 16105
rect 4212 16068 4257 16096
rect 4212 16056 4218 16068
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16096 4859 16099
rect 4847 16068 7420 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 4356 16028 4384 16059
rect 4356 16000 5028 16028
rect 4338 15960 4344 15972
rect 4080 15932 4344 15960
rect 4338 15920 4344 15932
rect 4396 15920 4402 15972
rect 3694 15892 3700 15904
rect 3655 15864 3700 15892
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 5000 15901 5028 16000
rect 7392 15960 7420 16068
rect 7466 16056 7472 16108
rect 7524 16096 7530 16108
rect 7852 16105 7880 16136
rect 7929 16133 7941 16167
rect 7975 16164 7987 16167
rect 8018 16164 8024 16176
rect 7975 16136 8024 16164
rect 7975 16133 7987 16136
rect 7929 16127 7987 16133
rect 8018 16124 8024 16136
rect 8076 16124 8082 16176
rect 8478 16124 8484 16176
rect 8536 16164 8542 16176
rect 9125 16167 9183 16173
rect 9125 16164 9137 16167
rect 8536 16136 9137 16164
rect 8536 16124 8542 16136
rect 9125 16133 9137 16136
rect 9171 16133 9183 16167
rect 9125 16127 9183 16133
rect 7721 16099 7779 16105
rect 7721 16096 7733 16099
rect 7524 16068 7733 16096
rect 7524 16056 7530 16068
rect 7721 16065 7733 16068
rect 7767 16065 7779 16099
rect 7721 16059 7779 16065
rect 7829 16099 7887 16105
rect 7829 16065 7841 16099
rect 7875 16065 7887 16099
rect 7829 16059 7887 16065
rect 8113 16099 8171 16105
rect 8113 16065 8125 16099
rect 8159 16096 8171 16099
rect 9306 16096 9312 16108
rect 8159 16068 9312 16096
rect 8159 16065 8171 16068
rect 8113 16059 8171 16065
rect 7650 15960 7656 15972
rect 7392 15932 7656 15960
rect 7650 15920 7656 15932
rect 7708 15960 7714 15972
rect 8128 15960 8156 16059
rect 9306 16056 9312 16068
rect 9364 16096 9370 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 9364 16068 9413 16096
rect 9364 16056 9370 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 9217 16031 9275 16037
rect 9217 16028 9229 16031
rect 8260 16000 9229 16028
rect 8260 15988 8266 16000
rect 9217 15997 9229 16000
rect 9263 16028 9275 16031
rect 9508 16028 9536 16204
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 19150 16192 19156 16244
rect 19208 16232 19214 16244
rect 20990 16232 20996 16244
rect 19208 16204 20996 16232
rect 19208 16192 19214 16204
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 22094 16232 22100 16244
rect 22055 16204 22100 16232
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 25225 16235 25283 16241
rect 25225 16201 25237 16235
rect 25271 16232 25283 16235
rect 25958 16232 25964 16244
rect 25271 16204 25964 16232
rect 25271 16201 25283 16204
rect 25225 16195 25283 16201
rect 25958 16192 25964 16204
rect 26016 16232 26022 16244
rect 27525 16235 27583 16241
rect 27525 16232 27537 16235
rect 26016 16204 27537 16232
rect 26016 16192 26022 16204
rect 27525 16201 27537 16204
rect 27571 16201 27583 16235
rect 27525 16195 27583 16201
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 11974 16164 11980 16176
rect 9732 16136 11980 16164
rect 9732 16124 9738 16136
rect 11974 16124 11980 16136
rect 12032 16124 12038 16176
rect 12342 16124 12348 16176
rect 12400 16124 12406 16176
rect 15381 16167 15439 16173
rect 15381 16133 15393 16167
rect 15427 16164 15439 16167
rect 15746 16164 15752 16176
rect 15427 16136 15752 16164
rect 15427 16133 15439 16136
rect 15381 16127 15439 16133
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 18690 16124 18696 16176
rect 18748 16164 18754 16176
rect 27246 16164 27252 16176
rect 18748 16136 27252 16164
rect 18748 16124 18754 16136
rect 27246 16124 27252 16136
rect 27304 16124 27310 16176
rect 10042 16096 10048 16108
rect 10003 16068 10048 16096
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 15194 16096 15200 16108
rect 14884 16068 15200 16096
rect 14884 16056 14890 16068
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 20530 16056 20536 16108
rect 20588 16096 20594 16108
rect 21913 16099 21971 16105
rect 21913 16096 21925 16099
rect 20588 16068 21925 16096
rect 20588 16056 20594 16068
rect 21913 16065 21925 16068
rect 21959 16065 21971 16099
rect 21913 16059 21971 16065
rect 25041 16099 25099 16105
rect 25041 16065 25053 16099
rect 25087 16096 25099 16099
rect 25498 16096 25504 16108
rect 25087 16068 25504 16096
rect 25087 16065 25099 16068
rect 25041 16059 25099 16065
rect 25498 16056 25504 16068
rect 25556 16056 25562 16108
rect 26513 16099 26571 16105
rect 26513 16065 26525 16099
rect 26559 16096 26571 16099
rect 27617 16099 27675 16105
rect 26559 16068 27200 16096
rect 26559 16065 26571 16068
rect 26513 16059 26571 16065
rect 9263 16000 9536 16028
rect 9263 15997 9275 16000
rect 9217 15991 9275 15997
rect 9950 15988 9956 16040
rect 10008 16028 10014 16040
rect 10413 16031 10471 16037
rect 10413 16028 10425 16031
rect 10008 16000 10425 16028
rect 10008 15988 10014 16000
rect 10413 15997 10425 16000
rect 10459 16028 10471 16031
rect 11054 16028 11060 16040
rect 10459 16000 11060 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 11606 16028 11612 16040
rect 11567 16000 11612 16028
rect 11606 15988 11612 16000
rect 11664 15988 11670 16040
rect 11882 16028 11888 16040
rect 11843 16000 11888 16028
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 13357 16031 13415 16037
rect 13357 16028 13369 16031
rect 12400 16000 13369 16028
rect 12400 15988 12406 16000
rect 13357 15997 13369 16000
rect 13403 15997 13415 16031
rect 13357 15991 13415 15997
rect 7708 15932 8156 15960
rect 9585 15963 9643 15969
rect 7708 15920 7714 15932
rect 9585 15929 9597 15963
rect 9631 15960 9643 15963
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 9631 15932 10517 15960
rect 9631 15929 9643 15932
rect 9585 15923 9643 15929
rect 10505 15929 10517 15932
rect 10551 15960 10563 15963
rect 10965 15963 11023 15969
rect 10551 15932 10824 15960
rect 10551 15929 10563 15932
rect 10505 15923 10563 15929
rect 4985 15895 5043 15901
rect 4985 15861 4997 15895
rect 5031 15892 5043 15895
rect 5166 15892 5172 15904
rect 5031 15864 5172 15892
rect 5031 15861 5043 15864
rect 4985 15855 5043 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5258 15852 5264 15904
rect 5316 15892 5322 15904
rect 7561 15895 7619 15901
rect 5316 15864 5361 15892
rect 5316 15852 5322 15864
rect 7561 15861 7573 15895
rect 7607 15892 7619 15895
rect 7834 15892 7840 15904
rect 7607 15864 7840 15892
rect 7607 15861 7619 15864
rect 7561 15855 7619 15861
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 9122 15892 9128 15904
rect 9083 15864 9128 15892
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 10594 15892 10600 15904
rect 10555 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 10796 15892 10824 15932
rect 10965 15929 10977 15963
rect 11011 15960 11023 15963
rect 11238 15960 11244 15972
rect 11011 15932 11244 15960
rect 11011 15929 11023 15932
rect 10965 15923 11023 15929
rect 11238 15920 11244 15932
rect 11296 15920 11302 15972
rect 27172 15969 27200 16068
rect 27617 16065 27629 16099
rect 27663 16096 27675 16099
rect 28166 16096 28172 16108
rect 27663 16068 28172 16096
rect 27663 16065 27675 16068
rect 27617 16059 27675 16065
rect 28166 16056 28172 16068
rect 28224 16056 28230 16108
rect 27246 15988 27252 16040
rect 27304 16028 27310 16040
rect 27709 16031 27767 16037
rect 27709 16028 27721 16031
rect 27304 16000 27721 16028
rect 27304 15988 27310 16000
rect 27709 15997 27721 16000
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 27157 15963 27215 15969
rect 27157 15929 27169 15963
rect 27203 15929 27215 15963
rect 27157 15923 27215 15929
rect 12434 15892 12440 15904
rect 10796 15864 12440 15892
rect 12434 15852 12440 15864
rect 12492 15852 12498 15904
rect 18049 15895 18107 15901
rect 18049 15861 18061 15895
rect 18095 15892 18107 15895
rect 18138 15892 18144 15904
rect 18095 15864 18144 15892
rect 18095 15861 18107 15864
rect 18049 15855 18107 15861
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 26697 15895 26755 15901
rect 26697 15861 26709 15895
rect 26743 15892 26755 15895
rect 26878 15892 26884 15904
rect 26743 15864 26884 15892
rect 26743 15861 26755 15864
rect 26697 15855 26755 15861
rect 26878 15852 26884 15864
rect 26936 15852 26942 15904
rect 1104 15802 28888 15824
rect 1104 15750 3350 15802
rect 3402 15750 3414 15802
rect 3466 15750 3478 15802
rect 3530 15750 3542 15802
rect 3594 15750 3606 15802
rect 3658 15750 8150 15802
rect 8202 15750 8214 15802
rect 8266 15750 8278 15802
rect 8330 15750 8342 15802
rect 8394 15750 8406 15802
rect 8458 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 17750 15802
rect 17802 15750 17814 15802
rect 17866 15750 17878 15802
rect 17930 15750 17942 15802
rect 17994 15750 18006 15802
rect 18058 15750 22550 15802
rect 22602 15750 22614 15802
rect 22666 15750 22678 15802
rect 22730 15750 22742 15802
rect 22794 15750 22806 15802
rect 22858 15750 27350 15802
rect 27402 15750 27414 15802
rect 27466 15750 27478 15802
rect 27530 15750 27542 15802
rect 27594 15750 27606 15802
rect 27658 15750 28888 15802
rect 1104 15728 28888 15750
rect 1765 15691 1823 15697
rect 1765 15657 1777 15691
rect 1811 15688 1823 15691
rect 2590 15688 2596 15700
rect 1811 15660 2596 15688
rect 1811 15657 1823 15660
rect 1765 15651 1823 15657
rect 2590 15648 2596 15660
rect 2648 15648 2654 15700
rect 3255 15691 3313 15697
rect 3255 15657 3267 15691
rect 3301 15688 3313 15691
rect 3694 15688 3700 15700
rect 3301 15660 3700 15688
rect 3301 15657 3313 15660
rect 3255 15651 3313 15657
rect 3694 15648 3700 15660
rect 3752 15648 3758 15700
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 5258 15688 5264 15700
rect 4212 15660 5264 15688
rect 4212 15648 4218 15660
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 8628 15660 9137 15688
rect 8628 15648 8634 15660
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9125 15651 9183 15657
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 11146 15688 11152 15700
rect 10652 15660 11152 15688
rect 10652 15648 10658 15660
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11606 15648 11612 15700
rect 11664 15688 11670 15700
rect 11701 15691 11759 15697
rect 11701 15688 11713 15691
rect 11664 15660 11713 15688
rect 11664 15648 11670 15660
rect 11701 15657 11713 15660
rect 11747 15688 11759 15691
rect 11747 15660 12434 15688
rect 11747 15657 11759 15660
rect 11701 15651 11759 15657
rect 3234 15512 3240 15564
rect 3292 15552 3298 15564
rect 3513 15555 3571 15561
rect 3513 15552 3525 15555
rect 3292 15524 3525 15552
rect 3292 15512 3298 15524
rect 3513 15521 3525 15524
rect 3559 15552 3571 15555
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 3559 15524 5273 15552
rect 3559 15521 3571 15524
rect 3513 15515 3571 15521
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 12406 15552 12434 15660
rect 19426 15648 19432 15700
rect 19484 15688 19490 15700
rect 20349 15691 20407 15697
rect 20349 15688 20361 15691
rect 19484 15660 20361 15688
rect 19484 15648 19490 15660
rect 20349 15657 20361 15660
rect 20395 15657 20407 15691
rect 20530 15688 20536 15700
rect 20491 15660 20536 15688
rect 20349 15651 20407 15657
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 28166 15648 28172 15700
rect 28224 15688 28230 15700
rect 28353 15691 28411 15697
rect 28353 15688 28365 15691
rect 28224 15660 28365 15688
rect 28224 15648 28230 15660
rect 28353 15657 28365 15660
rect 28399 15657 28411 15691
rect 28353 15651 28411 15657
rect 19334 15620 19340 15632
rect 19247 15592 19340 15620
rect 19334 15580 19340 15592
rect 19392 15620 19398 15632
rect 19981 15623 20039 15629
rect 19981 15620 19993 15623
rect 19392 15592 19993 15620
rect 19392 15580 19398 15592
rect 19981 15589 19993 15592
rect 20027 15620 20039 15623
rect 20070 15620 20076 15632
rect 20027 15592 20076 15620
rect 20027 15589 20039 15592
rect 19981 15583 20039 15589
rect 20070 15580 20076 15592
rect 20128 15580 20134 15632
rect 24489 15623 24547 15629
rect 24489 15589 24501 15623
rect 24535 15620 24547 15623
rect 24854 15620 24860 15632
rect 24535 15592 24860 15620
rect 24535 15589 24547 15592
rect 24489 15583 24547 15589
rect 24854 15580 24860 15592
rect 24912 15580 24918 15632
rect 15102 15552 15108 15564
rect 12406 15524 15108 15552
rect 5261 15515 5319 15521
rect 15102 15512 15108 15524
rect 15160 15512 15166 15564
rect 19794 15552 19800 15564
rect 19536 15524 19800 15552
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 7055 15456 7389 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 7377 15453 7389 15456
rect 7423 15484 7435 15487
rect 7423 15456 10456 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 2682 15376 2688 15428
rect 2740 15376 2746 15428
rect 10428 15425 10456 15456
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 19536 15493 19564 15524
rect 19794 15512 19800 15524
rect 19852 15552 19858 15564
rect 21542 15552 21548 15564
rect 19852 15524 21548 15552
rect 19852 15512 19858 15524
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 22557 15555 22615 15561
rect 22557 15521 22569 15555
rect 22603 15552 22615 15555
rect 26326 15552 26332 15564
rect 22603 15524 26332 15552
rect 22603 15521 22615 15524
rect 22557 15515 22615 15521
rect 26326 15512 26332 15524
rect 26384 15512 26390 15564
rect 26878 15552 26884 15564
rect 26839 15524 26884 15552
rect 26878 15512 26884 15524
rect 26936 15512 26942 15564
rect 19521 15487 19579 15493
rect 11112 15456 12112 15484
rect 11112 15444 11118 15456
rect 12084 15428 12112 15456
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15484 19763 15487
rect 21450 15484 21456 15496
rect 19751 15456 21456 15484
rect 19751 15453 19763 15456
rect 19705 15447 19763 15453
rect 21450 15444 21456 15456
rect 21508 15444 21514 15496
rect 24946 15484 24952 15496
rect 24886 15470 24952 15484
rect 24872 15456 24952 15470
rect 9401 15419 9459 15425
rect 9401 15385 9413 15419
rect 9447 15416 9459 15419
rect 10413 15419 10471 15425
rect 9447 15388 9481 15416
rect 9447 15385 9459 15388
rect 9401 15379 9459 15385
rect 10413 15385 10425 15419
rect 10459 15416 10471 15419
rect 10459 15388 11836 15416
rect 10459 15385 10471 15388
rect 10413 15379 10471 15385
rect 8665 15351 8723 15357
rect 8665 15317 8677 15351
rect 8711 15348 8723 15351
rect 9416 15348 9444 15379
rect 9766 15348 9772 15360
rect 8711 15320 9772 15348
rect 8711 15317 8723 15320
rect 8665 15311 8723 15317
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 11808 15348 11836 15388
rect 12066 15376 12072 15428
rect 12124 15416 12130 15428
rect 15746 15416 15752 15428
rect 12124 15388 15752 15416
rect 12124 15376 12130 15388
rect 15746 15376 15752 15388
rect 15804 15376 15810 15428
rect 20806 15416 20812 15428
rect 20767 15388 20812 15416
rect 20806 15376 20812 15388
rect 20864 15376 20870 15428
rect 12529 15351 12587 15357
rect 12529 15348 12541 15351
rect 11808 15320 12541 15348
rect 12529 15317 12541 15320
rect 12575 15348 12587 15351
rect 15930 15348 15936 15360
rect 12575 15320 15936 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 20349 15351 20407 15357
rect 20349 15317 20361 15351
rect 20395 15348 20407 15351
rect 21910 15348 21916 15360
rect 20395 15320 21916 15348
rect 20395 15317 20407 15320
rect 20349 15311 20407 15317
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 24872 15348 24900 15456
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 26237 15487 26295 15493
rect 26237 15453 26249 15487
rect 26283 15484 26295 15487
rect 26602 15484 26608 15496
rect 26283 15456 26608 15484
rect 26283 15453 26295 15456
rect 26237 15447 26295 15453
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 27890 15444 27896 15496
rect 27948 15484 27954 15496
rect 27948 15470 28014 15484
rect 27948 15456 28028 15470
rect 27948 15444 27954 15456
rect 25958 15416 25964 15428
rect 25919 15388 25964 15416
rect 25958 15376 25964 15388
rect 26016 15376 26022 15428
rect 25314 15348 25320 15360
rect 24872 15320 25320 15348
rect 25314 15308 25320 15320
rect 25372 15348 25378 15360
rect 28000 15348 28028 15456
rect 25372 15320 28028 15348
rect 25372 15308 25378 15320
rect 1104 15258 28888 15280
rect 1104 15206 5750 15258
rect 5802 15206 5814 15258
rect 5866 15206 5878 15258
rect 5930 15206 5942 15258
rect 5994 15206 6006 15258
rect 6058 15206 10550 15258
rect 10602 15206 10614 15258
rect 10666 15206 10678 15258
rect 10730 15206 10742 15258
rect 10794 15206 10806 15258
rect 10858 15206 15350 15258
rect 15402 15206 15414 15258
rect 15466 15206 15478 15258
rect 15530 15206 15542 15258
rect 15594 15206 15606 15258
rect 15658 15206 20150 15258
rect 20202 15206 20214 15258
rect 20266 15206 20278 15258
rect 20330 15206 20342 15258
rect 20394 15206 20406 15258
rect 20458 15206 24950 15258
rect 25002 15206 25014 15258
rect 25066 15206 25078 15258
rect 25130 15206 25142 15258
rect 25194 15206 25206 15258
rect 25258 15206 28888 15258
rect 1104 15184 28888 15206
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 11606 15144 11612 15156
rect 7616 15116 11612 15144
rect 7616 15104 7622 15116
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 12158 15144 12164 15156
rect 11808 15116 12164 15144
rect 3970 15036 3976 15088
rect 4028 15036 4034 15088
rect 5626 15076 5632 15088
rect 5587 15048 5632 15076
rect 5626 15036 5632 15048
rect 5684 15036 5690 15088
rect 7834 15076 7840 15088
rect 7795 15048 7840 15076
rect 7834 15036 7840 15048
rect 7892 15036 7898 15088
rect 8570 15036 8576 15088
rect 8628 15036 8634 15088
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11808 15076 11836 15116
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 17586 15104 17592 15156
rect 17644 15144 17650 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 17644 15116 18797 15144
rect 17644 15104 17650 15116
rect 18785 15113 18797 15116
rect 18831 15144 18843 15147
rect 20717 15147 20775 15153
rect 18831 15116 19472 15144
rect 18831 15113 18843 15116
rect 18785 15107 18843 15113
rect 11204 15048 11836 15076
rect 11885 15079 11943 15085
rect 11204 15036 11210 15048
rect 11885 15045 11897 15079
rect 11931 15076 11943 15079
rect 12066 15076 12072 15088
rect 11931 15048 12072 15076
rect 11931 15045 11943 15048
rect 11885 15039 11943 15045
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 3142 15008 3148 15020
rect 3103 14980 3148 15008
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 5810 15008 5816 15020
rect 5771 14980 5816 15008
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 14977 7067 15011
rect 7558 15008 7564 15020
rect 7519 14980 7564 15008
rect 7009 14971 7067 14977
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14940 3479 14943
rect 3878 14940 3884 14952
rect 3467 14912 3884 14940
rect 3467 14909 3479 14912
rect 3421 14903 3479 14909
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 6840 14940 6868 14971
rect 4908 14912 6868 14940
rect 7024 14940 7052 14971
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11296 14980 11805 15008
rect 11296 14968 11302 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11974 15008 11980 15020
rect 11935 14980 11980 15008
rect 11793 14971 11851 14977
rect 7466 14940 7472 14952
rect 7024 14912 7472 14940
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 4154 14804 4160 14816
rect 2648 14776 4160 14804
rect 2648 14764 2654 14776
rect 4154 14764 4160 14776
rect 4212 14804 4218 14816
rect 4908 14813 4936 14912
rect 7466 14900 7472 14912
rect 7524 14940 7530 14952
rect 9122 14940 9128 14952
rect 7524 14912 9128 14940
rect 7524 14900 7530 14912
rect 9122 14900 9128 14912
rect 9180 14940 9186 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 9180 14912 9321 14940
rect 9180 14900 9186 14912
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 11808 14940 11836 14971
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12176 15017 12204 15104
rect 18601 15079 18659 15085
rect 18601 15045 18613 15079
rect 18647 15076 18659 15079
rect 19153 15079 19211 15085
rect 19153 15076 19165 15079
rect 18647 15048 19165 15076
rect 18647 15045 18659 15048
rect 18601 15039 18659 15045
rect 19153 15045 19165 15048
rect 19199 15045 19211 15079
rect 19153 15039 19211 15045
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 14977 12219 15011
rect 12434 15008 12440 15020
rect 12395 14980 12440 15008
rect 12161 14971 12219 14977
rect 12176 14940 12204 14971
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 18877 15011 18935 15017
rect 18877 14977 18889 15011
rect 18923 15008 18935 15011
rect 19334 15008 19340 15020
rect 18923 14980 19340 15008
rect 18923 14977 18935 14980
rect 18877 14971 18935 14977
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 19444 15017 19472 15116
rect 20717 15113 20729 15147
rect 20763 15144 20775 15147
rect 20806 15144 20812 15156
rect 20763 15116 20812 15144
rect 20763 15113 20775 15116
rect 20717 15107 20775 15113
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 21910 15144 21916 15156
rect 21871 15116 21916 15144
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 24854 15104 24860 15156
rect 24912 15144 24918 15156
rect 25041 15147 25099 15153
rect 25041 15144 25053 15147
rect 24912 15116 25053 15144
rect 24912 15104 24918 15116
rect 25041 15113 25053 15116
rect 25087 15113 25099 15147
rect 25498 15144 25504 15156
rect 25459 15116 25504 15144
rect 25041 15107 25099 15113
rect 25498 15104 25504 15116
rect 25556 15104 25562 15156
rect 22278 15076 22284 15088
rect 22191 15048 22284 15076
rect 22278 15036 22284 15048
rect 22336 15076 22342 15088
rect 22336 15048 24256 15076
rect 22336 15036 22342 15048
rect 24228 15020 24256 15048
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 15008 19487 15011
rect 20714 15008 20720 15020
rect 19475 14980 20720 15008
rect 19475 14977 19487 14980
rect 19429 14971 19487 14977
rect 20714 14968 20720 14980
rect 20772 15008 20778 15020
rect 21266 15008 21272 15020
rect 20772 14980 21272 15008
rect 20772 14968 20778 14980
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22186 15008 22192 15020
rect 22143 14980 22192 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22186 14968 22192 14980
rect 22244 14968 22250 15020
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 12529 14943 12587 14949
rect 12529 14940 12541 14943
rect 11808 14912 12020 14940
rect 12176 14912 12541 14940
rect 9309 14903 9367 14909
rect 11609 14875 11667 14881
rect 11609 14841 11621 14875
rect 11655 14872 11667 14875
rect 11882 14872 11888 14884
rect 11655 14844 11888 14872
rect 11655 14841 11667 14844
rect 11609 14835 11667 14841
rect 11882 14832 11888 14844
rect 11940 14832 11946 14884
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 4212 14776 4905 14804
rect 4212 14764 4218 14776
rect 4893 14773 4905 14776
rect 4939 14773 4951 14807
rect 4893 14767 4951 14773
rect 5997 14807 6055 14813
rect 5997 14773 6009 14807
rect 6043 14804 6055 14807
rect 6546 14804 6552 14816
rect 6043 14776 6552 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 7193 14807 7251 14813
rect 7193 14773 7205 14807
rect 7239 14804 7251 14807
rect 8478 14804 8484 14816
rect 7239 14776 8484 14804
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 11992 14804 12020 14912
rect 12529 14909 12541 14912
rect 12575 14909 12587 14943
rect 19150 14940 19156 14952
rect 19111 14912 19156 14940
rect 12529 14903 12587 14909
rect 19150 14900 19156 14912
rect 19208 14900 19214 14952
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 22388 14940 22416 14971
rect 24210 14968 24216 15020
rect 24268 15008 24274 15020
rect 25133 15011 25191 15017
rect 25133 15008 25145 15011
rect 24268 14980 25145 15008
rect 24268 14968 24274 14980
rect 25133 14977 25145 14980
rect 25179 14977 25191 15011
rect 25133 14971 25191 14977
rect 21968 14912 22416 14940
rect 21968 14900 21974 14912
rect 24118 14900 24124 14952
rect 24176 14940 24182 14952
rect 24857 14943 24915 14949
rect 24857 14940 24869 14943
rect 24176 14912 24869 14940
rect 24176 14900 24182 14912
rect 17129 14875 17187 14881
rect 17129 14841 17141 14875
rect 17175 14872 17187 14875
rect 17218 14872 17224 14884
rect 17175 14844 17224 14872
rect 17175 14841 17187 14844
rect 17129 14835 17187 14841
rect 17218 14832 17224 14844
rect 17276 14872 17282 14884
rect 19702 14872 19708 14884
rect 17276 14844 19708 14872
rect 17276 14832 17282 14844
rect 19702 14832 19708 14844
rect 19760 14872 19766 14884
rect 23106 14872 23112 14884
rect 19760 14844 23112 14872
rect 19760 14832 19766 14844
rect 23106 14832 23112 14844
rect 23164 14832 23170 14884
rect 24412 14816 24440 14912
rect 24857 14909 24869 14912
rect 24903 14909 24915 14943
rect 24857 14903 24915 14909
rect 12342 14804 12348 14816
rect 11992 14776 12348 14804
rect 12342 14764 12348 14776
rect 12400 14804 12406 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12400 14776 12449 14804
rect 12400 14764 12406 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 12805 14807 12863 14813
rect 12805 14773 12817 14807
rect 12851 14804 12863 14807
rect 15746 14804 15752 14816
rect 12851 14776 15752 14804
rect 12851 14773 12863 14776
rect 12805 14767 12863 14773
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 18601 14807 18659 14813
rect 18601 14804 18613 14807
rect 18472 14776 18613 14804
rect 18472 14764 18478 14776
rect 18601 14773 18613 14776
rect 18647 14773 18659 14807
rect 24394 14804 24400 14816
rect 24355 14776 24400 14804
rect 18601 14767 18659 14773
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 1104 14714 28888 14736
rect 1104 14662 3350 14714
rect 3402 14662 3414 14714
rect 3466 14662 3478 14714
rect 3530 14662 3542 14714
rect 3594 14662 3606 14714
rect 3658 14662 8150 14714
rect 8202 14662 8214 14714
rect 8266 14662 8278 14714
rect 8330 14662 8342 14714
rect 8394 14662 8406 14714
rect 8458 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 17750 14714
rect 17802 14662 17814 14714
rect 17866 14662 17878 14714
rect 17930 14662 17942 14714
rect 17994 14662 18006 14714
rect 18058 14662 22550 14714
rect 22602 14662 22614 14714
rect 22666 14662 22678 14714
rect 22730 14662 22742 14714
rect 22794 14662 22806 14714
rect 22858 14662 27350 14714
rect 27402 14662 27414 14714
rect 27466 14662 27478 14714
rect 27530 14662 27542 14714
rect 27594 14662 27606 14714
rect 27658 14662 28888 14714
rect 1104 14640 28888 14662
rect 3878 14600 3884 14612
rect 3839 14572 3884 14600
rect 3878 14560 3884 14572
rect 3936 14560 3942 14612
rect 18325 14603 18383 14609
rect 18325 14569 18337 14603
rect 18371 14600 18383 14603
rect 19426 14600 19432 14612
rect 18371 14572 19432 14600
rect 18371 14569 18383 14572
rect 18325 14563 18383 14569
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 21542 14600 21548 14612
rect 21503 14572 21548 14600
rect 21542 14560 21548 14572
rect 21600 14560 21606 14612
rect 4338 14492 4344 14544
rect 4396 14492 4402 14544
rect 21266 14492 21272 14544
rect 21324 14532 21330 14544
rect 21910 14532 21916 14544
rect 21324 14504 21916 14532
rect 21324 14492 21330 14504
rect 21910 14492 21916 14504
rect 21968 14492 21974 14544
rect 4356 14464 4384 14492
rect 8478 14464 8484 14476
rect 4277 14436 4384 14464
rect 4540 14436 8484 14464
rect 4154 14405 4160 14408
rect 4137 14399 4160 14405
rect 4137 14365 4149 14399
rect 4137 14359 4160 14365
rect 4154 14356 4160 14359
rect 4212 14356 4218 14408
rect 4277 14399 4305 14436
rect 4540 14405 4568 14436
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 14921 14467 14979 14473
rect 14921 14464 14933 14467
rect 12308 14436 14933 14464
rect 12308 14424 12314 14436
rect 14921 14433 14933 14436
rect 14967 14464 14979 14467
rect 16206 14464 16212 14476
rect 14967 14436 16212 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 17405 14467 17463 14473
rect 17405 14464 17417 14467
rect 16868 14436 17417 14464
rect 4262 14393 4320 14399
rect 4262 14359 4274 14393
rect 4308 14359 4320 14393
rect 4262 14353 4320 14359
rect 4362 14396 4420 14402
rect 4362 14362 4374 14396
rect 4408 14362 4420 14396
rect 4362 14356 4420 14362
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 5166 14396 5172 14408
rect 5127 14368 5172 14396
rect 4525 14359 4583 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6328 14368 6469 14396
rect 6328 14356 6334 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 4377 14328 4405 14356
rect 5258 14328 5264 14340
rect 4377 14300 5264 14328
rect 4816 14272 4844 14300
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 5353 14331 5411 14337
rect 5353 14297 5365 14331
rect 5399 14328 5411 14331
rect 5810 14328 5816 14340
rect 5399 14300 5816 14328
rect 5399 14297 5411 14300
rect 5353 14291 5411 14297
rect 5810 14288 5816 14300
rect 5868 14328 5874 14340
rect 6638 14328 6644 14340
rect 5868 14300 6644 14328
rect 5868 14288 5874 14300
rect 6638 14288 6644 14300
rect 6696 14288 6702 14340
rect 6825 14331 6883 14337
rect 6825 14297 6837 14331
rect 6871 14328 6883 14331
rect 7098 14328 7104 14340
rect 6871 14300 7104 14328
rect 6871 14297 6883 14300
rect 6825 14291 6883 14297
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 15102 14288 15108 14340
rect 15160 14328 15166 14340
rect 15197 14331 15255 14337
rect 15197 14328 15209 14331
rect 15160 14300 15209 14328
rect 15160 14288 15166 14300
rect 15197 14297 15209 14300
rect 15243 14297 15255 14331
rect 16574 14328 16580 14340
rect 16422 14300 16580 14328
rect 15197 14291 15255 14297
rect 16574 14288 16580 14300
rect 16632 14328 16638 14340
rect 16868 14328 16896 14436
rect 17405 14433 17417 14436
rect 17451 14433 17463 14467
rect 22278 14464 22284 14476
rect 17405 14427 17463 14433
rect 21744 14436 22284 14464
rect 17218 14396 17224 14408
rect 17179 14368 17224 14396
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 21744 14405 21772 14436
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 17552 14368 18153 14396
rect 17552 14356 17558 14368
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 21729 14399 21787 14405
rect 21729 14365 21741 14399
rect 21775 14365 21787 14399
rect 21729 14359 21787 14365
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 22186 14396 22192 14408
rect 21867 14368 22192 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 22186 14356 22192 14368
rect 22244 14356 22250 14408
rect 16632 14300 16896 14328
rect 16632 14288 16638 14300
rect 16942 14288 16948 14340
rect 17000 14328 17006 14340
rect 17957 14331 18015 14337
rect 17000 14300 17045 14328
rect 17000 14288 17006 14300
rect 17957 14297 17969 14331
rect 18003 14297 18015 14331
rect 22094 14328 22100 14340
rect 22055 14300 22100 14328
rect 17957 14291 18015 14297
rect 4798 14260 4804 14272
rect 4759 14232 4804 14260
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 16666 14220 16672 14272
rect 16724 14260 16730 14272
rect 17972 14260 18000 14291
rect 22094 14288 22100 14300
rect 22152 14288 22158 14340
rect 16724 14232 18000 14260
rect 16724 14220 16730 14232
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 21913 14263 21971 14269
rect 21913 14260 21925 14263
rect 21876 14232 21925 14260
rect 21876 14220 21882 14232
rect 21913 14229 21925 14232
rect 21959 14229 21971 14263
rect 21913 14223 21971 14229
rect 1104 14170 28888 14192
rect 1104 14118 5750 14170
rect 5802 14118 5814 14170
rect 5866 14118 5878 14170
rect 5930 14118 5942 14170
rect 5994 14118 6006 14170
rect 6058 14118 10550 14170
rect 10602 14118 10614 14170
rect 10666 14118 10678 14170
rect 10730 14118 10742 14170
rect 10794 14118 10806 14170
rect 10858 14118 15350 14170
rect 15402 14118 15414 14170
rect 15466 14118 15478 14170
rect 15530 14118 15542 14170
rect 15594 14118 15606 14170
rect 15658 14118 20150 14170
rect 20202 14118 20214 14170
rect 20266 14118 20278 14170
rect 20330 14118 20342 14170
rect 20394 14118 20406 14170
rect 20458 14118 24950 14170
rect 25002 14118 25014 14170
rect 25066 14118 25078 14170
rect 25130 14118 25142 14170
rect 25194 14118 25206 14170
rect 25258 14118 28888 14170
rect 1104 14096 28888 14118
rect 15746 14056 15752 14068
rect 15396 14028 15752 14056
rect 6546 13988 6552 14000
rect 6507 13960 6552 13988
rect 6546 13948 6552 13960
rect 6604 13948 6610 14000
rect 15396 13988 15424 14028
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 21446 14059 21504 14065
rect 21446 14025 21458 14059
rect 21492 14056 21504 14059
rect 24210 14056 24216 14068
rect 21492 14028 22784 14056
rect 24171 14028 24216 14056
rect 21492 14025 21504 14028
rect 21446 14019 21504 14025
rect 16666 13988 16672 14000
rect 15304 13960 15424 13988
rect 15580 13960 16672 13988
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13920 12771 13923
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12759 13892 13093 13920
rect 12759 13889 12771 13892
rect 12713 13883 12771 13889
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 13538 13920 13544 13932
rect 13499 13892 13544 13920
rect 13081 13883 13139 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14090 13920 14096 13932
rect 14051 13892 14096 13920
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 15304 13929 15332 13960
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 15378 13880 15384 13932
rect 15436 13920 15442 13932
rect 15580 13929 15608 13960
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 18414 13988 18420 14000
rect 18375 13960 18420 13988
rect 18414 13948 18420 13960
rect 18472 13948 18478 14000
rect 22756 13997 22784 14028
rect 24210 14016 24216 14028
rect 24268 14016 24274 14068
rect 21545 13991 21603 13997
rect 21545 13957 21557 13991
rect 21591 13988 21603 13991
rect 21913 13991 21971 13997
rect 21913 13988 21925 13991
rect 21591 13960 21925 13988
rect 21591 13957 21603 13960
rect 21545 13951 21603 13957
rect 21913 13957 21925 13960
rect 21959 13957 21971 13991
rect 21913 13951 21971 13957
rect 22741 13991 22799 13997
rect 22741 13957 22753 13991
rect 22787 13957 22799 13991
rect 24949 13991 25007 13997
rect 24949 13988 24961 13991
rect 23966 13960 24961 13988
rect 22741 13951 22799 13957
rect 24949 13957 24961 13960
rect 24995 13988 25007 13991
rect 25314 13988 25320 14000
rect 24995 13960 25320 13988
rect 24995 13957 25007 13960
rect 24949 13951 25007 13957
rect 25314 13948 25320 13960
rect 25372 13948 25378 14000
rect 15565 13923 15623 13929
rect 15436 13892 15481 13920
rect 15436 13880 15442 13892
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13889 15715 13923
rect 17313 13923 17371 13929
rect 17313 13920 17325 13923
rect 15657 13883 15715 13889
rect 15856 13892 17325 13920
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 12492 13824 13921 13852
rect 12492 13812 12498 13824
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 15672 13852 15700 13883
rect 15746 13852 15752 13864
rect 13909 13815 13967 13821
rect 14936 13824 15752 13852
rect 6730 13784 6736 13796
rect 6691 13756 6736 13784
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 14182 13744 14188 13796
rect 14240 13784 14246 13796
rect 14936 13784 14964 13824
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 15102 13784 15108 13796
rect 14240 13756 14964 13784
rect 15063 13756 15108 13784
rect 14240 13744 14246 13756
rect 15102 13744 15108 13756
rect 15160 13744 15166 13796
rect 15856 13784 15884 13892
rect 17313 13889 17325 13892
rect 17359 13889 17371 13923
rect 17494 13920 17500 13932
rect 17455 13892 17500 13920
rect 17313 13883 17371 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 20165 13923 20223 13929
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 18141 13855 18199 13861
rect 18141 13852 18153 13855
rect 16264 13824 18153 13852
rect 16264 13812 16270 13824
rect 18141 13821 18153 13824
rect 18187 13821 18199 13855
rect 19536 13852 19564 13906
rect 20165 13889 20177 13923
rect 20211 13920 20223 13923
rect 20714 13920 20720 13932
rect 20211 13892 20720 13920
rect 20211 13889 20223 13892
rect 20165 13883 20223 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 21266 13920 21272 13932
rect 21227 13892 21272 13920
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 21361 13923 21419 13929
rect 21361 13889 21373 13923
rect 21407 13920 21419 13923
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 21407 13918 21496 13920
rect 21560 13918 22201 13920
rect 21407 13892 22201 13918
rect 21407 13889 21419 13892
rect 21468 13890 21588 13892
rect 21361 13883 21419 13889
rect 22189 13889 22201 13892
rect 22235 13920 22247 13923
rect 22278 13920 22284 13932
rect 22235 13892 22284 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 24581 13923 24639 13929
rect 24581 13889 24593 13923
rect 24627 13889 24639 13923
rect 27246 13920 27252 13932
rect 27207 13892 27252 13920
rect 24581 13883 24639 13889
rect 19536 13824 20944 13852
rect 18141 13815 18199 13821
rect 15764 13756 15884 13784
rect 12526 13716 12532 13728
rect 12487 13688 12532 13716
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 15764 13716 15792 13756
rect 14884 13688 15792 13716
rect 20916 13716 20944 13824
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 21913 13855 21971 13861
rect 21048 13844 21588 13852
rect 21652 13844 21772 13852
rect 21913 13844 21925 13855
rect 21048 13824 21925 13844
rect 21048 13812 21054 13824
rect 21560 13816 21680 13824
rect 21744 13821 21925 13824
rect 21959 13821 21971 13855
rect 21744 13816 21971 13821
rect 21913 13815 21971 13816
rect 22002 13812 22008 13864
rect 22060 13852 22066 13864
rect 22465 13855 22523 13861
rect 22465 13852 22477 13855
rect 22060 13824 22477 13852
rect 22060 13812 22066 13824
rect 22465 13821 22477 13824
rect 22511 13821 22523 13855
rect 24596 13852 24624 13883
rect 27246 13880 27252 13892
rect 27304 13880 27310 13932
rect 28166 13920 28172 13932
rect 28127 13892 28172 13920
rect 28166 13880 28172 13892
rect 28224 13880 28230 13932
rect 22465 13815 22523 13821
rect 22572 13824 24624 13852
rect 22572 13784 22600 13824
rect 21836 13756 22600 13784
rect 21174 13716 21180 13728
rect 20916 13688 21180 13716
rect 14884 13676 14890 13688
rect 21174 13676 21180 13688
rect 21232 13716 21238 13728
rect 21836 13716 21864 13756
rect 21232 13688 21864 13716
rect 21232 13676 21238 13688
rect 21910 13676 21916 13728
rect 21968 13716 21974 13728
rect 22097 13719 22155 13725
rect 22097 13716 22109 13719
rect 21968 13688 22109 13716
rect 21968 13676 21974 13688
rect 22097 13685 22109 13688
rect 22143 13685 22155 13719
rect 22097 13679 22155 13685
rect 26878 13676 26884 13728
rect 26936 13716 26942 13728
rect 27065 13719 27123 13725
rect 27065 13716 27077 13719
rect 26936 13688 27077 13716
rect 26936 13676 26942 13688
rect 27065 13685 27077 13688
rect 27111 13685 27123 13719
rect 28350 13716 28356 13728
rect 28311 13688 28356 13716
rect 27065 13679 27123 13685
rect 28350 13676 28356 13688
rect 28408 13676 28414 13728
rect 1104 13626 28888 13648
rect 1104 13574 3350 13626
rect 3402 13574 3414 13626
rect 3466 13574 3478 13626
rect 3530 13574 3542 13626
rect 3594 13574 3606 13626
rect 3658 13574 8150 13626
rect 8202 13574 8214 13626
rect 8266 13574 8278 13626
rect 8330 13574 8342 13626
rect 8394 13574 8406 13626
rect 8458 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 17750 13626
rect 17802 13574 17814 13626
rect 17866 13574 17878 13626
rect 17930 13574 17942 13626
rect 17994 13574 18006 13626
rect 18058 13574 22550 13626
rect 22602 13574 22614 13626
rect 22666 13574 22678 13626
rect 22730 13574 22742 13626
rect 22794 13574 22806 13626
rect 22858 13574 27350 13626
rect 27402 13574 27414 13626
rect 27466 13574 27478 13626
rect 27530 13574 27542 13626
rect 27594 13574 27606 13626
rect 27658 13574 28888 13626
rect 1104 13552 28888 13574
rect 9766 13512 9772 13524
rect 8496 13484 9772 13512
rect 2406 13308 2412 13320
rect 2367 13280 2412 13308
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 4982 13268 4988 13320
rect 5040 13308 5046 13320
rect 8496 13308 8524 13484
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 10781 13515 10839 13521
rect 10781 13481 10793 13515
rect 10827 13512 10839 13515
rect 10962 13512 10968 13524
rect 10827 13484 10968 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 10962 13472 10968 13484
rect 11020 13512 11026 13524
rect 11149 13515 11207 13521
rect 11149 13512 11161 13515
rect 11020 13484 11161 13512
rect 11020 13472 11026 13484
rect 11149 13481 11161 13484
rect 11195 13481 11207 13515
rect 11149 13475 11207 13481
rect 13538 13472 13544 13524
rect 13596 13512 13602 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 13596 13484 13737 13512
rect 13596 13472 13602 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 14148 13484 14657 13512
rect 14148 13472 14154 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 14645 13475 14703 13481
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 15378 13512 15384 13524
rect 14884 13484 14977 13512
rect 15339 13484 15384 13512
rect 14884 13472 14890 13484
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 20530 13512 20536 13524
rect 20443 13484 20536 13512
rect 20530 13472 20536 13484
rect 20588 13512 20594 13524
rect 20806 13512 20812 13524
rect 20588 13484 20812 13512
rect 20588 13472 20594 13484
rect 20806 13472 20812 13484
rect 20864 13472 20870 13524
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 22060 13484 22109 13512
rect 22060 13472 22066 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 14844 13444 14872 13472
rect 15396 13444 15424 13472
rect 17405 13447 17463 13453
rect 17405 13444 17417 13447
rect 12584 13416 14872 13444
rect 14936 13416 15424 13444
rect 16546 13416 17417 13444
rect 12584 13404 12590 13416
rect 8570 13336 8576 13388
rect 8628 13376 8634 13388
rect 13725 13379 13783 13385
rect 8628 13348 13492 13376
rect 8628 13336 8634 13348
rect 8665 13311 8723 13317
rect 8665 13308 8677 13311
rect 5040 13280 8677 13308
rect 5040 13268 5046 13280
rect 8665 13277 8677 13280
rect 8711 13277 8723 13311
rect 9030 13308 9036 13320
rect 8991 13280 9036 13308
rect 8665 13271 8723 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 11164 13317 11192 13348
rect 11149 13311 11207 13317
rect 11149 13277 11161 13311
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 11296 13280 11341 13308
rect 13004 13280 13369 13308
rect 11296 13268 11302 13280
rect 2958 13200 2964 13252
rect 3016 13240 3022 13252
rect 3970 13240 3976 13252
rect 3016 13212 3976 13240
rect 3016 13200 3022 13212
rect 3970 13200 3976 13212
rect 4028 13240 4034 13252
rect 4709 13243 4767 13249
rect 4709 13240 4721 13243
rect 4028 13212 4721 13240
rect 4028 13200 4034 13212
rect 4709 13209 4721 13212
rect 4755 13209 4767 13243
rect 4709 13203 4767 13209
rect 4893 13243 4951 13249
rect 4893 13209 4905 13243
rect 4939 13240 4951 13243
rect 9309 13243 9367 13249
rect 4939 13212 9260 13240
rect 4939 13209 4951 13212
rect 4893 13203 4951 13209
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 2225 13175 2283 13181
rect 2225 13172 2237 13175
rect 1820 13144 2237 13172
rect 1820 13132 1826 13144
rect 2225 13141 2237 13144
rect 2271 13141 2283 13175
rect 5074 13172 5080 13184
rect 5035 13144 5080 13172
rect 2225 13135 2283 13141
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 9232 13172 9260 13212
rect 9309 13209 9321 13243
rect 9355 13240 9367 13243
rect 9582 13240 9588 13252
rect 9355 13212 9588 13240
rect 9355 13209 9367 13212
rect 9309 13203 9367 13209
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 9766 13200 9772 13252
rect 9824 13200 9830 13252
rect 11146 13172 11152 13184
rect 9232 13144 11152 13172
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11517 13175 11575 13181
rect 11517 13141 11529 13175
rect 11563 13172 11575 13175
rect 12250 13172 12256 13184
rect 11563 13144 12256 13172
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12802 13132 12808 13184
rect 12860 13172 12866 13184
rect 13004 13181 13032 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13464 13308 13492 13348
rect 13725 13345 13737 13379
rect 13771 13376 13783 13379
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 13771 13348 14289 13376
rect 13771 13345 13783 13348
rect 13725 13339 13783 13345
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 14182 13308 14188 13320
rect 13464 13280 14188 13308
rect 13357 13271 13415 13277
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13308 14427 13311
rect 14936 13308 14964 13416
rect 15194 13376 15200 13388
rect 14415 13280 14964 13308
rect 15028 13348 15200 13376
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 15028 13249 15056 13348
rect 15194 13336 15200 13348
rect 15252 13376 15258 13388
rect 16546 13376 16574 13416
rect 17405 13413 17417 13416
rect 17451 13444 17463 13447
rect 17586 13444 17592 13456
rect 17451 13416 17592 13444
rect 17451 13413 17463 13416
rect 17405 13407 17463 13413
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 15252 13348 16574 13376
rect 16853 13379 16911 13385
rect 15252 13336 15258 13348
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 16942 13376 16948 13388
rect 16899 13348 16948 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 16942 13336 16948 13348
rect 17000 13376 17006 13388
rect 17310 13376 17316 13388
rect 17000 13348 17316 13376
rect 17000 13336 17006 13348
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 26878 13376 26884 13388
rect 26839 13348 26884 13376
rect 26878 13336 26884 13348
rect 26936 13336 26942 13388
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13308 15531 13311
rect 16666 13308 16672 13320
rect 15519 13280 15976 13308
rect 16579 13280 16672 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 15013 13243 15071 13249
rect 15013 13209 15025 13243
rect 15059 13209 15071 13243
rect 15013 13203 15071 13209
rect 15749 13243 15807 13249
rect 15749 13209 15761 13243
rect 15795 13240 15807 13243
rect 15838 13240 15844 13252
rect 15795 13212 15844 13240
rect 15795 13209 15807 13212
rect 15749 13203 15807 13209
rect 15838 13200 15844 13212
rect 15896 13200 15902 13252
rect 15948 13249 15976 13280
rect 16666 13268 16672 13280
rect 16724 13308 16730 13320
rect 17218 13308 17224 13320
rect 16724 13280 17224 13308
rect 16724 13268 16730 13280
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 20806 13308 20812 13320
rect 20767 13280 20812 13308
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22833 13311 22891 13317
rect 22833 13308 22845 13311
rect 21968 13280 22845 13308
rect 21968 13268 21974 13280
rect 22833 13277 22845 13280
rect 22879 13277 22891 13311
rect 22833 13271 22891 13277
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13308 25007 13311
rect 25406 13308 25412 13320
rect 24995 13280 25412 13308
rect 24995 13277 25007 13280
rect 24949 13271 25007 13277
rect 25406 13268 25412 13280
rect 25464 13268 25470 13320
rect 26602 13308 26608 13320
rect 26563 13280 26608 13308
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 15933 13243 15991 13249
rect 15933 13209 15945 13243
rect 15979 13240 15991 13243
rect 16758 13240 16764 13252
rect 15979 13212 16764 13240
rect 15979 13209 15991 13212
rect 15933 13203 15991 13209
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17405 13243 17463 13249
rect 17405 13240 17417 13243
rect 17092 13212 17417 13240
rect 17092 13200 17098 13212
rect 17405 13209 17417 13212
rect 17451 13209 17463 13243
rect 17405 13203 17463 13209
rect 25314 13200 25320 13252
rect 25372 13240 25378 13252
rect 25372 13212 27370 13240
rect 25372 13200 25378 13212
rect 12989 13175 13047 13181
rect 12989 13172 13001 13175
rect 12860 13144 13001 13172
rect 12860 13132 12866 13144
rect 12989 13141 13001 13144
rect 13035 13141 13047 13175
rect 12989 13135 13047 13141
rect 14813 13175 14871 13181
rect 14813 13141 14825 13175
rect 14859 13172 14871 13175
rect 15194 13172 15200 13184
rect 14859 13144 15200 13172
rect 14859 13141 14871 13144
rect 14813 13135 14871 13141
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 16117 13175 16175 13181
rect 16117 13141 16129 13175
rect 16163 13172 16175 13175
rect 16574 13172 16580 13184
rect 16163 13144 16580 13172
rect 16163 13141 16175 13144
rect 16117 13135 16175 13141
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 16942 13132 16948 13184
rect 17000 13172 17006 13184
rect 23014 13172 23020 13184
rect 17000 13144 17045 13172
rect 22975 13144 23020 13172
rect 17000 13132 17006 13144
rect 23014 13132 23020 13144
rect 23072 13132 23078 13184
rect 25133 13175 25191 13181
rect 25133 13141 25145 13175
rect 25179 13172 25191 13175
rect 25866 13172 25872 13184
rect 25179 13144 25872 13172
rect 25179 13141 25191 13144
rect 25133 13135 25191 13141
rect 25866 13132 25872 13144
rect 25924 13132 25930 13184
rect 27706 13132 27712 13184
rect 27764 13172 27770 13184
rect 28166 13172 28172 13184
rect 27764 13144 28172 13172
rect 27764 13132 27770 13144
rect 28166 13132 28172 13144
rect 28224 13172 28230 13184
rect 28353 13175 28411 13181
rect 28353 13172 28365 13175
rect 28224 13144 28365 13172
rect 28224 13132 28230 13144
rect 28353 13141 28365 13144
rect 28399 13141 28411 13175
rect 28353 13135 28411 13141
rect 1104 13082 28888 13104
rect 1104 13030 5750 13082
rect 5802 13030 5814 13082
rect 5866 13030 5878 13082
rect 5930 13030 5942 13082
rect 5994 13030 6006 13082
rect 6058 13030 10550 13082
rect 10602 13030 10614 13082
rect 10666 13030 10678 13082
rect 10730 13030 10742 13082
rect 10794 13030 10806 13082
rect 10858 13030 15350 13082
rect 15402 13030 15414 13082
rect 15466 13030 15478 13082
rect 15530 13030 15542 13082
rect 15594 13030 15606 13082
rect 15658 13030 20150 13082
rect 20202 13030 20214 13082
rect 20266 13030 20278 13082
rect 20330 13030 20342 13082
rect 20394 13030 20406 13082
rect 20458 13030 24950 13082
rect 25002 13030 25014 13082
rect 25066 13030 25078 13082
rect 25130 13030 25142 13082
rect 25194 13030 25206 13082
rect 25258 13030 28888 13082
rect 1104 13008 28888 13030
rect 8478 12968 8484 12980
rect 8312 12940 8484 12968
rect 1762 12900 1768 12912
rect 1723 12872 1768 12900
rect 1762 12860 1768 12872
rect 1820 12860 1826 12912
rect 3142 12900 3148 12912
rect 2990 12872 3148 12900
rect 3142 12860 3148 12872
rect 3200 12860 3206 12912
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 4798 12900 4804 12912
rect 4028 12872 4108 12900
rect 4028 12860 4034 12872
rect 4080 12841 4108 12872
rect 4377 12872 4804 12900
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 4154 12838 4212 12844
rect 4154 12804 4166 12838
rect 4200 12804 4212 12838
rect 4154 12798 4212 12804
rect 4270 12835 4328 12841
rect 4270 12801 4282 12835
rect 4316 12832 4328 12835
rect 4377 12832 4405 12872
rect 4798 12860 4804 12872
rect 4856 12860 4862 12912
rect 5721 12903 5779 12909
rect 5721 12869 5733 12903
rect 5767 12900 5779 12903
rect 6638 12900 6644 12912
rect 5767 12872 6644 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 6638 12860 6644 12872
rect 6696 12900 6702 12912
rect 8312 12909 8340 12940
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 9582 12968 9588 12980
rect 9543 12940 9588 12968
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 11238 12968 11244 12980
rect 10091 12940 11244 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 12434 12968 12440 12980
rect 11388 12940 12440 12968
rect 11388 12928 11394 12940
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 16758 12968 16764 12980
rect 16719 12940 16764 12968
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 20559 12971 20617 12977
rect 20559 12937 20571 12971
rect 20605 12968 20617 12971
rect 23014 12968 23020 12980
rect 20605 12940 23020 12968
rect 20605 12937 20617 12940
rect 20559 12931 20617 12937
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 27246 12968 27252 12980
rect 27207 12940 27252 12968
rect 27246 12928 27252 12940
rect 27304 12928 27310 12980
rect 27706 12968 27712 12980
rect 27667 12940 27712 12968
rect 27706 12928 27712 12940
rect 27764 12928 27770 12980
rect 8297 12903 8355 12909
rect 6696 12872 7972 12900
rect 6696 12860 6702 12872
rect 4316 12804 4405 12832
rect 4433 12835 4491 12841
rect 4316 12801 4328 12804
rect 1489 12767 1547 12773
rect 1489 12733 1501 12767
rect 1535 12764 1547 12767
rect 1762 12764 1768 12776
rect 1535 12736 1768 12764
rect 1535 12733 1547 12736
rect 1489 12727 1547 12733
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 3234 12628 3240 12640
rect 3195 12600 3240 12628
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 3789 12631 3847 12637
rect 3789 12597 3801 12631
rect 3835 12628 3847 12631
rect 3970 12628 3976 12640
rect 3835 12600 3976 12628
rect 3835 12597 3847 12600
rect 3789 12591 3847 12597
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4172 12628 4200 12798
rect 4270 12795 4328 12801
rect 4433 12801 4445 12835
rect 4479 12832 4491 12835
rect 5074 12832 5080 12844
rect 4479 12804 5080 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 5074 12792 5080 12804
rect 5132 12832 5138 12844
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5132 12804 5549 12832
rect 5132 12792 5138 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12832 5963 12835
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 5951 12804 6837 12832
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 6825 12801 6837 12804
rect 6871 12832 6883 12835
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6871 12804 7297 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7944 12832 7972 12872
rect 8297 12869 8309 12903
rect 8343 12869 8355 12903
rect 8297 12863 8355 12869
rect 10781 12903 10839 12909
rect 10781 12869 10793 12903
rect 10827 12900 10839 12903
rect 12526 12900 12532 12912
rect 10827 12872 12532 12900
rect 10827 12869 10839 12872
rect 10781 12863 10839 12869
rect 12526 12860 12532 12872
rect 12584 12860 12590 12912
rect 20349 12903 20407 12909
rect 20349 12869 20361 12903
rect 20395 12900 20407 12903
rect 20990 12900 20996 12912
rect 20395 12872 20996 12900
rect 20395 12869 20407 12872
rect 20349 12863 20407 12869
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 21361 12903 21419 12909
rect 21361 12869 21373 12903
rect 21407 12900 21419 12903
rect 21818 12900 21824 12912
rect 21407 12872 21824 12900
rect 21407 12869 21419 12872
rect 21361 12863 21419 12869
rect 21818 12860 21824 12872
rect 21876 12860 21882 12912
rect 22065 12903 22123 12909
rect 22065 12900 22077 12903
rect 21928 12872 22077 12900
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 7944 12804 8493 12832
rect 7285 12795 7343 12801
rect 8481 12801 8493 12804
rect 8527 12832 8539 12835
rect 8570 12832 8576 12844
rect 8527 12804 8576 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 8570 12792 8576 12804
rect 8628 12792 8634 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9674 12832 9680 12844
rect 9635 12804 9680 12832
rect 9493 12795 9551 12801
rect 6730 12764 6736 12776
rect 6691 12736 6736 12764
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 9508 12764 9536 12795
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 10239 12835 10297 12841
rect 10239 12801 10251 12835
rect 10285 12832 10297 12835
rect 10962 12832 10968 12844
rect 10285 12804 10968 12832
rect 10285 12801 10297 12804
rect 10239 12795 10297 12801
rect 9858 12764 9864 12776
rect 9508 12736 9864 12764
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 9968 12764 9996 12795
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 12250 12832 12256 12844
rect 12211 12804 12256 12832
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13872 12804 14197 12832
rect 13872 12792 13878 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 17034 12832 17040 12844
rect 16995 12804 17040 12832
rect 14185 12795 14243 12801
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17310 12832 17316 12844
rect 17271 12804 17316 12832
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 21177 12835 21235 12841
rect 21177 12801 21189 12835
rect 21223 12801 21235 12835
rect 21450 12832 21456 12844
rect 21411 12804 21456 12832
rect 21177 12795 21235 12801
rect 15930 12764 15936 12776
rect 9968 12736 10364 12764
rect 15843 12736 15936 12764
rect 4338 12656 4344 12708
rect 4396 12696 4402 12708
rect 9968 12696 9996 12736
rect 4396 12668 9996 12696
rect 10229 12699 10287 12705
rect 4396 12656 4402 12668
rect 10229 12665 10241 12699
rect 10275 12665 10287 12699
rect 10336 12696 10364 12736
rect 15930 12724 15936 12736
rect 15988 12764 15994 12776
rect 16482 12764 16488 12776
rect 15988 12736 16488 12764
rect 15988 12724 15994 12736
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 21192 12764 21220 12795
rect 21450 12792 21456 12804
rect 21508 12832 21514 12844
rect 21928 12832 21956 12872
rect 22065 12869 22077 12872
rect 22111 12869 22123 12903
rect 22278 12900 22284 12912
rect 22239 12872 22284 12900
rect 22065 12863 22123 12869
rect 22278 12860 22284 12872
rect 22336 12860 22342 12912
rect 25314 12860 25320 12912
rect 25372 12860 25378 12912
rect 25866 12900 25872 12912
rect 25827 12872 25872 12900
rect 25866 12860 25872 12872
rect 25924 12900 25930 12912
rect 27617 12903 27675 12909
rect 27617 12900 27629 12903
rect 25924 12872 27629 12900
rect 25924 12860 25930 12872
rect 27617 12869 27629 12872
rect 27663 12869 27675 12903
rect 27617 12863 27675 12869
rect 21508 12804 21956 12832
rect 26145 12835 26203 12841
rect 21508 12792 21514 12804
rect 26145 12801 26157 12835
rect 26191 12832 26203 12835
rect 26602 12832 26608 12844
rect 26191 12804 26608 12832
rect 26191 12801 26203 12804
rect 26145 12795 26203 12801
rect 26602 12792 26608 12804
rect 26660 12792 26666 12844
rect 22094 12764 22100 12776
rect 21192 12736 22100 12764
rect 22094 12724 22100 12736
rect 22152 12764 22158 12776
rect 22278 12764 22284 12776
rect 22152 12736 22284 12764
rect 22152 12724 22158 12736
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 27801 12767 27859 12773
rect 27801 12764 27813 12767
rect 26712 12736 27813 12764
rect 11330 12696 11336 12708
rect 10336 12668 11336 12696
rect 10229 12659 10287 12665
rect 4356 12628 4384 12656
rect 4798 12628 4804 12640
rect 4172 12600 4384 12628
rect 4759 12600 4804 12628
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 6457 12631 6515 12637
rect 6457 12628 6469 12631
rect 6420 12600 6469 12628
rect 6420 12588 6426 12600
rect 6457 12597 6469 12600
rect 6503 12597 6515 12631
rect 7374 12628 7380 12640
rect 7335 12600 7380 12628
rect 6457 12591 6515 12597
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 8662 12628 8668 12640
rect 8623 12600 8668 12628
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10244 12628 10272 12659
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 20993 12699 21051 12705
rect 20993 12696 21005 12699
rect 20548 12668 21005 12696
rect 9732 12600 10272 12628
rect 9732 12588 9738 12600
rect 10410 12588 10416 12640
rect 10468 12628 10474 12640
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 10468 12600 10609 12628
rect 10468 12588 10474 12600
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 12342 12628 12348 12640
rect 12303 12600 12348 12628
rect 10597 12591 10655 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 13814 12628 13820 12640
rect 13775 12600 13820 12628
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 16942 12628 16948 12640
rect 16903 12600 16948 12628
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 20548 12637 20576 12668
rect 20993 12665 21005 12668
rect 21039 12665 21051 12699
rect 21910 12696 21916 12708
rect 21871 12668 21916 12696
rect 20993 12659 21051 12665
rect 21910 12656 21916 12668
rect 21968 12656 21974 12708
rect 26712 12640 26740 12736
rect 27801 12733 27813 12736
rect 27847 12733 27859 12767
rect 27801 12727 27859 12733
rect 20533 12631 20591 12637
rect 20533 12597 20545 12631
rect 20579 12597 20591 12631
rect 20533 12591 20591 12597
rect 20717 12631 20775 12637
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 20806 12628 20812 12640
rect 20763 12600 20812 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 21818 12588 21824 12640
rect 21876 12628 21882 12640
rect 22097 12631 22155 12637
rect 22097 12628 22109 12631
rect 21876 12600 22109 12628
rect 21876 12588 21882 12600
rect 22097 12597 22109 12600
rect 22143 12597 22155 12631
rect 22097 12591 22155 12597
rect 24397 12631 24455 12637
rect 24397 12597 24409 12631
rect 24443 12628 24455 12631
rect 24854 12628 24860 12640
rect 24443 12600 24860 12628
rect 24443 12597 24455 12600
rect 24397 12591 24455 12597
rect 24854 12588 24860 12600
rect 24912 12588 24918 12640
rect 26694 12628 26700 12640
rect 26655 12600 26700 12628
rect 26694 12588 26700 12600
rect 26752 12588 26758 12640
rect 1104 12538 28888 12560
rect 1104 12486 3350 12538
rect 3402 12486 3414 12538
rect 3466 12486 3478 12538
rect 3530 12486 3542 12538
rect 3594 12486 3606 12538
rect 3658 12486 8150 12538
rect 8202 12486 8214 12538
rect 8266 12486 8278 12538
rect 8330 12486 8342 12538
rect 8394 12486 8406 12538
rect 8458 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 17750 12538
rect 17802 12486 17814 12538
rect 17866 12486 17878 12538
rect 17930 12486 17942 12538
rect 17994 12486 18006 12538
rect 18058 12486 22550 12538
rect 22602 12486 22614 12538
rect 22666 12486 22678 12538
rect 22730 12486 22742 12538
rect 22794 12486 22806 12538
rect 22858 12486 27350 12538
rect 27402 12486 27414 12538
rect 27466 12486 27478 12538
rect 27530 12486 27542 12538
rect 27594 12486 27606 12538
rect 27658 12486 28888 12538
rect 1104 12464 28888 12486
rect 1486 12384 1492 12436
rect 1544 12424 1550 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1544 12396 1593 12424
rect 1544 12384 1550 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2406 12424 2412 12436
rect 2271 12396 2412 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15473 12427 15531 12433
rect 15473 12424 15485 12427
rect 15252 12396 15485 12424
rect 15252 12384 15258 12396
rect 15473 12393 15485 12396
rect 15519 12393 15531 12427
rect 15473 12387 15531 12393
rect 15657 12427 15715 12433
rect 15657 12393 15669 12427
rect 15703 12424 15715 12427
rect 25406 12424 25412 12436
rect 15703 12396 16896 12424
rect 25367 12396 25412 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 6730 12316 6736 12368
rect 6788 12356 6794 12368
rect 12342 12356 12348 12368
rect 6788 12328 9628 12356
rect 12303 12328 12348 12356
rect 6788 12316 6794 12328
rect 9600 12300 9628 12328
rect 12342 12316 12348 12328
rect 12400 12316 12406 12368
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3878 12288 3884 12300
rect 2915 12260 3884 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 7374 12288 7380 12300
rect 7055 12260 7380 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 7374 12248 7380 12260
rect 7432 12288 7438 12300
rect 7653 12291 7711 12297
rect 7653 12288 7665 12291
rect 7432 12260 7665 12288
rect 7432 12248 7438 12260
rect 7653 12257 7665 12260
rect 7699 12257 7711 12291
rect 7653 12251 7711 12257
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 11609 12291 11667 12297
rect 11609 12288 11621 12291
rect 9640 12260 11621 12288
rect 9640 12248 9646 12260
rect 11609 12257 11621 12260
rect 11655 12257 11667 12291
rect 11609 12251 11667 12257
rect 12069 12291 12127 12297
rect 12069 12257 12081 12291
rect 12115 12288 12127 12291
rect 12713 12291 12771 12297
rect 12115 12260 12434 12288
rect 12115 12257 12127 12260
rect 12069 12251 12127 12257
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12220 1823 12223
rect 2685 12223 2743 12229
rect 2685 12220 2697 12223
rect 1811 12192 2697 12220
rect 1811 12189 1823 12192
rect 1765 12183 1823 12189
rect 2685 12189 2697 12192
rect 2731 12220 2743 12223
rect 3234 12220 3240 12232
rect 2731 12192 3240 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12189 6239 12223
rect 6362 12220 6368 12232
rect 6323 12192 6368 12220
rect 6181 12183 6239 12189
rect 2590 12152 2596 12164
rect 2551 12124 2596 12152
rect 2590 12112 2596 12124
rect 2648 12112 2654 12164
rect 3142 12044 3148 12096
rect 3200 12084 3206 12096
rect 3421 12087 3479 12093
rect 3421 12084 3433 12087
rect 3200 12056 3433 12084
rect 3200 12044 3206 12056
rect 3421 12053 3433 12056
rect 3467 12084 3479 12087
rect 3694 12084 3700 12096
rect 3467 12056 3700 12084
rect 3467 12053 3479 12056
rect 3421 12047 3479 12053
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 3878 12084 3884 12096
rect 3839 12056 3884 12084
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 5905 12087 5963 12093
rect 5905 12053 5917 12087
rect 5951 12084 5963 12087
rect 6196 12084 6224 12183
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6687 12192 7297 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12220 11759 12223
rect 12250 12220 12256 12232
rect 11747 12192 12256 12220
rect 11747 12189 11759 12192
rect 11701 12183 11759 12189
rect 6273 12155 6331 12161
rect 6273 12121 6285 12155
rect 6319 12152 6331 12155
rect 6656 12152 6684 12183
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 12406 12220 12434 12260
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 13081 12291 13139 12297
rect 13081 12288 13093 12291
rect 12759 12260 13093 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 13081 12257 13093 12260
rect 13127 12257 13139 12291
rect 16868 12288 16896 12396
rect 25406 12384 25412 12396
rect 25464 12384 25470 12436
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 17092 12328 17724 12356
rect 17092 12316 17098 12328
rect 16942 12288 16948 12300
rect 16868 12260 16948 12288
rect 13081 12251 13139 12257
rect 16942 12248 16948 12260
rect 17000 12288 17006 12300
rect 17696 12297 17724 12328
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 17000 12260 17601 12288
rect 17000 12248 17006 12260
rect 17589 12257 17601 12260
rect 17635 12257 17647 12291
rect 17589 12251 17647 12257
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12257 17739 12291
rect 19978 12288 19984 12300
rect 19939 12260 19984 12288
rect 17681 12251 17739 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 21729 12291 21787 12297
rect 21729 12257 21741 12291
rect 21775 12288 21787 12291
rect 21775 12260 22094 12288
rect 21775 12257 21787 12260
rect 21729 12251 21787 12257
rect 12894 12220 12900 12232
rect 12406 12192 12900 12220
rect 12894 12180 12900 12192
rect 12952 12220 12958 12232
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12952 12192 13001 12220
rect 12952 12180 12958 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12220 13231 12223
rect 16025 12223 16083 12229
rect 13219 12192 13584 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 9858 12152 9864 12164
rect 6319 12124 6684 12152
rect 9771 12124 9864 12152
rect 6319 12121 6331 12124
rect 6273 12115 6331 12121
rect 9858 12112 9864 12124
rect 9916 12152 9922 12164
rect 10962 12152 10968 12164
rect 9916 12124 10968 12152
rect 9916 12112 9922 12124
rect 10962 12112 10968 12124
rect 11020 12152 11026 12164
rect 13188 12152 13216 12183
rect 11020 12124 13216 12152
rect 11020 12112 11026 12124
rect 13556 12096 13584 12192
rect 16025 12189 16037 12223
rect 16071 12220 16083 12223
rect 16758 12220 16764 12232
rect 16071 12192 16764 12220
rect 16071 12189 16083 12192
rect 16025 12183 16083 12189
rect 16758 12180 16764 12192
rect 16816 12220 16822 12232
rect 17034 12220 17040 12232
rect 16816 12192 17040 12220
rect 16816 12180 16822 12192
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 17310 12180 17316 12232
rect 17368 12220 17374 12232
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 17368 12192 17509 12220
rect 17368 12180 17374 12192
rect 17497 12189 17509 12192
rect 17543 12189 17555 12223
rect 22066 12220 22094 12260
rect 24210 12248 24216 12300
rect 24268 12288 24274 12300
rect 24394 12288 24400 12300
rect 24268 12260 24400 12288
rect 24268 12248 24274 12260
rect 24394 12248 24400 12260
rect 24452 12288 24458 12300
rect 24765 12291 24823 12297
rect 24765 12288 24777 12291
rect 24452 12260 24777 12288
rect 24452 12248 24458 12260
rect 24765 12257 24777 12260
rect 24811 12257 24823 12291
rect 24765 12251 24823 12257
rect 24854 12248 24860 12300
rect 24912 12288 24918 12300
rect 24949 12291 25007 12297
rect 24949 12288 24961 12291
rect 24912 12260 24961 12288
rect 24912 12248 24918 12260
rect 24949 12257 24961 12260
rect 24995 12257 25007 12291
rect 24949 12251 25007 12257
rect 22278 12220 22284 12232
rect 22066 12192 22284 12220
rect 17497 12183 17555 12189
rect 22278 12180 22284 12192
rect 22336 12220 22342 12232
rect 25041 12223 25099 12229
rect 25041 12220 25053 12223
rect 22336 12192 25053 12220
rect 22336 12180 22342 12192
rect 25041 12189 25053 12192
rect 25087 12189 25099 12223
rect 25041 12183 25099 12189
rect 15657 12155 15715 12161
rect 15657 12121 15669 12155
rect 15703 12152 15715 12155
rect 17328 12152 17356 12180
rect 15703 12124 17356 12152
rect 20257 12155 20315 12161
rect 15703 12121 15715 12124
rect 15657 12115 15715 12121
rect 20257 12121 20269 12155
rect 20303 12121 20315 12155
rect 23382 12152 23388 12164
rect 21482 12124 23388 12152
rect 20257 12115 20315 12121
rect 6822 12084 6828 12096
rect 5951 12056 6828 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7006 12084 7012 12096
rect 6967 12056 7012 12084
rect 7006 12044 7012 12056
rect 7064 12084 7070 12096
rect 7653 12087 7711 12093
rect 7653 12084 7665 12087
rect 7064 12056 7665 12084
rect 7064 12044 7070 12056
rect 7653 12053 7665 12056
rect 7699 12053 7711 12087
rect 7653 12047 7711 12053
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 12345 12087 12403 12093
rect 12345 12084 12357 12087
rect 10192 12056 12357 12084
rect 10192 12044 10198 12056
rect 12345 12053 12357 12056
rect 12391 12084 12403 12087
rect 12802 12084 12808 12096
rect 12391 12056 12808 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 13538 12084 13544 12096
rect 13499 12056 13544 12084
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 17313 12087 17371 12093
rect 17313 12053 17325 12087
rect 17359 12084 17371 12087
rect 17494 12084 17500 12096
rect 17359 12056 17500 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 17494 12044 17500 12056
rect 17552 12084 17558 12096
rect 17770 12084 17776 12096
rect 17552 12056 17776 12084
rect 17552 12044 17558 12056
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 20272 12084 20300 12115
rect 23382 12112 23388 12124
rect 23440 12112 23446 12164
rect 20622 12084 20628 12096
rect 20272 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 24121 12087 24179 12093
rect 24121 12053 24133 12087
rect 24167 12084 24179 12087
rect 24210 12084 24216 12096
rect 24167 12056 24216 12084
rect 24167 12053 24179 12056
rect 24121 12047 24179 12053
rect 24210 12044 24216 12056
rect 24268 12044 24274 12096
rect 1104 11994 28888 12016
rect 1104 11942 5750 11994
rect 5802 11942 5814 11994
rect 5866 11942 5878 11994
rect 5930 11942 5942 11994
rect 5994 11942 6006 11994
rect 6058 11942 10550 11994
rect 10602 11942 10614 11994
rect 10666 11942 10678 11994
rect 10730 11942 10742 11994
rect 10794 11942 10806 11994
rect 10858 11942 15350 11994
rect 15402 11942 15414 11994
rect 15466 11942 15478 11994
rect 15530 11942 15542 11994
rect 15594 11942 15606 11994
rect 15658 11942 20150 11994
rect 20202 11942 20214 11994
rect 20266 11942 20278 11994
rect 20330 11942 20342 11994
rect 20394 11942 20406 11994
rect 20458 11942 24950 11994
rect 25002 11942 25014 11994
rect 25066 11942 25078 11994
rect 25130 11942 25142 11994
rect 25194 11942 25206 11994
rect 25258 11942 28888 11994
rect 1104 11920 28888 11942
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 3712 11852 4537 11880
rect 3712 11824 3740 11852
rect 4525 11849 4537 11852
rect 4571 11880 4583 11883
rect 4982 11880 4988 11892
rect 4571 11852 4988 11880
rect 4571 11849 4583 11852
rect 4525 11843 4583 11849
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 16666 11840 16672 11892
rect 16724 11880 16730 11892
rect 17126 11880 17132 11892
rect 16724 11852 17132 11880
rect 16724 11840 16730 11852
rect 17126 11840 17132 11852
rect 17184 11880 17190 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 17184 11852 17417 11880
rect 17184 11840 17190 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 20533 11883 20591 11889
rect 20533 11849 20545 11883
rect 20579 11880 20591 11883
rect 20622 11880 20628 11892
rect 20579 11852 20628 11880
rect 20579 11849 20591 11852
rect 20533 11843 20591 11849
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 3694 11812 3700 11824
rect 3542 11784 3700 11812
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 3970 11812 3976 11824
rect 3931 11784 3976 11812
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 13538 11772 13544 11824
rect 13596 11812 13602 11824
rect 18230 11812 18236 11824
rect 13596 11784 18236 11812
rect 13596 11772 13602 11784
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6420 11716 6837 11744
rect 6420 11704 6426 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11744 7067 11747
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 7055 11716 7297 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 12894 11744 12900 11756
rect 12855 11716 12900 11744
rect 7285 11707 7343 11713
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 13127 11716 13369 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13357 11713 13369 11716
rect 13403 11713 13415 11747
rect 17770 11744 17776 11756
rect 17731 11716 17776 11744
rect 13357 11707 13415 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 20806 11744 20812 11756
rect 20763 11716 20812 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 23477 11747 23535 11753
rect 23477 11713 23489 11747
rect 23523 11744 23535 11747
rect 23934 11744 23940 11756
rect 23523 11716 23940 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 23934 11704 23940 11716
rect 23992 11704 23998 11756
rect 27154 11704 27160 11756
rect 27212 11744 27218 11756
rect 27249 11747 27307 11753
rect 27249 11744 27261 11747
rect 27212 11716 27261 11744
rect 27212 11704 27218 11716
rect 27249 11713 27261 11716
rect 27295 11713 27307 11747
rect 28166 11744 28172 11756
rect 28127 11716 28172 11744
rect 27249 11707 27307 11713
rect 28166 11704 28172 11716
rect 28224 11704 28230 11756
rect 1762 11636 1768 11688
rect 1820 11676 1826 11688
rect 4249 11679 4307 11685
rect 4249 11676 4261 11679
rect 1820 11648 4261 11676
rect 1820 11636 1826 11648
rect 4249 11645 4261 11648
rect 4295 11645 4307 11679
rect 4249 11639 4307 11645
rect 4264 11608 4292 11639
rect 4798 11636 4804 11688
rect 4856 11676 4862 11688
rect 6641 11679 6699 11685
rect 6641 11676 6653 11679
rect 4856 11648 6653 11676
rect 4856 11636 4862 11648
rect 6641 11645 6653 11648
rect 6687 11676 6699 11679
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 6687 11648 7849 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 7837 11645 7849 11648
rect 7883 11676 7895 11679
rect 8754 11676 8760 11688
rect 7883 11648 8760 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8754 11636 8760 11648
rect 8812 11676 8818 11688
rect 12713 11679 12771 11685
rect 8812 11648 12434 11676
rect 8812 11636 8818 11648
rect 9030 11608 9036 11620
rect 4264 11580 9036 11608
rect 9030 11568 9036 11580
rect 9088 11568 9094 11620
rect 12406 11608 12434 11648
rect 12713 11645 12725 11679
rect 12759 11676 12771 11679
rect 17865 11679 17923 11685
rect 12759 11648 13952 11676
rect 12759 11645 12771 11648
rect 12713 11639 12771 11645
rect 12728 11608 12756 11639
rect 12406 11580 12756 11608
rect 13924 11552 13952 11648
rect 17865 11645 17877 11679
rect 17911 11645 17923 11679
rect 26694 11676 26700 11688
rect 17865 11639 17923 11645
rect 22066 11648 26700 11676
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2958 11540 2964 11552
rect 2547 11512 2964 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 7469 11543 7527 11549
rect 7469 11509 7481 11543
rect 7515 11540 7527 11543
rect 7558 11540 7564 11552
rect 7515 11512 7564 11540
rect 7515 11509 7527 11512
rect 7469 11503 7527 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 13541 11543 13599 11549
rect 13541 11540 13553 11543
rect 13412 11512 13553 11540
rect 13412 11500 13418 11512
rect 13541 11509 13553 11512
rect 13587 11509 13599 11543
rect 13906 11540 13912 11552
rect 13867 11512 13912 11540
rect 13541 11503 13599 11509
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 17880 11540 17908 11639
rect 18049 11611 18107 11617
rect 18049 11577 18061 11611
rect 18095 11608 18107 11611
rect 19242 11608 19248 11620
rect 18095 11580 19248 11608
rect 18095 11577 18107 11580
rect 18049 11571 18107 11577
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 18138 11540 18144 11552
rect 17880 11512 18144 11540
rect 18138 11500 18144 11512
rect 18196 11540 18202 11552
rect 18414 11540 18420 11552
rect 18196 11512 18420 11540
rect 18196 11500 18202 11512
rect 18414 11500 18420 11512
rect 18472 11540 18478 11552
rect 22066 11540 22094 11648
rect 26694 11636 26700 11648
rect 26752 11636 26758 11688
rect 18472 11512 22094 11540
rect 23661 11543 23719 11549
rect 18472 11500 18478 11512
rect 23661 11509 23673 11543
rect 23707 11540 23719 11543
rect 23842 11540 23848 11552
rect 23707 11512 23848 11540
rect 23707 11509 23719 11512
rect 23661 11503 23719 11509
rect 23842 11500 23848 11512
rect 23900 11500 23906 11552
rect 26786 11500 26792 11552
rect 26844 11540 26850 11552
rect 27065 11543 27123 11549
rect 27065 11540 27077 11543
rect 26844 11512 27077 11540
rect 26844 11500 26850 11512
rect 27065 11509 27077 11512
rect 27111 11509 27123 11543
rect 28350 11540 28356 11552
rect 28311 11512 28356 11540
rect 27065 11503 27123 11509
rect 28350 11500 28356 11512
rect 28408 11500 28414 11552
rect 1104 11450 28888 11472
rect 1104 11398 3350 11450
rect 3402 11398 3414 11450
rect 3466 11398 3478 11450
rect 3530 11398 3542 11450
rect 3594 11398 3606 11450
rect 3658 11398 8150 11450
rect 8202 11398 8214 11450
rect 8266 11398 8278 11450
rect 8330 11398 8342 11450
rect 8394 11398 8406 11450
rect 8458 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 17750 11450
rect 17802 11398 17814 11450
rect 17866 11398 17878 11450
rect 17930 11398 17942 11450
rect 17994 11398 18006 11450
rect 18058 11398 22550 11450
rect 22602 11398 22614 11450
rect 22666 11398 22678 11450
rect 22730 11398 22742 11450
rect 22794 11398 22806 11450
rect 22858 11398 27350 11450
rect 27402 11398 27414 11450
rect 27466 11398 27478 11450
rect 27530 11398 27542 11450
rect 27594 11398 27606 11450
rect 27658 11398 28888 11450
rect 1104 11376 28888 11398
rect 7929 11339 7987 11345
rect 7929 11305 7941 11339
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 7558 11200 7564 11212
rect 7331 11172 7564 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4614 11132 4620 11144
rect 4575 11104 4620 11132
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 7006 11132 7012 11144
rect 6963 11104 7012 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 6549 11067 6607 11073
rect 6549 11064 6561 11067
rect 4632 11036 6561 11064
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 4632 11005 4660 11036
rect 6549 11033 6561 11036
rect 6595 11064 6607 11067
rect 6932 11064 6960 11095
rect 7006 11092 7012 11104
rect 7064 11132 7070 11144
rect 7944 11141 7972 11299
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 11020 11308 11345 11336
rect 11020 11296 11026 11308
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 12989 11339 13047 11345
rect 12989 11336 13001 11339
rect 12860 11308 13001 11336
rect 12860 11296 12866 11308
rect 12989 11305 13001 11308
rect 13035 11336 13047 11339
rect 13725 11339 13783 11345
rect 13725 11336 13737 11339
rect 13035 11308 13737 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13725 11305 13737 11308
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 9582 11200 9588 11212
rect 9543 11172 9588 11200
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 9861 11203 9919 11209
rect 9861 11169 9873 11203
rect 9907 11200 9919 11203
rect 11054 11200 11060 11212
rect 9907 11172 11060 11200
rect 9907 11169 9919 11172
rect 9861 11163 9919 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 13354 11200 13360 11212
rect 13315 11172 13360 11200
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 13740 11209 13768 11299
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11169 13783 11203
rect 16298 11200 16304 11212
rect 13725 11163 13783 11169
rect 16040 11172 16304 11200
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7064 11104 7941 11132
rect 7064 11092 7070 11104
rect 7929 11101 7941 11104
rect 7975 11132 7987 11135
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 7975 11104 8217 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8205 11101 8217 11104
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 16040 11141 16068 11172
rect 16298 11160 16304 11172
rect 16356 11200 16362 11212
rect 22373 11203 22431 11209
rect 16356 11172 17264 11200
rect 16356 11160 16362 11172
rect 9493 11135 9551 11141
rect 9493 11132 9505 11135
rect 8720 11104 9505 11132
rect 8720 11092 8726 11104
rect 9493 11101 9505 11104
rect 9539 11132 9551 11135
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9539 11104 10149 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 16025 11135 16083 11141
rect 16025 11101 16037 11135
rect 16071 11101 16083 11135
rect 16025 11095 16083 11101
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11101 16543 11135
rect 16485 11095 16543 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 16758 11132 16764 11144
rect 16715 11104 16764 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 6595 11036 6960 11064
rect 16500 11064 16528 11095
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 17236 11141 17264 11172
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 23474 11200 23480 11212
rect 22419 11172 23480 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 26786 11200 26792 11212
rect 26747 11172 26792 11200
rect 26786 11160 26792 11172
rect 26844 11160 26850 11212
rect 17221 11135 17279 11141
rect 17221 11101 17233 11135
rect 17267 11132 17279 11135
rect 17310 11132 17316 11144
rect 17267 11104 17316 11132
rect 17267 11101 17279 11104
rect 17221 11095 17279 11101
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17586 11132 17592 11144
rect 17547 11104 17592 11132
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 17773 11135 17831 11141
rect 17773 11101 17785 11135
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 24121 11135 24179 11141
rect 24121 11101 24133 11135
rect 24167 11132 24179 11135
rect 26510 11132 26516 11144
rect 24167 11104 26516 11132
rect 24167 11101 24179 11104
rect 24121 11095 24179 11101
rect 17788 11064 17816 11095
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 18230 11064 18236 11076
rect 16500 11036 17816 11064
rect 17972 11036 18236 11064
rect 6595 11033 6607 11036
rect 6549 11027 6607 11033
rect 6932 11005 6960 11036
rect 16684 11008 16712 11036
rect 4617 10999 4675 11005
rect 4617 10996 4629 10999
rect 4580 10968 4629 10996
rect 4580 10956 4586 10968
rect 4617 10965 4629 10968
rect 4663 10965 4675 10999
rect 4617 10959 4675 10965
rect 6917 10999 6975 11005
rect 6917 10965 6929 10999
rect 6963 10996 6975 10999
rect 10229 10999 10287 11005
rect 6963 10968 6997 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 10229 10965 10241 10999
rect 10275 10996 10287 10999
rect 10410 10996 10416 11008
rect 10275 10968 10416 10996
rect 10275 10965 10287 10968
rect 10229 10959 10287 10965
rect 10410 10956 10416 10968
rect 10468 10956 10474 11008
rect 15381 10999 15439 11005
rect 15381 10965 15393 10999
rect 15427 10996 15439 10999
rect 15746 10996 15752 11008
rect 15427 10968 15752 10996
rect 15427 10965 15439 10968
rect 15381 10959 15439 10965
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 16666 10956 16672 11008
rect 16724 10956 16730 11008
rect 16758 10956 16764 11008
rect 16816 10996 16822 11008
rect 16942 10996 16948 11008
rect 16816 10968 16948 10996
rect 16816 10956 16822 10968
rect 16942 10956 16948 10968
rect 17000 10996 17006 11008
rect 17586 10996 17592 11008
rect 17000 10968 17592 10996
rect 17000 10956 17006 10968
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 17972 11005 18000 11036
rect 18230 11024 18236 11036
rect 18288 11024 18294 11076
rect 23382 11024 23388 11076
rect 23440 11024 23446 11076
rect 23842 11064 23848 11076
rect 23755 11036 23848 11064
rect 23842 11024 23848 11036
rect 23900 11064 23906 11076
rect 23900 11036 27200 11064
rect 23900 11024 23906 11036
rect 17957 10999 18015 11005
rect 17957 10965 17969 10999
rect 18003 10965 18015 10999
rect 27172 10996 27200 11036
rect 27798 11024 27804 11076
rect 27856 11024 27862 11076
rect 27614 10996 27620 11008
rect 27172 10968 27620 10996
rect 17957 10959 18015 10965
rect 27614 10956 27620 10968
rect 27672 10956 27678 11008
rect 27706 10956 27712 11008
rect 27764 10996 27770 11008
rect 28166 10996 28172 11008
rect 27764 10968 28172 10996
rect 27764 10956 27770 10968
rect 28166 10956 28172 10968
rect 28224 10996 28230 11008
rect 28261 10999 28319 11005
rect 28261 10996 28273 10999
rect 28224 10968 28273 10996
rect 28224 10956 28230 10968
rect 28261 10965 28273 10968
rect 28307 10965 28319 10999
rect 28261 10959 28319 10965
rect 1104 10906 28888 10928
rect 1104 10854 5750 10906
rect 5802 10854 5814 10906
rect 5866 10854 5878 10906
rect 5930 10854 5942 10906
rect 5994 10854 6006 10906
rect 6058 10854 10550 10906
rect 10602 10854 10614 10906
rect 10666 10854 10678 10906
rect 10730 10854 10742 10906
rect 10794 10854 10806 10906
rect 10858 10854 15350 10906
rect 15402 10854 15414 10906
rect 15466 10854 15478 10906
rect 15530 10854 15542 10906
rect 15594 10854 15606 10906
rect 15658 10854 20150 10906
rect 20202 10854 20214 10906
rect 20266 10854 20278 10906
rect 20330 10854 20342 10906
rect 20394 10854 20406 10906
rect 20458 10854 24950 10906
rect 25002 10854 25014 10906
rect 25066 10854 25078 10906
rect 25130 10854 25142 10906
rect 25194 10854 25206 10906
rect 25258 10854 28888 10906
rect 1104 10832 28888 10854
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 4580 10764 4629 10792
rect 4580 10752 4586 10764
rect 4617 10761 4629 10764
rect 4663 10792 4675 10795
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 4663 10764 5273 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 5261 10761 5273 10764
rect 5307 10761 5319 10795
rect 5261 10755 5319 10761
rect 9030 10752 9036 10804
rect 9088 10792 9094 10804
rect 9125 10795 9183 10801
rect 9125 10792 9137 10795
rect 9088 10764 9137 10792
rect 9088 10752 9094 10764
rect 9125 10761 9137 10764
rect 9171 10761 9183 10795
rect 9125 10755 9183 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12860 10764 13185 10792
rect 12860 10752 12866 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 10962 10724 10968 10736
rect 9548 10696 10968 10724
rect 9548 10684 9554 10696
rect 10962 10684 10968 10696
rect 11020 10724 11026 10736
rect 11020 10696 11284 10724
rect 11020 10684 11026 10696
rect 4614 10656 4620 10668
rect 4575 10628 4620 10656
rect 4614 10616 4620 10628
rect 4672 10656 4678 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 4672 10628 5273 10656
rect 4672 10616 4678 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 4246 10588 4252 10600
rect 4159 10560 4252 10588
rect 4246 10548 4252 10560
rect 4304 10588 4310 10600
rect 4893 10591 4951 10597
rect 4893 10588 4905 10591
rect 4304 10560 4905 10588
rect 4304 10548 4310 10560
rect 4893 10557 4905 10560
rect 4939 10588 4951 10591
rect 4982 10588 4988 10600
rect 4939 10560 4988 10588
rect 4939 10557 4951 10560
rect 4893 10551 4951 10557
rect 4982 10548 4988 10560
rect 5040 10548 5046 10600
rect 5276 10520 5304 10619
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5592 10628 5641 10656
rect 5592 10616 5598 10628
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 7883 10628 9873 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 9861 10625 9873 10628
rect 9907 10656 9919 10659
rect 10318 10656 10324 10668
rect 9907 10628 10324 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 11054 10656 11060 10668
rect 10468 10628 10513 10656
rect 11015 10628 11060 10656
rect 10468 10616 10474 10628
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11256 10665 11284 10696
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10625 11299 10659
rect 11241 10619 11299 10625
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10656 11943 10659
rect 11974 10656 11980 10668
rect 11931 10628 11980 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 13188 10665 13216 10755
rect 16206 10752 16212 10804
rect 16264 10792 16270 10804
rect 19978 10792 19984 10804
rect 16264 10764 19984 10792
rect 16264 10752 16270 10764
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 23474 10792 23480 10804
rect 23435 10764 23480 10792
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 23934 10792 23940 10804
rect 23895 10764 23940 10792
rect 23934 10752 23940 10764
rect 23992 10752 23998 10804
rect 27154 10752 27160 10804
rect 27212 10792 27218 10804
rect 27249 10795 27307 10801
rect 27249 10792 27261 10795
rect 27212 10764 27261 10792
rect 27212 10752 27218 10764
rect 27249 10761 27261 10764
rect 27295 10761 27307 10795
rect 27614 10792 27620 10804
rect 27575 10764 27620 10792
rect 27249 10755 27307 10761
rect 27614 10752 27620 10764
rect 27672 10752 27678 10804
rect 27706 10752 27712 10804
rect 27764 10792 27770 10804
rect 27764 10764 27809 10792
rect 27764 10752 27770 10764
rect 19242 10724 19248 10736
rect 19203 10696 19248 10724
rect 19242 10684 19248 10696
rect 19300 10684 19306 10736
rect 20717 10727 20775 10733
rect 20717 10693 20729 10727
rect 20763 10724 20775 10727
rect 20993 10727 21051 10733
rect 20993 10724 21005 10727
rect 20763 10696 21005 10724
rect 20763 10693 20775 10696
rect 20717 10687 20775 10693
rect 20993 10693 21005 10696
rect 21039 10693 21051 10727
rect 20993 10687 21051 10693
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12636 10628 12817 10656
rect 9950 10548 9956 10600
rect 10008 10588 10014 10600
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10008 10560 10793 10588
rect 10008 10548 10014 10560
rect 10781 10557 10793 10560
rect 10827 10588 10839 10591
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 10827 10560 11161 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 12636 10532 12664 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 13219 10628 13461 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10656 15715 10659
rect 15746 10656 15752 10668
rect 15703 10628 15752 10656
rect 15703 10625 15715 10628
rect 15657 10619 15715 10625
rect 15488 10588 15516 10619
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 16298 10656 16304 10668
rect 16259 10628 16304 10656
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 18138 10616 18144 10668
rect 18196 10616 18202 10668
rect 20441 10659 20499 10665
rect 20441 10625 20453 10659
rect 20487 10625 20499 10659
rect 20441 10619 20499 10625
rect 20533 10659 20591 10665
rect 20533 10625 20545 10659
rect 20579 10656 20591 10659
rect 21269 10659 21327 10665
rect 21269 10656 21281 10659
rect 20579 10628 21281 10656
rect 20579 10625 20591 10628
rect 20533 10619 20591 10625
rect 21269 10625 21281 10628
rect 21315 10656 21327 10659
rect 21818 10656 21824 10668
rect 21315 10628 21824 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 16209 10591 16267 10597
rect 16209 10588 16221 10591
rect 15488 10560 16221 10588
rect 16209 10557 16221 10560
rect 16255 10588 16267 10591
rect 16666 10588 16672 10600
rect 16255 10560 16672 10588
rect 16255 10557 16267 10560
rect 16209 10551 16267 10557
rect 16666 10548 16672 10560
rect 16724 10588 16730 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 16724 10560 17509 10588
rect 16724 10548 16730 10560
rect 17497 10557 17509 10560
rect 17543 10557 17555 10591
rect 17497 10551 17555 10557
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 20070 10588 20076 10600
rect 19567 10560 20076 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 5629 10523 5687 10529
rect 5629 10520 5641 10523
rect 5276 10492 5641 10520
rect 5629 10489 5641 10492
rect 5675 10489 5687 10523
rect 5629 10483 5687 10489
rect 12069 10523 12127 10529
rect 12069 10489 12081 10523
rect 12115 10520 12127 10523
rect 12618 10520 12624 10532
rect 12115 10492 12624 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 15657 10523 15715 10529
rect 15657 10489 15669 10523
rect 15703 10520 15715 10523
rect 16942 10520 16948 10532
rect 15703 10492 16948 10520
rect 15703 10489 15715 10492
rect 15657 10483 15715 10489
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 20456 10520 20484 10619
rect 21818 10616 21824 10628
rect 21876 10656 21882 10668
rect 23569 10659 23627 10665
rect 23569 10656 23581 10659
rect 21876 10628 23581 10656
rect 21876 10616 21882 10628
rect 23569 10625 23581 10628
rect 23615 10625 23627 10659
rect 23569 10619 23627 10625
rect 20990 10588 20996 10600
rect 20951 10560 20996 10588
rect 20990 10548 20996 10560
rect 21048 10548 21054 10600
rect 21177 10591 21235 10597
rect 21177 10557 21189 10591
rect 21223 10588 21235 10591
rect 21450 10588 21456 10600
rect 21223 10560 21456 10588
rect 21223 10557 21235 10560
rect 21177 10551 21235 10557
rect 20898 10520 20904 10532
rect 20456 10492 20904 10520
rect 20898 10480 20904 10492
rect 20956 10520 20962 10532
rect 21192 10520 21220 10551
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 22925 10591 22983 10597
rect 22925 10557 22937 10591
rect 22971 10588 22983 10591
rect 23385 10591 23443 10597
rect 23385 10588 23397 10591
rect 22971 10560 23397 10588
rect 22971 10557 22983 10560
rect 22925 10551 22983 10557
rect 23385 10557 23397 10560
rect 23431 10588 23443 10591
rect 24210 10588 24216 10600
rect 23431 10560 24216 10588
rect 23431 10557 23443 10560
rect 23385 10551 23443 10557
rect 24210 10548 24216 10560
rect 24268 10548 24274 10600
rect 27801 10591 27859 10597
rect 27801 10588 27813 10591
rect 26712 10560 27813 10588
rect 20956 10492 21220 10520
rect 20956 10480 20962 10492
rect 26712 10464 26740 10560
rect 27801 10557 27813 10560
rect 27847 10557 27859 10591
rect 27801 10551 27859 10557
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10413 10455 10471 10461
rect 10413 10452 10425 10455
rect 10192 10424 10425 10452
rect 10192 10412 10198 10424
rect 10413 10421 10425 10424
rect 10459 10421 10471 10455
rect 15930 10452 15936 10464
rect 15891 10424 15936 10452
rect 10413 10415 10471 10421
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 16301 10455 16359 10461
rect 16301 10421 16313 10455
rect 16347 10452 16359 10455
rect 16758 10452 16764 10464
rect 16347 10424 16764 10452
rect 16347 10421 16359 10424
rect 16301 10415 16359 10421
rect 16758 10412 16764 10424
rect 16816 10412 16822 10464
rect 20346 10412 20352 10464
rect 20404 10452 20410 10464
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 20404 10424 20729 10452
rect 20404 10412 20410 10424
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 26694 10452 26700 10464
rect 26655 10424 26700 10452
rect 20717 10415 20775 10421
rect 26694 10412 26700 10424
rect 26752 10412 26758 10464
rect 1104 10362 28888 10384
rect 1104 10310 3350 10362
rect 3402 10310 3414 10362
rect 3466 10310 3478 10362
rect 3530 10310 3542 10362
rect 3594 10310 3606 10362
rect 3658 10310 8150 10362
rect 8202 10310 8214 10362
rect 8266 10310 8278 10362
rect 8330 10310 8342 10362
rect 8394 10310 8406 10362
rect 8458 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 17750 10362
rect 17802 10310 17814 10362
rect 17866 10310 17878 10362
rect 17930 10310 17942 10362
rect 17994 10310 18006 10362
rect 18058 10310 22550 10362
rect 22602 10310 22614 10362
rect 22666 10310 22678 10362
rect 22730 10310 22742 10362
rect 22794 10310 22806 10362
rect 22858 10310 27350 10362
rect 27402 10310 27414 10362
rect 27466 10310 27478 10362
rect 27530 10310 27542 10362
rect 27594 10310 27606 10362
rect 27658 10310 28888 10362
rect 1104 10288 28888 10310
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12710 10248 12716 10260
rect 12575 10220 12716 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12710 10208 12716 10220
rect 12768 10248 12774 10260
rect 13170 10248 13176 10260
rect 12768 10220 13176 10248
rect 12768 10208 12774 10220
rect 13170 10208 13176 10220
rect 13228 10248 13234 10260
rect 13722 10248 13728 10260
rect 13228 10220 13728 10248
rect 13228 10208 13234 10220
rect 13722 10208 13728 10220
rect 13780 10248 13786 10260
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 13780 10220 13829 10248
rect 13780 10208 13786 10220
rect 13817 10217 13829 10220
rect 13863 10217 13875 10251
rect 13817 10211 13875 10217
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 13964 10220 14933 10248
rect 13964 10208 13970 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 21818 10248 21824 10260
rect 21779 10220 21824 10248
rect 14921 10211 14979 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 4614 10180 4620 10192
rect 4575 10152 4620 10180
rect 4614 10140 4620 10152
rect 4672 10180 4678 10192
rect 5261 10183 5319 10189
rect 5261 10180 5273 10183
rect 4672 10152 5273 10180
rect 4672 10140 4678 10152
rect 5261 10149 5273 10152
rect 5307 10149 5319 10183
rect 6730 10180 6736 10192
rect 5261 10143 5319 10149
rect 5920 10152 6736 10180
rect 4893 10115 4951 10121
rect 4893 10081 4905 10115
rect 4939 10112 4951 10115
rect 4982 10112 4988 10124
rect 4939 10084 4988 10112
rect 4939 10081 4951 10084
rect 4893 10075 4951 10081
rect 4982 10072 4988 10084
rect 5040 10072 5046 10124
rect 5920 10121 5948 10152
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 9493 10183 9551 10189
rect 9493 10149 9505 10183
rect 9539 10180 9551 10183
rect 9766 10180 9772 10192
rect 9539 10152 9772 10180
rect 9539 10149 9551 10152
rect 9493 10143 9551 10149
rect 9766 10140 9772 10152
rect 9824 10180 9830 10192
rect 10137 10183 10195 10189
rect 10137 10180 10149 10183
rect 9824 10152 10149 10180
rect 9824 10140 9830 10152
rect 10137 10149 10149 10152
rect 10183 10180 10195 10183
rect 10410 10180 10416 10192
rect 10183 10152 10416 10180
rect 10183 10149 10195 10152
rect 10137 10143 10195 10149
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 12161 10115 12219 10121
rect 12161 10081 12173 10115
rect 12207 10112 12219 10115
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 12207 10084 15761 10112
rect 12207 10081 12219 10084
rect 12161 10075 12219 10081
rect 15749 10081 15761 10084
rect 15795 10112 15807 10115
rect 16114 10112 16120 10124
rect 15795 10084 16120 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 4246 10044 4252 10056
rect 4207 10016 4252 10044
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5592 10016 5825 10044
rect 5592 10004 5598 10016
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 6196 10044 6224 10075
rect 16114 10072 16120 10084
rect 16172 10072 16178 10124
rect 17586 10072 17592 10124
rect 17644 10112 17650 10124
rect 17773 10115 17831 10121
rect 17773 10112 17785 10115
rect 17644 10084 17785 10112
rect 17644 10072 17650 10084
rect 17773 10081 17785 10084
rect 17819 10081 17831 10115
rect 20346 10112 20352 10124
rect 20307 10084 20352 10112
rect 17773 10075 17831 10081
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 6641 10047 6699 10053
rect 6641 10044 6653 10047
rect 6196 10016 6653 10044
rect 5813 10007 5871 10013
rect 6641 10013 6653 10016
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 4982 9936 4988 9988
rect 5040 9976 5046 9988
rect 6457 9979 6515 9985
rect 6457 9976 6469 9979
rect 5040 9948 6469 9976
rect 5040 9936 5046 9948
rect 6457 9945 6469 9948
rect 6503 9945 6515 9979
rect 6656 9976 6684 10007
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 9125 10047 9183 10053
rect 6880 10016 7236 10044
rect 6880 10004 6886 10016
rect 6914 9976 6920 9988
rect 6656 9948 6920 9976
rect 6457 9939 6515 9945
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 7208 9917 7236 10016
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 9171 10016 9781 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9769 10013 9781 10016
rect 9815 10044 9827 10047
rect 9950 10044 9956 10056
rect 9815 10016 9956 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 9950 10004 9956 10016
rect 10008 10004 10014 10056
rect 10318 10004 10324 10056
rect 10376 10044 10382 10056
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 10376 10016 10425 10044
rect 10376 10004 10382 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12676 10016 12817 10044
rect 12676 10004 12682 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 13170 10044 13176 10056
rect 13131 10016 13176 10044
rect 12805 10007 12863 10013
rect 12820 9976 12848 10007
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13078 9976 13084 9988
rect 12820 9948 13084 9976
rect 13078 9936 13084 9948
rect 13136 9976 13142 9988
rect 13464 9976 13492 10007
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 13780 10016 13829 10044
rect 13780 10004 13786 10016
rect 13817 10013 13829 10016
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 15105 10047 15163 10053
rect 15105 10013 15117 10047
rect 15151 10013 15163 10047
rect 18138 10044 18144 10056
rect 17158 10016 18144 10044
rect 15105 10007 15163 10013
rect 13136 9948 13492 9976
rect 15120 9976 15148 10007
rect 18138 10004 18144 10016
rect 18196 10044 18202 10056
rect 19426 10044 19432 10056
rect 18196 10016 19432 10044
rect 18196 10004 18202 10016
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 20070 10044 20076 10056
rect 20031 10016 20076 10044
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 15930 9976 15936 9988
rect 15120 9948 15936 9976
rect 13136 9936 13142 9948
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 16025 9979 16083 9985
rect 16025 9945 16037 9979
rect 16071 9945 16083 9979
rect 19444 9976 19472 10004
rect 23382 9976 23388 9988
rect 19444 9948 20838 9976
rect 22066 9948 23388 9976
rect 16025 9939 16083 9945
rect 4617 9911 4675 9917
rect 4617 9908 4629 9911
rect 4580 9880 4629 9908
rect 4580 9868 4586 9880
rect 4617 9877 4629 9880
rect 4663 9908 4675 9911
rect 5261 9911 5319 9917
rect 5261 9908 5273 9911
rect 4663 9880 5273 9908
rect 4663 9877 4675 9880
rect 4617 9871 4675 9877
rect 5261 9877 5273 9880
rect 5307 9877 5319 9911
rect 5261 9871 5319 9877
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9908 7251 9911
rect 8294 9908 8300 9920
rect 7239 9880 8300 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9908 9551 9911
rect 9674 9908 9680 9920
rect 9539 9880 9680 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 9674 9868 9680 9880
rect 9732 9908 9738 9920
rect 10134 9908 10140 9920
rect 9732 9880 10140 9908
rect 9732 9868 9738 9880
rect 10134 9868 10140 9880
rect 10192 9868 10198 9920
rect 16040 9908 16068 9939
rect 16758 9908 16764 9920
rect 16040 9880 16764 9908
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 20732 9908 20760 9948
rect 22066 9908 22094 9948
rect 23382 9936 23388 9948
rect 23440 9936 23446 9988
rect 20732 9880 22094 9908
rect 1104 9818 28888 9840
rect 1104 9766 5750 9818
rect 5802 9766 5814 9818
rect 5866 9766 5878 9818
rect 5930 9766 5942 9818
rect 5994 9766 6006 9818
rect 6058 9766 10550 9818
rect 10602 9766 10614 9818
rect 10666 9766 10678 9818
rect 10730 9766 10742 9818
rect 10794 9766 10806 9818
rect 10858 9766 15350 9818
rect 15402 9766 15414 9818
rect 15466 9766 15478 9818
rect 15530 9766 15542 9818
rect 15594 9766 15606 9818
rect 15658 9766 20150 9818
rect 20202 9766 20214 9818
rect 20266 9766 20278 9818
rect 20330 9766 20342 9818
rect 20394 9766 20406 9818
rect 20458 9766 24950 9818
rect 25002 9766 25014 9818
rect 25066 9766 25078 9818
rect 25130 9766 25142 9818
rect 25194 9766 25206 9818
rect 25258 9766 28888 9818
rect 1104 9744 28888 9766
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 4580 9676 4629 9704
rect 4580 9664 4586 9676
rect 4617 9673 4629 9676
rect 4663 9704 4675 9707
rect 5261 9707 5319 9713
rect 5261 9704 5273 9707
rect 4663 9676 5273 9704
rect 4663 9673 4675 9676
rect 4617 9667 4675 9673
rect 5261 9673 5273 9676
rect 5307 9673 5319 9707
rect 5261 9667 5319 9673
rect 9125 9707 9183 9713
rect 9125 9673 9137 9707
rect 9171 9704 9183 9707
rect 9674 9704 9680 9716
rect 9171 9676 9680 9704
rect 9171 9673 9183 9676
rect 9125 9667 9183 9673
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 10318 9664 10324 9716
rect 10376 9704 10382 9716
rect 10376 9676 12296 9704
rect 10376 9664 10382 9676
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 11974 9636 11980 9648
rect 6972 9608 10732 9636
rect 11935 9608 11980 9636
rect 6972 9596 6978 9608
rect 4614 9568 4620 9580
rect 4575 9540 4620 9568
rect 4614 9528 4620 9540
rect 4672 9568 4678 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 4672 9540 5273 9568
rect 4672 9528 4678 9540
rect 5261 9537 5273 9540
rect 5307 9537 5319 9571
rect 8294 9568 8300 9580
rect 8207 9540 8300 9568
rect 5261 9531 5319 9537
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 9582 9568 9588 9580
rect 8536 9540 9588 9568
rect 8536 9528 8542 9540
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9766 9568 9772 9580
rect 9727 9540 9772 9568
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10704 9577 10732 9608
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 12268 9645 12296 9676
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 12805 9707 12863 9713
rect 12805 9704 12817 9707
rect 12768 9676 12817 9704
rect 12768 9664 12774 9676
rect 12805 9673 12817 9676
rect 12851 9704 12863 9707
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 12851 9676 13461 9704
rect 12851 9673 12863 9676
rect 12805 9667 12863 9673
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13449 9667 13507 9673
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12299 9608 12434 9636
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 10008 9540 10149 9568
rect 10008 9528 10014 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11112 9540 11805 9568
rect 11112 9528 11118 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 12406 9568 12434 9608
rect 15930 9596 15936 9648
rect 15988 9636 15994 9648
rect 17589 9639 17647 9645
rect 17589 9636 17601 9639
rect 15988 9608 17601 9636
rect 15988 9596 15994 9608
rect 17589 9605 17601 9608
rect 17635 9605 17647 9639
rect 17589 9599 17647 9605
rect 16574 9568 16580 9580
rect 12406 9540 16580 9568
rect 11793 9531 11851 9537
rect 16574 9528 16580 9540
rect 16632 9528 16638 9580
rect 16942 9568 16948 9580
rect 16903 9540 16948 9568
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 17218 9568 17224 9580
rect 17179 9540 17224 9568
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 17773 9571 17831 9577
rect 17773 9537 17785 9571
rect 17819 9568 17831 9571
rect 18506 9568 18512 9580
rect 17819 9540 18512 9568
rect 17819 9537 17831 9540
rect 17773 9531 17831 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 24673 9571 24731 9577
rect 24673 9537 24685 9571
rect 24719 9568 24731 9571
rect 24854 9568 24860 9580
rect 24719 9540 24860 9568
rect 24719 9537 24731 9540
rect 24673 9531 24731 9537
rect 24854 9528 24860 9540
rect 24912 9528 24918 9580
rect 27154 9528 27160 9580
rect 27212 9568 27218 9580
rect 27249 9571 27307 9577
rect 27249 9568 27261 9571
rect 27212 9540 27261 9568
rect 27212 9528 27218 9540
rect 27249 9537 27261 9540
rect 27295 9537 27307 9571
rect 27249 9531 27307 9537
rect 28169 9571 28227 9577
rect 28169 9537 28181 9571
rect 28215 9568 28227 9571
rect 28258 9568 28264 9580
rect 28215 9540 28264 9568
rect 28215 9537 28227 9540
rect 28169 9531 28227 9537
rect 28258 9528 28264 9540
rect 28316 9528 28322 9580
rect 4246 9500 4252 9512
rect 4159 9472 4252 9500
rect 4246 9460 4252 9472
rect 4304 9500 4310 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4304 9472 4905 9500
rect 4304 9460 4310 9472
rect 4893 9469 4905 9472
rect 4939 9500 4951 9503
rect 4982 9500 4988 9512
rect 4939 9472 4988 9500
rect 4939 9469 4951 9472
rect 4893 9463 4951 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 8312 9432 8340 9528
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 8435 9472 8769 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 9490 9500 9496 9512
rect 8757 9463 8815 9469
rect 8864 9472 9496 9500
rect 8570 9432 8576 9444
rect 8312 9404 8576 9432
rect 8570 9392 8576 9404
rect 8628 9432 8634 9444
rect 8864 9432 8892 9472
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 9600 9472 10517 9500
rect 9122 9432 9128 9444
rect 8628 9404 8892 9432
rect 9083 9404 9128 9432
rect 8628 9392 8634 9404
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 9600 9364 9628 9472
rect 10505 9469 10517 9472
rect 10551 9500 10563 9503
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10551 9472 11161 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 11149 9469 11161 9472
rect 11195 9500 11207 9503
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 11195 9472 11621 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11609 9469 11621 9472
rect 11655 9500 11667 9503
rect 12250 9500 12256 9512
rect 11655 9472 12256 9500
rect 11655 9469 11667 9472
rect 11609 9463 11667 9469
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12768 9472 12817 9500
rect 12768 9460 12774 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 13078 9460 13084 9512
rect 13136 9500 13142 9512
rect 13173 9503 13231 9509
rect 13173 9500 13185 9503
rect 13136 9472 13185 9500
rect 13136 9460 13142 9472
rect 13173 9469 13185 9472
rect 13219 9469 13231 9503
rect 16758 9500 16764 9512
rect 16719 9472 16764 9500
rect 13173 9463 13231 9469
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 17037 9503 17095 9509
rect 17037 9469 17049 9503
rect 17083 9469 17095 9503
rect 17037 9463 17095 9469
rect 17052 9432 17080 9463
rect 17126 9460 17132 9512
rect 17184 9500 17190 9512
rect 17184 9472 17229 9500
rect 17184 9460 17190 9472
rect 17957 9435 18015 9441
rect 17957 9432 17969 9435
rect 17052 9404 17969 9432
rect 17957 9401 17969 9404
rect 18003 9401 18015 9435
rect 17957 9395 18015 9401
rect 8812 9336 9628 9364
rect 8812 9324 8818 9336
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9769 9367 9827 9373
rect 9769 9364 9781 9367
rect 9732 9336 9781 9364
rect 9732 9324 9738 9336
rect 9769 9333 9781 9336
rect 9815 9333 9827 9367
rect 10870 9364 10876 9376
rect 10831 9336 10876 9364
rect 9769 9327 9827 9333
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 24857 9367 24915 9373
rect 24857 9333 24869 9367
rect 24903 9364 24915 9367
rect 25958 9364 25964 9376
rect 24903 9336 25964 9364
rect 24903 9333 24915 9336
rect 24857 9327 24915 9333
rect 25958 9324 25964 9336
rect 26016 9324 26022 9376
rect 26786 9324 26792 9376
rect 26844 9364 26850 9376
rect 27065 9367 27123 9373
rect 27065 9364 27077 9367
rect 26844 9336 27077 9364
rect 26844 9324 26850 9336
rect 27065 9333 27077 9336
rect 27111 9333 27123 9367
rect 28350 9364 28356 9376
rect 28311 9336 28356 9364
rect 27065 9327 27123 9333
rect 28350 9324 28356 9336
rect 28408 9324 28414 9376
rect 1104 9274 28888 9296
rect 1104 9222 3350 9274
rect 3402 9222 3414 9274
rect 3466 9222 3478 9274
rect 3530 9222 3542 9274
rect 3594 9222 3606 9274
rect 3658 9222 8150 9274
rect 8202 9222 8214 9274
rect 8266 9222 8278 9274
rect 8330 9222 8342 9274
rect 8394 9222 8406 9274
rect 8458 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 17750 9274
rect 17802 9222 17814 9274
rect 17866 9222 17878 9274
rect 17930 9222 17942 9274
rect 17994 9222 18006 9274
rect 18058 9222 22550 9274
rect 22602 9222 22614 9274
rect 22666 9222 22678 9274
rect 22730 9222 22742 9274
rect 22794 9222 22806 9274
rect 22858 9222 27350 9274
rect 27402 9222 27414 9274
rect 27466 9222 27478 9274
rect 27530 9222 27542 9274
rect 27594 9222 27606 9274
rect 27658 9222 28888 9274
rect 1104 9200 28888 9222
rect 12250 9160 12256 9172
rect 12211 9132 12256 9160
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12710 9160 12716 9172
rect 12671 9132 12716 9160
rect 12710 9120 12716 9132
rect 12768 9160 12774 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12768 9132 13001 9160
rect 12768 9120 12774 9132
rect 12989 9129 13001 9132
rect 13035 9160 13047 9163
rect 13078 9160 13084 9172
rect 13035 9132 13084 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 13078 9120 13084 9132
rect 13136 9160 13142 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 13136 9132 13369 9160
rect 13136 9120 13142 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9129 14243 9163
rect 14185 9123 14243 9129
rect 4614 9092 4620 9104
rect 4575 9064 4620 9092
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 4246 9024 4252 9036
rect 4207 8996 4252 9024
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 13372 9033 13400 9123
rect 14200 9033 14228 9123
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 9180 8996 9413 9024
rect 9180 8984 9186 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 13357 9027 13415 9033
rect 13357 8993 13369 9027
rect 13403 9024 13415 9027
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13403 8996 14197 9024
rect 13403 8993 13415 8996
rect 13357 8987 13415 8993
rect 14185 8993 14197 8996
rect 14231 9024 14243 9027
rect 14829 9027 14887 9033
rect 14829 9024 14841 9027
rect 14231 8996 14841 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 14829 8993 14841 8996
rect 14875 8993 14887 9027
rect 25958 9024 25964 9036
rect 25919 8996 25964 9024
rect 14829 8987 14887 8993
rect 25958 8984 25964 8996
rect 26016 8984 26022 9036
rect 26786 9024 26792 9036
rect 26747 8996 26792 9024
rect 26786 8984 26792 8996
rect 26844 8984 26850 9036
rect 7098 8956 7104 8968
rect 7059 8928 7104 8956
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 8478 8956 8484 8968
rect 7774 8928 8484 8956
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 10928 8928 11805 8956
rect 10928 8916 10934 8928
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 8110 8888 8116 8900
rect 8071 8860 8116 8888
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 11977 8891 12035 8897
rect 11977 8857 11989 8891
rect 12023 8888 12035 8891
rect 12710 8888 12716 8900
rect 12023 8860 12716 8888
rect 12023 8857 12035 8860
rect 11977 8851 12035 8857
rect 12710 8848 12716 8860
rect 12768 8888 12774 8900
rect 13740 8888 13768 8919
rect 14568 8888 14596 8919
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 20070 8956 20076 8968
rect 19392 8928 20076 8956
rect 19392 8916 19398 8928
rect 20070 8916 20076 8928
rect 20128 8956 20134 8968
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 20128 8928 21557 8956
rect 20128 8916 20134 8928
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 21545 8919 21603 8925
rect 23382 8916 23388 8968
rect 23440 8956 23446 8968
rect 26237 8959 26295 8965
rect 23440 8928 24886 8956
rect 23440 8916 23446 8928
rect 26237 8925 26249 8959
rect 26283 8956 26295 8959
rect 26510 8956 26516 8968
rect 26283 8928 26516 8956
rect 26283 8925 26295 8928
rect 26237 8919 26295 8925
rect 26510 8916 26516 8928
rect 26568 8916 26574 8968
rect 21818 8888 21824 8900
rect 12768 8860 14596 8888
rect 21779 8860 21824 8888
rect 12768 8848 12774 8860
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 23934 8888 23940 8900
rect 23046 8860 23940 8888
rect 23934 8848 23940 8860
rect 23992 8848 23998 8900
rect 27798 8848 27804 8900
rect 27856 8848 27862 8900
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4617 8823 4675 8829
rect 4617 8820 4629 8823
rect 4580 8792 4629 8820
rect 4580 8780 4586 8792
rect 4617 8789 4629 8792
rect 4663 8820 4675 8823
rect 5442 8820 5448 8832
rect 4663 8792 5448 8820
rect 4663 8789 4675 8792
rect 4617 8783 4675 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 23290 8820 23296 8832
rect 23251 8792 23296 8820
rect 23290 8780 23296 8792
rect 23348 8780 23354 8832
rect 24486 8820 24492 8832
rect 24447 8792 24492 8820
rect 24486 8780 24492 8792
rect 24544 8780 24550 8832
rect 25958 8780 25964 8832
rect 26016 8820 26022 8832
rect 27614 8820 27620 8832
rect 26016 8792 27620 8820
rect 26016 8780 26022 8792
rect 27614 8780 27620 8792
rect 27672 8780 27678 8832
rect 28258 8820 28264 8832
rect 28219 8792 28264 8820
rect 28258 8780 28264 8792
rect 28316 8780 28322 8832
rect 1104 8730 28888 8752
rect 1104 8678 5750 8730
rect 5802 8678 5814 8730
rect 5866 8678 5878 8730
rect 5930 8678 5942 8730
rect 5994 8678 6006 8730
rect 6058 8678 10550 8730
rect 10602 8678 10614 8730
rect 10666 8678 10678 8730
rect 10730 8678 10742 8730
rect 10794 8678 10806 8730
rect 10858 8678 15350 8730
rect 15402 8678 15414 8730
rect 15466 8678 15478 8730
rect 15530 8678 15542 8730
rect 15594 8678 15606 8730
rect 15658 8678 20150 8730
rect 20202 8678 20214 8730
rect 20266 8678 20278 8730
rect 20330 8678 20342 8730
rect 20394 8678 20406 8730
rect 20458 8678 24950 8730
rect 25002 8678 25014 8730
rect 25066 8678 25078 8730
rect 25130 8678 25142 8730
rect 25194 8678 25206 8730
rect 25258 8678 28888 8730
rect 1104 8656 28888 8678
rect 2958 8616 2964 8628
rect 2919 8588 2964 8616
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 8110 8576 8116 8628
rect 8168 8576 8174 8628
rect 13078 8616 13084 8628
rect 13039 8588 13084 8616
rect 13078 8576 13084 8588
rect 13136 8616 13142 8628
rect 13725 8619 13783 8625
rect 13725 8616 13737 8619
rect 13136 8588 13737 8616
rect 13136 8576 13142 8588
rect 13725 8585 13737 8588
rect 13771 8616 13783 8619
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 13771 8588 14381 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 14369 8585 14381 8588
rect 14415 8616 14427 8619
rect 15013 8619 15071 8625
rect 15013 8616 15025 8619
rect 14415 8588 15025 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 15013 8585 15025 8588
rect 15059 8585 15071 8619
rect 15013 8579 15071 8585
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 17957 8619 18015 8625
rect 17957 8616 17969 8619
rect 16632 8588 17969 8616
rect 16632 8576 16638 8588
rect 17957 8585 17969 8588
rect 18003 8585 18015 8619
rect 17957 8579 18015 8585
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 8128 8548 8156 8576
rect 17972 8548 18000 8579
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 7944 8520 8892 8548
rect 17972 8520 18245 8548
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 3053 8483 3111 8489
rect 2363 8452 2636 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 2608 8353 2636 8452
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3234 8480 3240 8492
rect 3099 8452 3240 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7944 8489 7972 8520
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 7156 8452 7205 8480
rect 7156 8440 7162 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8480 8447 8483
rect 8570 8480 8576 8492
rect 8435 8452 8576 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 8754 8480 8760 8492
rect 8715 8452 8760 8480
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 8864 8489 8892 8520
rect 18233 8517 18245 8520
rect 18279 8548 18291 8551
rect 20438 8548 20444 8560
rect 18279 8520 20444 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 20438 8508 20444 8520
rect 20496 8508 20502 8560
rect 21174 8548 21180 8560
rect 21135 8520 21180 8548
rect 21174 8508 21180 8520
rect 21232 8508 21238 8560
rect 21376 8548 21404 8579
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 21876 8588 22477 8616
rect 21876 8576 21882 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 22465 8579 22523 8585
rect 24486 8576 24492 8628
rect 24544 8616 24550 8628
rect 24765 8619 24823 8625
rect 24765 8616 24777 8619
rect 24544 8588 24777 8616
rect 24544 8576 24550 8588
rect 24765 8585 24777 8588
rect 24811 8585 24823 8619
rect 24765 8579 24823 8585
rect 24854 8576 24860 8628
rect 24912 8616 24918 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 24912 8588 25237 8616
rect 24912 8576 24918 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 25225 8579 25283 8585
rect 27154 8576 27160 8628
rect 27212 8616 27218 8628
rect 27249 8619 27307 8625
rect 27249 8616 27261 8619
rect 27212 8588 27261 8616
rect 27212 8576 27218 8588
rect 27249 8585 27261 8588
rect 27295 8585 27307 8619
rect 27614 8616 27620 8628
rect 27575 8588 27620 8616
rect 27249 8579 27307 8585
rect 27614 8576 27620 8588
rect 27672 8576 27678 8628
rect 27709 8619 27767 8625
rect 27709 8585 27721 8619
rect 27755 8616 27767 8619
rect 28258 8616 28264 8628
rect 27755 8588 28264 8616
rect 27755 8585 27767 8588
rect 27709 8579 27767 8585
rect 28258 8576 28264 8588
rect 28316 8576 28322 8628
rect 21376 8520 22692 8548
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8449 8907 8483
rect 12710 8480 12716 8492
rect 12671 8452 12716 8480
rect 8849 8443 8907 8449
rect 12710 8440 12716 8452
rect 12768 8480 12774 8492
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 12768 8452 13369 8480
rect 12768 8440 12774 8452
rect 13357 8449 13369 8452
rect 13403 8480 13415 8483
rect 13722 8480 13728 8492
rect 13403 8452 13728 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 13722 8440 13728 8452
rect 13780 8480 13786 8492
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 13780 8452 14013 8480
rect 13780 8440 13786 8452
rect 14001 8449 14013 8452
rect 14047 8480 14059 8483
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 14047 8452 14657 8480
rect 14047 8449 14059 8452
rect 14001 8443 14059 8449
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8480 20867 8483
rect 20898 8480 20904 8492
rect 20855 8452 20904 8480
rect 20855 8449 20867 8452
rect 20809 8443 20867 8449
rect 20898 8440 20904 8452
rect 20956 8480 20962 8492
rect 21913 8483 21971 8489
rect 21913 8480 21925 8483
rect 20956 8452 21925 8480
rect 20956 8440 20962 8452
rect 21913 8449 21925 8452
rect 21959 8449 21971 8483
rect 22094 8480 22100 8492
rect 22055 8452 22100 8480
rect 21913 8443 21971 8449
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 22664 8489 22692 8520
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 23290 8440 23296 8492
rect 23348 8480 23354 8492
rect 24857 8483 24915 8489
rect 24857 8480 24869 8483
rect 23348 8452 24869 8480
rect 23348 8440 23354 8452
rect 24857 8449 24869 8452
rect 24903 8449 24915 8483
rect 24857 8443 24915 8449
rect 3142 8412 3148 8424
rect 3103 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8412 3206 8424
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3200 8384 3617 8412
rect 3200 8372 3206 8384
rect 3605 8381 3617 8384
rect 3651 8412 3663 8415
rect 3878 8412 3884 8424
rect 3651 8384 3884 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 7282 8372 7288 8424
rect 7340 8412 7346 8424
rect 7653 8415 7711 8421
rect 7653 8412 7665 8415
rect 7340 8384 7665 8412
rect 7340 8372 7346 8384
rect 7653 8381 7665 8384
rect 7699 8381 7711 8415
rect 8772 8412 8800 8440
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8772 8384 9321 8412
rect 7653 8375 7711 8381
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12618 8412 12624 8424
rect 12483 8384 12624 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12618 8372 12624 8384
rect 12676 8412 12682 8424
rect 13078 8412 13084 8424
rect 12676 8384 13084 8412
rect 12676 8372 12682 8384
rect 13078 8372 13084 8384
rect 13136 8412 13142 8424
rect 24210 8412 24216 8424
rect 13136 8384 13768 8412
rect 24123 8384 24216 8412
rect 13136 8372 13142 8384
rect 13740 8353 13768 8384
rect 24210 8372 24216 8384
rect 24268 8412 24274 8424
rect 24670 8412 24676 8424
rect 24268 8384 24676 8412
rect 24268 8372 24274 8384
rect 24670 8372 24676 8384
rect 24728 8372 24734 8424
rect 26694 8412 26700 8424
rect 26607 8384 26700 8412
rect 26694 8372 26700 8384
rect 26752 8412 26758 8424
rect 27706 8412 27712 8424
rect 26752 8384 27712 8412
rect 26752 8372 26758 8384
rect 27706 8372 27712 8384
rect 27764 8412 27770 8424
rect 27801 8415 27859 8421
rect 27801 8412 27813 8415
rect 27764 8384 27813 8412
rect 27764 8372 27770 8384
rect 27801 8381 27813 8384
rect 27847 8381 27859 8415
rect 27801 8375 27859 8381
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8313 2651 8347
rect 2593 8307 2651 8313
rect 13725 8347 13783 8353
rect 13725 8313 13737 8347
rect 13771 8344 13783 8347
rect 14369 8347 14427 8353
rect 14369 8344 14381 8347
rect 13771 8316 14381 8344
rect 13771 8313 13783 8316
rect 13725 8307 13783 8313
rect 14369 8313 14381 8316
rect 14415 8344 14427 8347
rect 15013 8347 15071 8353
rect 15013 8344 15025 8347
rect 14415 8316 15025 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 15013 8313 15025 8316
rect 15059 8344 15071 8347
rect 15289 8347 15347 8353
rect 15289 8344 15301 8347
rect 15059 8316 15301 8344
rect 15059 8313 15071 8316
rect 15013 8307 15071 8313
rect 15289 8313 15301 8316
rect 15335 8313 15347 8347
rect 15289 8307 15347 8313
rect 1946 8236 1952 8288
rect 2004 8276 2010 8288
rect 2133 8279 2191 8285
rect 2133 8276 2145 8279
rect 2004 8248 2145 8276
rect 2004 8236 2010 8248
rect 2133 8245 2145 8248
rect 2179 8245 2191 8279
rect 7098 8276 7104 8288
rect 7059 8248 7104 8276
rect 2133 8239 2191 8245
rect 7098 8236 7104 8248
rect 7156 8236 7162 8288
rect 9030 8276 9036 8288
rect 8991 8248 9036 8276
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 19521 8279 19579 8285
rect 19521 8276 19533 8279
rect 19392 8248 19533 8276
rect 19392 8236 19398 8248
rect 19521 8245 19533 8248
rect 19567 8245 19579 8279
rect 19521 8239 19579 8245
rect 20990 8236 20996 8288
rect 21048 8276 21054 8288
rect 21177 8279 21235 8285
rect 21177 8276 21189 8279
rect 21048 8248 21189 8276
rect 21048 8236 21054 8248
rect 21177 8245 21189 8248
rect 21223 8245 21235 8279
rect 21177 8239 21235 8245
rect 1104 8186 28888 8208
rect 1104 8134 3350 8186
rect 3402 8134 3414 8186
rect 3466 8134 3478 8186
rect 3530 8134 3542 8186
rect 3594 8134 3606 8186
rect 3658 8134 8150 8186
rect 8202 8134 8214 8186
rect 8266 8134 8278 8186
rect 8330 8134 8342 8186
rect 8394 8134 8406 8186
rect 8458 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 17750 8186
rect 17802 8134 17814 8186
rect 17866 8134 17878 8186
rect 17930 8134 17942 8186
rect 17994 8134 18006 8186
rect 18058 8134 22550 8186
rect 22602 8134 22614 8186
rect 22666 8134 22678 8186
rect 22730 8134 22742 8186
rect 22794 8134 22806 8186
rect 22858 8134 27350 8186
rect 27402 8134 27414 8186
rect 27466 8134 27478 8186
rect 27530 8134 27542 8186
rect 27594 8134 27606 8186
rect 27658 8134 28888 8186
rect 1104 8112 28888 8134
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 7009 8075 7067 8081
rect 7009 8072 7021 8075
rect 5592 8044 7021 8072
rect 5592 8032 5598 8044
rect 7009 8041 7021 8044
rect 7055 8072 7067 8075
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7055 8044 7665 8072
rect 7055 8041 7067 8044
rect 7009 8035 7067 8041
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 8570 8072 8576 8084
rect 8531 8044 8576 8072
rect 7653 8035 7711 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 12618 8072 12624 8084
rect 12579 8044 12624 8072
rect 12618 8032 12624 8044
rect 12676 8072 12682 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12676 8044 13001 8072
rect 12676 8032 12682 8044
rect 12989 8041 13001 8044
rect 13035 8072 13047 8075
rect 13357 8075 13415 8081
rect 13357 8072 13369 8075
rect 13035 8044 13369 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13357 8041 13369 8044
rect 13403 8041 13415 8075
rect 20438 8072 20444 8084
rect 20399 8044 20444 8072
rect 13357 8035 13415 8041
rect 13372 8004 13400 8035
rect 20438 8032 20444 8044
rect 20496 8032 20502 8084
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 23385 8075 23443 8081
rect 23385 8072 23397 8075
rect 22152 8044 23397 8072
rect 22152 8032 22158 8044
rect 23385 8041 23397 8044
rect 23431 8041 23443 8075
rect 23385 8035 23443 8041
rect 14182 8004 14188 8016
rect 13372 7976 14188 8004
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 1946 7936 1952 7948
rect 1907 7908 1952 7936
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 7282 7936 7288 7948
rect 6687 7908 7288 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 13372 7945 13400 7976
rect 14182 7964 14188 7976
rect 14240 8004 14246 8016
rect 14829 8007 14887 8013
rect 14829 8004 14841 8007
rect 14240 7976 14841 8004
rect 14240 7964 14246 7976
rect 14829 7973 14841 7976
rect 14875 7973 14887 8007
rect 14829 7967 14887 7973
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7905 13415 7939
rect 13722 7936 13728 7948
rect 13683 7908 13728 7936
rect 13357 7899 13415 7905
rect 13722 7896 13728 7908
rect 13780 7936 13786 7948
rect 14553 7939 14611 7945
rect 14553 7936 14565 7939
rect 13780 7908 14565 7936
rect 13780 7896 13786 7908
rect 14553 7905 14565 7908
rect 14599 7905 14611 7939
rect 14553 7899 14611 7905
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7098 7868 7104 7880
rect 7055 7840 7104 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7098 7828 7104 7840
rect 7156 7868 7162 7880
rect 7650 7868 7656 7880
rect 7156 7840 7656 7868
rect 7156 7828 7162 7840
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9088 7840 9505 7868
rect 9088 7828 9094 7840
rect 9493 7837 9505 7840
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 20438 7828 20444 7880
rect 20496 7868 20502 7880
rect 20809 7871 20867 7877
rect 20809 7868 20821 7871
rect 20496 7840 20821 7868
rect 20496 7828 20502 7840
rect 20809 7837 20821 7840
rect 20855 7837 20867 7871
rect 20809 7831 20867 7837
rect 22094 7828 22100 7880
rect 22152 7868 22158 7880
rect 23201 7871 23259 7877
rect 23201 7868 23213 7871
rect 22152 7840 23213 7868
rect 22152 7828 22158 7840
rect 23201 7837 23213 7840
rect 23247 7868 23259 7871
rect 23382 7868 23388 7880
rect 23247 7840 23388 7868
rect 23247 7837 23259 7840
rect 23201 7831 23259 7837
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 3694 7800 3700 7812
rect 3174 7772 3700 7800
rect 3694 7760 3700 7772
rect 3752 7800 3758 7812
rect 9858 7800 9864 7812
rect 3752 7772 3924 7800
rect 9819 7772 9864 7800
rect 3752 7760 3758 7772
rect 3896 7744 3924 7772
rect 9858 7760 9864 7772
rect 9916 7760 9922 7812
rect 22002 7760 22008 7812
rect 22060 7800 22066 7812
rect 22833 7803 22891 7809
rect 22833 7800 22845 7803
rect 22060 7772 22845 7800
rect 22060 7760 22066 7772
rect 22833 7769 22845 7772
rect 22879 7769 22891 7803
rect 22833 7763 22891 7769
rect 23109 7803 23167 7809
rect 23109 7769 23121 7803
rect 23155 7800 23167 7803
rect 23290 7800 23296 7812
rect 23155 7772 23296 7800
rect 23155 7769 23167 7772
rect 23109 7763 23167 7769
rect 23290 7760 23296 7772
rect 23348 7760 23354 7812
rect 3418 7732 3424 7744
rect 3379 7704 3424 7732
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 3878 7732 3884 7744
rect 3839 7704 3884 7732
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 14182 7732 14188 7744
rect 14143 7704 14188 7732
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 22278 7732 22284 7744
rect 22239 7704 22284 7732
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 23014 7732 23020 7744
rect 22975 7704 23020 7732
rect 23014 7692 23020 7704
rect 23072 7692 23078 7744
rect 1104 7642 28888 7664
rect 1104 7590 5750 7642
rect 5802 7590 5814 7642
rect 5866 7590 5878 7642
rect 5930 7590 5942 7642
rect 5994 7590 6006 7642
rect 6058 7590 10550 7642
rect 10602 7590 10614 7642
rect 10666 7590 10678 7642
rect 10730 7590 10742 7642
rect 10794 7590 10806 7642
rect 10858 7590 15350 7642
rect 15402 7590 15414 7642
rect 15466 7590 15478 7642
rect 15530 7590 15542 7642
rect 15594 7590 15606 7642
rect 15658 7590 20150 7642
rect 20202 7590 20214 7642
rect 20266 7590 20278 7642
rect 20330 7590 20342 7642
rect 20394 7590 20406 7642
rect 20458 7590 24950 7642
rect 25002 7590 25014 7642
rect 25066 7590 25078 7642
rect 25130 7590 25142 7642
rect 25194 7590 25206 7642
rect 25258 7590 28888 7642
rect 1104 7568 28888 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 6089 7531 6147 7537
rect 6089 7528 6101 7531
rect 5592 7500 6101 7528
rect 5592 7488 5598 7500
rect 6089 7497 6101 7500
rect 6135 7528 6147 7531
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 6135 7500 7021 7528
rect 6135 7497 6147 7500
rect 6089 7491 6147 7497
rect 7009 7497 7021 7500
rect 7055 7528 7067 7531
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7055 7500 7665 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9732 7500 9873 7528
rect 9732 7488 9738 7500
rect 9861 7497 9873 7500
rect 9907 7528 9919 7531
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 9907 7500 10333 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 10321 7497 10333 7500
rect 10367 7528 10379 7531
rect 11057 7531 11115 7537
rect 11057 7528 11069 7531
rect 10367 7500 11069 7528
rect 10367 7497 10379 7500
rect 10321 7491 10379 7497
rect 11057 7497 11069 7500
rect 11103 7497 11115 7531
rect 11057 7491 11115 7497
rect 13909 7531 13967 7537
rect 13909 7497 13921 7531
rect 13955 7528 13967 7531
rect 14182 7528 14188 7540
rect 13955 7500 14188 7528
rect 13955 7497 13967 7500
rect 13909 7491 13967 7497
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 3418 7392 3424 7404
rect 1811 7364 3424 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 5767 7364 6653 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 6641 7361 6653 7364
rect 6687 7392 6699 7395
rect 7282 7392 7288 7404
rect 6687 7364 7288 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 11072 7401 11100 7491
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 19426 7528 19432 7540
rect 18892 7500 19432 7528
rect 18892 7460 18920 7500
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 21174 7488 21180 7540
rect 21232 7528 21238 7540
rect 21913 7531 21971 7537
rect 21913 7528 21925 7531
rect 21232 7500 21925 7528
rect 21232 7488 21238 7500
rect 21913 7497 21925 7500
rect 21959 7497 21971 7531
rect 21913 7491 21971 7497
rect 18814 7432 18920 7460
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7392 11115 7395
rect 11609 7395 11667 7401
rect 11609 7392 11621 7395
rect 11103 7364 11621 7392
rect 11103 7361 11115 7364
rect 11057 7355 11115 7361
rect 11609 7361 11621 7364
rect 11655 7361 11667 7395
rect 22186 7392 22192 7404
rect 22099 7364 22192 7392
rect 11609 7355 11667 7361
rect 22186 7352 22192 7364
rect 22244 7392 22250 7404
rect 23014 7392 23020 7404
rect 22244 7364 23020 7392
rect 22244 7352 22250 7364
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 9916 7296 10701 7324
rect 9916 7284 9922 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 19150 7324 19156 7336
rect 19111 7296 19156 7324
rect 10689 7287 10747 7293
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19521 7327 19579 7333
rect 19521 7324 19533 7327
rect 19392 7296 19533 7324
rect 19392 7284 19398 7296
rect 19521 7293 19533 7296
rect 19567 7293 19579 7327
rect 22094 7324 22100 7336
rect 22055 7296 22100 7324
rect 19521 7287 19579 7293
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7293 22339 7327
rect 22281 7287 22339 7293
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7324 22431 7327
rect 23290 7324 23296 7336
rect 22419 7296 23296 7324
rect 22419 7293 22431 7296
rect 22373 7287 22431 7293
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 7009 7259 7067 7265
rect 7009 7256 7021 7259
rect 6135 7228 7021 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 7009 7225 7021 7228
rect 7055 7256 7067 7259
rect 7650 7256 7656 7268
rect 7055 7228 7656 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 7650 7216 7656 7228
rect 7708 7216 7714 7268
rect 22002 7216 22008 7268
rect 22060 7256 22066 7268
rect 22296 7256 22324 7287
rect 23290 7284 23296 7296
rect 23348 7284 23354 7336
rect 22060 7228 22324 7256
rect 22060 7216 22066 7228
rect 17727 7191 17785 7197
rect 17727 7157 17739 7191
rect 17773 7188 17785 7191
rect 18598 7188 18604 7200
rect 17773 7160 18604 7188
rect 17773 7157 17785 7160
rect 17727 7151 17785 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 1104 7098 28888 7120
rect 1104 7046 3350 7098
rect 3402 7046 3414 7098
rect 3466 7046 3478 7098
rect 3530 7046 3542 7098
rect 3594 7046 3606 7098
rect 3658 7046 8150 7098
rect 8202 7046 8214 7098
rect 8266 7046 8278 7098
rect 8330 7046 8342 7098
rect 8394 7046 8406 7098
rect 8458 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 17750 7098
rect 17802 7046 17814 7098
rect 17866 7046 17878 7098
rect 17930 7046 17942 7098
rect 17994 7046 18006 7098
rect 18058 7046 22550 7098
rect 22602 7046 22614 7098
rect 22666 7046 22678 7098
rect 22730 7046 22742 7098
rect 22794 7046 22806 7098
rect 22858 7046 27350 7098
rect 27402 7046 27414 7098
rect 27466 7046 27478 7098
rect 27530 7046 27542 7098
rect 27594 7046 27606 7098
rect 27658 7046 28888 7098
rect 1104 7024 28888 7046
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5721 6987 5779 6993
rect 5721 6984 5733 6987
rect 5592 6956 5733 6984
rect 5592 6944 5598 6956
rect 5721 6953 5733 6956
rect 5767 6984 5779 6987
rect 6365 6987 6423 6993
rect 6365 6984 6377 6987
rect 5767 6956 6377 6984
rect 5767 6953 5779 6956
rect 5721 6947 5779 6953
rect 6365 6953 6377 6956
rect 6411 6984 6423 6987
rect 7009 6987 7067 6993
rect 7009 6984 7021 6987
rect 6411 6956 7021 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 7009 6953 7021 6956
rect 7055 6984 7067 6987
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 7055 6956 7665 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 7653 6953 7665 6956
rect 7699 6984 7711 6987
rect 8297 6987 8355 6993
rect 8297 6984 8309 6987
rect 7699 6956 8309 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 8297 6953 8309 6956
rect 8343 6984 8355 6987
rect 9674 6984 9680 6996
rect 8343 6956 9680 6984
rect 8343 6953 8355 6956
rect 8297 6947 8355 6953
rect 9674 6944 9680 6956
rect 9732 6984 9738 6996
rect 10410 6984 10416 6996
rect 9732 6956 10416 6984
rect 9732 6944 9738 6956
rect 10410 6944 10416 6956
rect 10468 6984 10474 6996
rect 11057 6987 11115 6993
rect 11057 6984 11069 6987
rect 10468 6956 11069 6984
rect 10468 6944 10474 6956
rect 11057 6953 11069 6956
rect 11103 6984 11115 6987
rect 11701 6987 11759 6993
rect 11701 6984 11713 6987
rect 11103 6956 11713 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11701 6953 11713 6956
rect 11747 6984 11759 6987
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 11747 6956 12357 6984
rect 11747 6953 11759 6956
rect 11701 6947 11759 6953
rect 12345 6953 12357 6956
rect 12391 6984 12403 6987
rect 12621 6987 12679 6993
rect 12621 6984 12633 6987
rect 12391 6956 12633 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 12621 6953 12633 6956
rect 12667 6953 12679 6987
rect 12621 6947 12679 6953
rect 18601 6987 18659 6993
rect 18601 6953 18613 6987
rect 18647 6984 18659 6987
rect 19150 6984 19156 6996
rect 18647 6956 19156 6984
rect 18647 6953 18659 6956
rect 18601 6947 18659 6953
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5997 6851 6055 6857
rect 5997 6848 6009 6851
rect 5399 6820 6009 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5997 6817 6009 6820
rect 6043 6848 6055 6851
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 6043 6820 6653 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 6641 6817 6653 6820
rect 6687 6848 6699 6851
rect 7282 6848 7288 6860
rect 6687 6820 7288 6848
rect 6687 6817 6699 6820
rect 6641 6811 6699 6817
rect 7282 6808 7288 6820
rect 7340 6848 7346 6860
rect 7929 6851 7987 6857
rect 7929 6848 7941 6851
rect 7340 6820 7941 6848
rect 7340 6808 7346 6820
rect 7929 6817 7941 6820
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 12360 6857 12388 6947
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 20990 6984 20996 6996
rect 20951 6956 20996 6984
rect 20990 6944 20996 6956
rect 21048 6944 21054 6996
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9916 6820 10057 6848
rect 9916 6808 9922 6820
rect 10045 6817 10057 6820
rect 10091 6848 10103 6851
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 10091 6820 10701 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 10689 6817 10701 6820
rect 10735 6848 10747 6851
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 10735 6820 11345 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 11333 6817 11345 6820
rect 11379 6848 11391 6851
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11379 6820 11989 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 12345 6851 12403 6857
rect 12345 6817 12357 6851
rect 12391 6817 12403 6851
rect 20990 6848 20996 6860
rect 12345 6811 12403 6817
rect 18340 6820 20996 6848
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5767 6752 6377 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 6365 6749 6377 6752
rect 6411 6780 6423 6783
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6411 6752 7021 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 7009 6749 7021 6752
rect 7055 6780 7067 6783
rect 7650 6780 7656 6792
rect 7055 6752 7656 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7650 6740 7656 6752
rect 7708 6780 7714 6792
rect 8202 6780 8208 6792
rect 7708 6752 8208 6780
rect 7708 6740 7714 6752
rect 8202 6740 8208 6752
rect 8260 6780 8266 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 8260 6752 8309 6780
rect 8260 6740 8266 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 10410 6780 10416 6792
rect 10371 6752 10416 6780
rect 8297 6743 8355 6749
rect 10410 6740 10416 6752
rect 10468 6780 10474 6792
rect 18340 6789 18368 6820
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 22094 6848 22100 6860
rect 21652 6820 22100 6848
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10468 6752 11069 6780
rect 10468 6740 10474 6752
rect 11057 6749 11069 6752
rect 11103 6780 11115 6783
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 11103 6752 11713 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18598 6780 18604 6792
rect 18559 6752 18604 6780
rect 18325 6743 18383 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 21652 6789 21680 6820
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 22278 6808 22284 6860
rect 22336 6848 22342 6860
rect 22373 6851 22431 6857
rect 22373 6848 22385 6851
rect 22336 6820 22385 6848
rect 22336 6808 22342 6820
rect 22373 6817 22385 6820
rect 22419 6817 22431 6851
rect 22373 6811 22431 6817
rect 21637 6783 21695 6789
rect 21637 6749 21649 6783
rect 21683 6749 21695 6783
rect 21637 6743 21695 6749
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6780 21971 6783
rect 22186 6780 22192 6792
rect 21959 6752 22192 6780
rect 21959 6749 21971 6752
rect 21913 6743 21971 6749
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 25225 6783 25283 6789
rect 25225 6749 25237 6783
rect 25271 6780 25283 6783
rect 25682 6780 25688 6792
rect 25271 6752 25688 6780
rect 25271 6749 25283 6752
rect 25225 6743 25283 6749
rect 25682 6740 25688 6752
rect 25740 6740 25746 6792
rect 27246 6780 27252 6792
rect 27207 6752 27252 6780
rect 27246 6740 27252 6752
rect 27304 6740 27310 6792
rect 28169 6783 28227 6789
rect 28169 6749 28181 6783
rect 28215 6780 28227 6783
rect 28258 6780 28264 6792
rect 28215 6752 28264 6780
rect 28215 6749 28227 6752
rect 28169 6743 28227 6749
rect 28258 6740 28264 6752
rect 28316 6740 28322 6792
rect 18414 6672 18420 6724
rect 18472 6712 18478 6724
rect 18509 6715 18567 6721
rect 18509 6712 18521 6715
rect 18472 6684 18521 6712
rect 18472 6672 18478 6684
rect 18509 6681 18521 6684
rect 18555 6681 18567 6715
rect 20806 6712 20812 6724
rect 20767 6684 20812 6712
rect 18509 6675 18567 6681
rect 18524 6644 18552 6675
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 21025 6715 21083 6721
rect 21025 6681 21037 6715
rect 21071 6712 21083 6715
rect 21453 6715 21511 6721
rect 21453 6712 21465 6715
rect 21071 6684 21465 6712
rect 21071 6681 21083 6684
rect 21025 6675 21083 6681
rect 21453 6681 21465 6684
rect 21499 6681 21511 6715
rect 21453 6675 21511 6681
rect 21542 6672 21548 6724
rect 21600 6712 21606 6724
rect 21821 6715 21879 6721
rect 21821 6712 21833 6715
rect 21600 6684 21833 6712
rect 21600 6672 21606 6684
rect 21821 6681 21833 6684
rect 21867 6712 21879 6715
rect 22002 6712 22008 6724
rect 21867 6684 22008 6712
rect 21867 6681 21879 6684
rect 21821 6675 21879 6681
rect 22002 6672 22008 6684
rect 22060 6672 22066 6724
rect 22646 6712 22652 6724
rect 22607 6684 22652 6712
rect 22646 6672 22652 6684
rect 22704 6672 22710 6724
rect 23934 6712 23940 6724
rect 23847 6684 23940 6712
rect 23934 6672 23940 6684
rect 23992 6712 23998 6724
rect 24578 6712 24584 6724
rect 23992 6684 24584 6712
rect 23992 6672 23998 6684
rect 24578 6672 24584 6684
rect 24636 6672 24642 6724
rect 18874 6644 18880 6656
rect 18524 6616 18880 6644
rect 18874 6604 18880 6616
rect 18932 6604 18938 6656
rect 21177 6647 21235 6653
rect 21177 6613 21189 6647
rect 21223 6644 21235 6647
rect 21634 6644 21640 6656
rect 21223 6616 21640 6644
rect 21223 6613 21235 6616
rect 21177 6607 21235 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 23382 6604 23388 6656
rect 23440 6644 23446 6656
rect 24118 6644 24124 6656
rect 23440 6616 24124 6644
rect 23440 6604 23446 6616
rect 24118 6604 24124 6616
rect 24176 6604 24182 6656
rect 25409 6647 25467 6653
rect 25409 6613 25421 6647
rect 25455 6644 25467 6647
rect 26234 6644 26240 6656
rect 25455 6616 26240 6644
rect 25455 6613 25467 6616
rect 25409 6607 25467 6613
rect 26234 6604 26240 6616
rect 26292 6604 26298 6656
rect 26878 6604 26884 6656
rect 26936 6644 26942 6656
rect 27065 6647 27123 6653
rect 27065 6644 27077 6647
rect 26936 6616 27077 6644
rect 26936 6604 26942 6616
rect 27065 6613 27077 6616
rect 27111 6613 27123 6647
rect 27065 6607 27123 6613
rect 27617 6647 27675 6653
rect 27617 6613 27629 6647
rect 27663 6644 27675 6647
rect 27798 6644 27804 6656
rect 27663 6616 27804 6644
rect 27663 6613 27675 6616
rect 27617 6607 27675 6613
rect 27798 6604 27804 6616
rect 27856 6604 27862 6656
rect 28350 6644 28356 6656
rect 28311 6616 28356 6644
rect 28350 6604 28356 6616
rect 28408 6604 28414 6656
rect 1104 6554 28888 6576
rect 1104 6502 5750 6554
rect 5802 6502 5814 6554
rect 5866 6502 5878 6554
rect 5930 6502 5942 6554
rect 5994 6502 6006 6554
rect 6058 6502 10550 6554
rect 10602 6502 10614 6554
rect 10666 6502 10678 6554
rect 10730 6502 10742 6554
rect 10794 6502 10806 6554
rect 10858 6502 15350 6554
rect 15402 6502 15414 6554
rect 15466 6502 15478 6554
rect 15530 6502 15542 6554
rect 15594 6502 15606 6554
rect 15658 6502 20150 6554
rect 20202 6502 20214 6554
rect 20266 6502 20278 6554
rect 20330 6502 20342 6554
rect 20394 6502 20406 6554
rect 20458 6502 24950 6554
rect 25002 6502 25014 6554
rect 25066 6502 25078 6554
rect 25130 6502 25142 6554
rect 25194 6502 25206 6554
rect 25258 6502 28888 6554
rect 1104 6480 28888 6502
rect 4065 6443 4123 6449
rect 4065 6409 4077 6443
rect 4111 6440 4123 6443
rect 5261 6443 5319 6449
rect 5261 6440 5273 6443
rect 4111 6412 5273 6440
rect 4111 6409 4123 6412
rect 4065 6403 4123 6409
rect 5261 6409 5273 6412
rect 5307 6440 5319 6443
rect 5534 6440 5540 6452
rect 5307 6412 5540 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 4080 6313 4108 6403
rect 5534 6400 5540 6412
rect 5592 6440 5598 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 5592 6412 6101 6440
rect 5592 6400 5598 6412
rect 6089 6409 6101 6412
rect 6135 6440 6147 6443
rect 6638 6440 6644 6452
rect 6135 6412 6644 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 6638 6400 6644 6412
rect 6696 6440 6702 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6696 6412 7021 6440
rect 6696 6400 6702 6412
rect 7009 6409 7021 6412
rect 7055 6440 7067 6443
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 7055 6412 7665 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 7653 6409 7665 6412
rect 7699 6440 7711 6443
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 7699 6412 8309 6440
rect 7699 6409 7711 6412
rect 7653 6403 7711 6409
rect 8297 6409 8309 6412
rect 8343 6440 8355 6443
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8343 6412 9045 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 9033 6409 9045 6412
rect 9079 6440 9091 6443
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 9079 6412 9413 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 9401 6403 9459 6409
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 5767 6276 6653 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 6641 6273 6653 6276
rect 6687 6304 6699 6307
rect 7282 6304 7288 6316
rect 6687 6276 7288 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 7282 6264 7288 6276
rect 7340 6304 7346 6316
rect 7650 6304 7656 6316
rect 7340 6276 7656 6304
rect 7340 6264 7346 6276
rect 7650 6264 7656 6276
rect 7708 6304 7714 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7708 6276 7941 6304
rect 7708 6264 7714 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 9416 6313 9444 6403
rect 20806 6400 20812 6452
rect 20864 6440 20870 6452
rect 21085 6443 21143 6449
rect 21085 6440 21097 6443
rect 20864 6412 21097 6440
rect 20864 6400 20870 6412
rect 21085 6409 21097 6412
rect 21131 6409 21143 6443
rect 22186 6440 22192 6452
rect 21085 6403 21143 6409
rect 21192 6412 22192 6440
rect 21192 6381 21220 6412
rect 22186 6400 22192 6412
rect 22244 6400 22250 6452
rect 22373 6443 22431 6449
rect 22373 6409 22385 6443
rect 22419 6440 22431 6443
rect 22646 6440 22652 6452
rect 22419 6412 22652 6440
rect 22419 6409 22431 6412
rect 22373 6403 22431 6409
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 27246 6440 27252 6452
rect 27207 6412 27252 6440
rect 27246 6400 27252 6412
rect 27304 6400 27310 6452
rect 21177 6375 21235 6381
rect 21177 6372 21189 6375
rect 19720 6344 21189 6372
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 8260 6276 8309 6304
rect 8260 6264 8266 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9769 6307 9827 6313
rect 9447 6276 9674 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4479 6208 4721 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4709 6205 4721 6208
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 6089 6171 6147 6177
rect 6089 6137 6101 6171
rect 6135 6168 6147 6171
rect 7009 6171 7067 6177
rect 7009 6168 7021 6171
rect 6135 6140 7021 6168
rect 6135 6137 6147 6140
rect 6089 6131 6147 6137
rect 7009 6137 7021 6140
rect 7055 6168 7067 6171
rect 7282 6168 7288 6180
rect 7055 6140 7288 6168
rect 7055 6137 7067 6140
rect 7009 6131 7067 6137
rect 7282 6128 7288 6140
rect 7340 6168 7346 6180
rect 7653 6171 7711 6177
rect 7653 6168 7665 6171
rect 7340 6140 7665 6168
rect 7340 6128 7346 6140
rect 7653 6137 7665 6140
rect 7699 6168 7711 6171
rect 8220 6168 8248 6264
rect 9646 6236 9674 6276
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 9858 6304 9864 6316
rect 9815 6276 9864 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 9858 6264 9864 6276
rect 9916 6304 9922 6316
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9916 6276 10057 6304
rect 9916 6264 9922 6276
rect 10045 6273 10057 6276
rect 10091 6304 10103 6307
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10091 6276 10701 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 10689 6273 10701 6276
rect 10735 6304 10747 6307
rect 11609 6307 11667 6313
rect 11609 6304 11621 6307
rect 10735 6276 11621 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 11609 6273 11621 6276
rect 11655 6304 11667 6307
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 11655 6276 12265 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 12253 6273 12265 6276
rect 12299 6304 12311 6307
rect 12621 6307 12679 6313
rect 12299 6276 12572 6304
rect 12299 6273 12311 6276
rect 12253 6267 12311 6273
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 9646 6208 10425 6236
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6205 12035 6239
rect 12544 6236 12572 6276
rect 12621 6273 12633 6307
rect 12667 6304 12679 6307
rect 12667 6276 13308 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 13280 6245 13308 6276
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 19242 6304 19248 6316
rect 18656 6276 19248 6304
rect 18656 6264 18662 6276
rect 19242 6264 19248 6276
rect 19300 6304 19306 6316
rect 19720 6313 19748 6344
rect 21177 6341 21189 6344
rect 21223 6341 21235 6375
rect 21177 6335 21235 6341
rect 21361 6375 21419 6381
rect 21361 6341 21373 6375
rect 21407 6372 21419 6375
rect 22094 6372 22100 6384
rect 21407 6344 22100 6372
rect 21407 6341 21419 6344
rect 21361 6335 21419 6341
rect 22094 6332 22100 6344
rect 22152 6332 22158 6384
rect 26234 6332 26240 6384
rect 26292 6372 26298 6384
rect 27617 6375 27675 6381
rect 27617 6372 27629 6375
rect 26292 6344 27629 6372
rect 26292 6332 26298 6344
rect 27617 6341 27629 6344
rect 27663 6341 27675 6375
rect 27617 6335 27675 6341
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 19300 6276 19717 6304
rect 19300 6264 19306 6276
rect 19705 6273 19717 6276
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6304 19855 6307
rect 20714 6304 20720 6316
rect 19843 6276 20720 6304
rect 19843 6273 19855 6276
rect 19797 6267 19855 6273
rect 20714 6264 20720 6276
rect 20772 6304 20778 6316
rect 21085 6307 21143 6313
rect 21085 6304 21097 6307
rect 20772 6276 21097 6304
rect 20772 6264 20778 6276
rect 21085 6273 21097 6276
rect 21131 6304 21143 6307
rect 21542 6304 21548 6316
rect 21131 6276 21548 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 21542 6264 21548 6276
rect 21600 6264 21606 6316
rect 21634 6264 21640 6316
rect 21692 6304 21698 6316
rect 22189 6307 22247 6313
rect 22189 6304 22201 6307
rect 21692 6276 22201 6304
rect 21692 6264 21698 6276
rect 22189 6273 22201 6276
rect 22235 6273 22247 6307
rect 22189 6267 22247 6273
rect 24578 6264 24584 6316
rect 24636 6304 24642 6316
rect 24636 6290 25162 6304
rect 24636 6276 25176 6290
rect 24636 6264 24642 6276
rect 12897 6239 12955 6245
rect 12897 6236 12909 6239
rect 12544 6208 12909 6236
rect 11977 6199 12035 6205
rect 12897 6205 12909 6208
rect 12943 6205 12955 6239
rect 12897 6199 12955 6205
rect 13265 6239 13323 6245
rect 13265 6205 13277 6239
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6236 19579 6239
rect 20990 6236 20996 6248
rect 19567 6208 20996 6236
rect 19567 6205 19579 6208
rect 19521 6199 19579 6205
rect 7699 6140 8248 6168
rect 7699 6137 7711 6140
rect 7653 6131 7711 6137
rect 10428 6109 10456 6199
rect 11072 6109 11100 6199
rect 11992 6109 12020 6199
rect 10413 6103 10471 6109
rect 10413 6069 10425 6103
rect 10459 6100 10471 6103
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 10459 6072 11069 6100
rect 10459 6069 10471 6072
rect 10413 6063 10471 6069
rect 11057 6069 11069 6072
rect 11103 6100 11115 6103
rect 11977 6103 12035 6109
rect 11977 6100 11989 6103
rect 11103 6072 11989 6100
rect 11103 6069 11115 6072
rect 11057 6063 11115 6069
rect 11977 6069 11989 6072
rect 12023 6100 12035 6103
rect 12618 6100 12624 6112
rect 12023 6072 12624 6100
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 12618 6060 12624 6072
rect 12676 6100 12682 6112
rect 13280 6109 13308 6199
rect 20990 6196 20996 6208
rect 21048 6196 21054 6248
rect 25148 6236 25176 6276
rect 26513 6239 26571 6245
rect 25148 6208 26464 6236
rect 13265 6103 13323 6109
rect 13265 6100 13277 6103
rect 12676 6072 13277 6100
rect 12676 6060 12682 6072
rect 13265 6069 13277 6072
rect 13311 6100 13323 6103
rect 13541 6103 13599 6109
rect 13541 6100 13553 6103
rect 13311 6072 13553 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 13541 6069 13553 6072
rect 13587 6069 13599 6103
rect 13541 6063 13599 6069
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 19613 6103 19671 6109
rect 19613 6100 19625 6103
rect 19576 6072 19625 6100
rect 19576 6060 19582 6072
rect 19613 6069 19625 6072
rect 19659 6069 19671 6103
rect 19613 6063 19671 6069
rect 24765 6103 24823 6109
rect 24765 6069 24777 6103
rect 24811 6100 24823 6103
rect 25222 6100 25228 6112
rect 24811 6072 25228 6100
rect 24811 6069 24823 6072
rect 24765 6063 24823 6069
rect 25222 6060 25228 6072
rect 25280 6060 25286 6112
rect 26436 6100 26464 6208
rect 26513 6205 26525 6239
rect 26559 6236 26571 6239
rect 26602 6236 26608 6248
rect 26559 6208 26608 6236
rect 26559 6205 26571 6208
rect 26513 6199 26571 6205
rect 26602 6196 26608 6208
rect 26660 6196 26666 6248
rect 27709 6239 27767 6245
rect 27709 6205 27721 6239
rect 27755 6205 27767 6239
rect 27709 6199 27767 6205
rect 27724 6168 27752 6199
rect 27798 6196 27804 6248
rect 27856 6236 27862 6248
rect 27856 6208 27901 6236
rect 27856 6196 27862 6208
rect 28350 6168 28356 6180
rect 27724 6140 28356 6168
rect 28350 6128 28356 6140
rect 28408 6128 28414 6180
rect 27890 6100 27896 6112
rect 26436 6072 27896 6100
rect 27890 6060 27896 6072
rect 27948 6060 27954 6112
rect 1104 6010 28888 6032
rect 1104 5958 3350 6010
rect 3402 5958 3414 6010
rect 3466 5958 3478 6010
rect 3530 5958 3542 6010
rect 3594 5958 3606 6010
rect 3658 5958 8150 6010
rect 8202 5958 8214 6010
rect 8266 5958 8278 6010
rect 8330 5958 8342 6010
rect 8394 5958 8406 6010
rect 8458 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 17750 6010
rect 17802 5958 17814 6010
rect 17866 5958 17878 6010
rect 17930 5958 17942 6010
rect 17994 5958 18006 6010
rect 18058 5958 22550 6010
rect 22602 5958 22614 6010
rect 22666 5958 22678 6010
rect 22730 5958 22742 6010
rect 22794 5958 22806 6010
rect 22858 5958 27350 6010
rect 27402 5958 27414 6010
rect 27466 5958 27478 6010
rect 27530 5958 27542 6010
rect 27594 5958 27606 6010
rect 27658 5958 28888 6010
rect 1104 5936 28888 5958
rect 9309 5899 9367 5905
rect 9309 5865 9321 5899
rect 9355 5896 9367 5899
rect 12345 5899 12403 5905
rect 9355 5868 9812 5896
rect 9355 5865 9367 5868
rect 9309 5859 9367 5865
rect 6641 5831 6699 5837
rect 6641 5797 6653 5831
rect 6687 5828 6699 5831
rect 7282 5828 7288 5840
rect 6687 5800 7288 5828
rect 6687 5797 6699 5800
rect 6641 5791 6699 5797
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 7650 5760 7656 5772
rect 7055 5732 7656 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 9784 5633 9812 5868
rect 12345 5865 12357 5899
rect 12391 5896 12403 5899
rect 12618 5896 12624 5908
rect 12391 5868 12624 5896
rect 12391 5865 12403 5868
rect 12345 5859 12403 5865
rect 11698 5828 11704 5840
rect 11611 5800 11704 5828
rect 11698 5788 11704 5800
rect 11756 5828 11762 5840
rect 12360 5828 12388 5859
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 24670 5896 24676 5908
rect 24631 5868 24676 5896
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 25682 5896 25688 5908
rect 25643 5868 25688 5896
rect 25682 5856 25688 5868
rect 25740 5856 25746 5908
rect 28350 5896 28356 5908
rect 28311 5868 28356 5896
rect 28350 5856 28356 5868
rect 28408 5856 28414 5908
rect 11756 5800 12388 5828
rect 11756 5788 11762 5800
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9916 5732 10057 5760
rect 9916 5720 9922 5732
rect 10045 5729 10057 5732
rect 10091 5760 10103 5763
rect 10689 5763 10747 5769
rect 10689 5760 10701 5763
rect 10091 5732 10701 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 10689 5729 10701 5732
rect 10735 5760 10747 5763
rect 10962 5760 10968 5772
rect 10735 5732 10968 5760
rect 10735 5729 10747 5732
rect 10689 5723 10747 5729
rect 10962 5720 10968 5732
rect 11020 5760 11026 5772
rect 12360 5769 12388 5800
rect 19337 5831 19395 5837
rect 19337 5797 19349 5831
rect 19383 5828 19395 5831
rect 19426 5828 19432 5840
rect 19383 5800 19432 5828
rect 19383 5797 19395 5800
rect 19337 5791 19395 5797
rect 19426 5788 19432 5800
rect 19484 5788 19490 5840
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11020 5732 11345 5760
rect 11020 5720 11026 5732
rect 11333 5729 11345 5732
rect 11379 5760 11391 5763
rect 11977 5763 12035 5769
rect 11977 5760 11989 5763
rect 11379 5732 11989 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 11977 5729 11989 5732
rect 12023 5729 12035 5763
rect 11977 5723 12035 5729
rect 12345 5763 12403 5769
rect 12345 5729 12357 5763
rect 12391 5729 12403 5763
rect 12345 5723 12403 5729
rect 19242 5720 19248 5772
rect 19300 5760 19306 5772
rect 24688 5760 24716 5856
rect 25041 5763 25099 5769
rect 25041 5760 25053 5763
rect 19300 5732 19656 5760
rect 24688 5732 25053 5760
rect 19300 5720 19306 5732
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 10459 5664 11069 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 11057 5661 11069 5664
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 19337 5695 19395 5701
rect 19337 5661 19349 5695
rect 19383 5692 19395 5695
rect 19518 5692 19524 5704
rect 19383 5664 19524 5692
rect 19383 5661 19395 5664
rect 19337 5655 19395 5661
rect 9769 5627 9827 5633
rect 9769 5593 9781 5627
rect 9815 5624 9827 5627
rect 10428 5624 10456 5655
rect 9815 5596 10456 5624
rect 9815 5593 9827 5596
rect 9769 5587 9827 5593
rect 6638 5556 6644 5568
rect 6599 5528 6644 5556
rect 6638 5516 6644 5528
rect 6696 5556 6702 5568
rect 10428 5565 10456 5596
rect 11072 5565 11100 5655
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 19628 5701 19656 5732
rect 25041 5729 25053 5732
rect 25087 5729 25099 5763
rect 25222 5760 25228 5772
rect 25183 5732 25228 5760
rect 25041 5723 25099 5729
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 26878 5760 26884 5772
rect 26839 5732 26884 5760
rect 26878 5720 26884 5732
rect 26936 5720 26942 5772
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 24118 5652 24124 5704
rect 24176 5692 24182 5704
rect 25317 5695 25375 5701
rect 25317 5692 25329 5695
rect 24176 5664 25329 5692
rect 24176 5652 24182 5664
rect 25317 5661 25329 5664
rect 25363 5661 25375 5695
rect 26602 5692 26608 5704
rect 26563 5664 26608 5692
rect 25317 5655 25375 5661
rect 26602 5652 26608 5664
rect 26660 5652 26666 5704
rect 27890 5584 27896 5636
rect 27948 5584 27954 5636
rect 7285 5559 7343 5565
rect 7285 5556 7297 5559
rect 6696 5528 7297 5556
rect 6696 5516 6702 5528
rect 7285 5525 7297 5528
rect 7331 5525 7343 5559
rect 7285 5519 7343 5525
rect 10413 5559 10471 5565
rect 10413 5525 10425 5559
rect 10459 5525 10471 5559
rect 10413 5519 10471 5525
rect 11057 5559 11115 5565
rect 11057 5525 11069 5559
rect 11103 5556 11115 5559
rect 11698 5556 11704 5568
rect 11103 5528 11704 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 19521 5559 19579 5565
rect 19521 5525 19533 5559
rect 19567 5556 19579 5559
rect 20714 5556 20720 5568
rect 19567 5528 20720 5556
rect 19567 5525 19579 5528
rect 19521 5519 19579 5525
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 1104 5466 28888 5488
rect 1104 5414 5750 5466
rect 5802 5414 5814 5466
rect 5866 5414 5878 5466
rect 5930 5414 5942 5466
rect 5994 5414 6006 5466
rect 6058 5414 10550 5466
rect 10602 5414 10614 5466
rect 10666 5414 10678 5466
rect 10730 5414 10742 5466
rect 10794 5414 10806 5466
rect 10858 5414 15350 5466
rect 15402 5414 15414 5466
rect 15466 5414 15478 5466
rect 15530 5414 15542 5466
rect 15594 5414 15606 5466
rect 15658 5414 20150 5466
rect 20202 5414 20214 5466
rect 20266 5414 20278 5466
rect 20330 5414 20342 5466
rect 20394 5414 20406 5466
rect 20458 5414 24950 5466
rect 25002 5414 25014 5466
rect 25066 5414 25078 5466
rect 25130 5414 25142 5466
rect 25194 5414 25206 5466
rect 25258 5414 28888 5466
rect 1104 5392 28888 5414
rect 9953 5355 10011 5361
rect 9953 5321 9965 5355
rect 9999 5352 10011 5355
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 9999 5324 10425 5352
rect 9999 5321 10011 5324
rect 9953 5315 10011 5321
rect 10413 5321 10425 5324
rect 10459 5352 10471 5355
rect 10689 5355 10747 5361
rect 10689 5352 10701 5355
rect 10459 5324 10701 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 10689 5321 10701 5324
rect 10735 5352 10747 5355
rect 11698 5352 11704 5364
rect 10735 5324 11704 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 10704 5225 10732 5315
rect 11698 5312 11704 5324
rect 11756 5352 11762 5364
rect 11977 5355 12035 5361
rect 11977 5352 11989 5355
rect 11756 5324 11989 5352
rect 11756 5312 11762 5324
rect 11977 5321 11989 5324
rect 12023 5321 12035 5355
rect 11977 5315 12035 5321
rect 20533 5355 20591 5361
rect 20533 5321 20545 5355
rect 20579 5352 20591 5355
rect 20714 5352 20720 5364
rect 20579 5324 20720 5352
rect 20579 5321 20591 5324
rect 20533 5315 20591 5321
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 19334 5284 19340 5296
rect 18800 5256 19340 5284
rect 10689 5219 10747 5225
rect 10689 5216 10701 5219
rect 10652 5188 10701 5216
rect 10652 5176 10658 5188
rect 10689 5185 10701 5188
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 18800 5225 18828 5256
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 19610 5244 19616 5296
rect 19668 5244 19674 5296
rect 11057 5219 11115 5225
rect 11057 5216 11069 5219
rect 11020 5188 11069 5216
rect 11020 5176 11026 5188
rect 11057 5185 11069 5188
rect 11103 5185 11115 5219
rect 11057 5179 11115 5185
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 19061 5151 19119 5157
rect 19061 5117 19073 5151
rect 19107 5148 19119 5151
rect 19426 5148 19432 5160
rect 19107 5120 19432 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 23017 5015 23075 5021
rect 23017 4981 23029 5015
rect 23063 5012 23075 5015
rect 23566 5012 23572 5024
rect 23063 4984 23572 5012
rect 23063 4981 23075 4984
rect 23017 4975 23075 4981
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 1104 4922 28888 4944
rect 1104 4870 3350 4922
rect 3402 4870 3414 4922
rect 3466 4870 3478 4922
rect 3530 4870 3542 4922
rect 3594 4870 3606 4922
rect 3658 4870 8150 4922
rect 8202 4870 8214 4922
rect 8266 4870 8278 4922
rect 8330 4870 8342 4922
rect 8394 4870 8406 4922
rect 8458 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 17750 4922
rect 17802 4870 17814 4922
rect 17866 4870 17878 4922
rect 17930 4870 17942 4922
rect 17994 4870 18006 4922
rect 18058 4870 22550 4922
rect 22602 4870 22614 4922
rect 22666 4870 22678 4922
rect 22730 4870 22742 4922
rect 22794 4870 22806 4922
rect 22858 4870 27350 4922
rect 27402 4870 27414 4922
rect 27466 4870 27478 4922
rect 27530 4870 27542 4922
rect 27594 4870 27606 4922
rect 27658 4870 28888 4922
rect 1104 4848 28888 4870
rect 10594 4808 10600 4820
rect 10555 4780 10600 4808
rect 10594 4768 10600 4780
rect 10652 4808 10658 4820
rect 11149 4811 11207 4817
rect 11149 4808 11161 4811
rect 10652 4780 11161 4808
rect 10652 4768 10658 4780
rect 11149 4777 11161 4780
rect 11195 4777 11207 4811
rect 11149 4771 11207 4777
rect 21821 4675 21879 4681
rect 21821 4641 21833 4675
rect 21867 4672 21879 4675
rect 22741 4675 22799 4681
rect 22741 4672 22753 4675
rect 21867 4644 22753 4672
rect 21867 4641 21879 4644
rect 21821 4635 21879 4641
rect 22741 4641 22753 4644
rect 22787 4672 22799 4675
rect 23566 4672 23572 4684
rect 22787 4644 23572 4672
rect 22787 4641 22799 4644
rect 22741 4635 22799 4641
rect 23566 4632 23572 4644
rect 23624 4672 23630 4684
rect 23753 4675 23811 4681
rect 23753 4672 23765 4675
rect 23624 4644 23765 4672
rect 23624 4632 23630 4644
rect 23753 4641 23765 4644
rect 23799 4672 23811 4675
rect 24670 4672 24676 4684
rect 23799 4644 24676 4672
rect 23799 4641 23811 4644
rect 23753 4635 23811 4641
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 22465 4607 22523 4613
rect 22465 4604 22477 4607
rect 20772 4576 22477 4604
rect 20772 4564 20778 4576
rect 22465 4573 22477 4576
rect 22511 4573 22523 4607
rect 22465 4567 22523 4573
rect 23014 4564 23020 4616
rect 23072 4604 23078 4616
rect 23477 4607 23535 4613
rect 23477 4604 23489 4607
rect 23072 4576 23489 4604
rect 23072 4564 23078 4576
rect 23477 4573 23489 4576
rect 23523 4573 23535 4607
rect 23477 4567 23535 4573
rect 26234 4564 26240 4616
rect 26292 4604 26298 4616
rect 26602 4604 26608 4616
rect 26292 4576 26608 4604
rect 26292 4564 26298 4576
rect 26602 4564 26608 4576
rect 26660 4604 26666 4616
rect 26697 4607 26755 4613
rect 26697 4604 26709 4607
rect 26660 4576 26709 4604
rect 26660 4564 26666 4576
rect 26697 4573 26709 4576
rect 26743 4573 26755 4607
rect 26697 4567 26755 4573
rect 26970 4536 26976 4548
rect 26931 4508 26976 4536
rect 26970 4496 26976 4508
rect 27028 4496 27034 4548
rect 27982 4496 27988 4548
rect 28040 4496 28046 4548
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3329 4471 3387 4477
rect 3329 4468 3341 4471
rect 3200 4440 3341 4468
rect 3200 4428 3206 4440
rect 3329 4437 3341 4440
rect 3375 4437 3387 4471
rect 22094 4468 22100 4480
rect 22055 4440 22100 4468
rect 3329 4431 3387 4437
rect 22094 4428 22100 4440
rect 22152 4428 22158 4480
rect 22557 4471 22615 4477
rect 22557 4437 22569 4471
rect 22603 4468 22615 4471
rect 23014 4468 23020 4480
rect 22603 4440 23020 4468
rect 22603 4437 22615 4440
rect 22557 4431 22615 4437
rect 23014 4428 23020 4440
rect 23072 4428 23078 4480
rect 23109 4471 23167 4477
rect 23109 4437 23121 4471
rect 23155 4468 23167 4471
rect 23198 4468 23204 4480
rect 23155 4440 23204 4468
rect 23155 4437 23167 4440
rect 23109 4431 23167 4437
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 23566 4428 23572 4480
rect 23624 4468 23630 4480
rect 28442 4468 28448 4480
rect 23624 4440 23669 4468
rect 28403 4440 28448 4468
rect 23624 4428 23630 4440
rect 28442 4428 28448 4440
rect 28500 4428 28506 4480
rect 1104 4378 28888 4400
rect 1104 4326 5750 4378
rect 5802 4326 5814 4378
rect 5866 4326 5878 4378
rect 5930 4326 5942 4378
rect 5994 4326 6006 4378
rect 6058 4326 10550 4378
rect 10602 4326 10614 4378
rect 10666 4326 10678 4378
rect 10730 4326 10742 4378
rect 10794 4326 10806 4378
rect 10858 4326 15350 4378
rect 15402 4326 15414 4378
rect 15466 4326 15478 4378
rect 15530 4326 15542 4378
rect 15594 4326 15606 4378
rect 15658 4326 20150 4378
rect 20202 4326 20214 4378
rect 20266 4326 20278 4378
rect 20330 4326 20342 4378
rect 20394 4326 20406 4378
rect 20458 4326 24950 4378
rect 25002 4326 25014 4378
rect 25066 4326 25078 4378
rect 25130 4326 25142 4378
rect 25194 4326 25206 4378
rect 25258 4326 28888 4378
rect 1104 4304 28888 4326
rect 2869 4267 2927 4273
rect 2869 4233 2881 4267
rect 2915 4264 2927 4267
rect 10226 4264 10232 4276
rect 2915 4236 10232 4264
rect 2915 4233 2927 4236
rect 2869 4227 2927 4233
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 27709 4267 27767 4273
rect 27709 4233 27721 4267
rect 27755 4264 27767 4267
rect 28442 4264 28448 4276
rect 27755 4236 28448 4264
rect 27755 4233 27767 4236
rect 27709 4227 27767 4233
rect 28442 4224 28448 4236
rect 28500 4224 28506 4276
rect 3881 4199 3939 4205
rect 3881 4165 3893 4199
rect 3927 4196 3939 4199
rect 11606 4196 11612 4208
rect 3927 4168 11612 4196
rect 3927 4165 3939 4168
rect 3881 4159 3939 4165
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 19610 4156 19616 4208
rect 19668 4196 19674 4208
rect 20070 4196 20076 4208
rect 19668 4168 20076 4196
rect 19668 4156 19674 4168
rect 20070 4156 20076 4168
rect 20128 4196 20134 4208
rect 22557 4199 22615 4205
rect 22557 4196 22569 4199
rect 20128 4168 22569 4196
rect 20128 4156 20134 4168
rect 22557 4165 22569 4168
rect 22603 4165 22615 4199
rect 22557 4159 22615 4165
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4128 20591 4131
rect 21082 4128 21088 4140
rect 20579 4100 21088 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 22094 4128 22100 4140
rect 22051 4100 22100 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 23198 4128 23204 4140
rect 23159 4100 23204 4128
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 25406 4128 25412 4140
rect 25367 4100 25412 4128
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 27617 4131 27675 4137
rect 27617 4128 27629 4131
rect 26206 4100 27629 4128
rect 2958 4060 2964 4072
rect 2919 4032 2964 4060
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3142 4060 3148 4072
rect 3103 4032 3148 4060
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 26206 4060 26234 4100
rect 27617 4097 27629 4100
rect 27663 4097 27675 4131
rect 27617 4091 27675 4097
rect 22204 4032 26234 4060
rect 26697 4063 26755 4069
rect 21634 3952 21640 4004
rect 21692 3992 21698 4004
rect 22204 4001 22232 4032
rect 26697 4029 26709 4063
rect 26743 4060 26755 4063
rect 27798 4060 27804 4072
rect 26743 4032 27804 4060
rect 26743 4029 26755 4032
rect 26697 4023 26755 4029
rect 27798 4020 27804 4032
rect 27856 4020 27862 4072
rect 22189 3995 22247 4001
rect 22189 3992 22201 3995
rect 21692 3964 22201 3992
rect 21692 3952 21698 3964
rect 22189 3961 22201 3964
rect 22235 3961 22247 3995
rect 23382 3992 23388 4004
rect 23295 3964 23388 3992
rect 22189 3955 22247 3961
rect 23382 3952 23388 3964
rect 23440 3992 23446 4004
rect 25774 3992 25780 4004
rect 23440 3964 25780 3992
rect 23440 3952 23446 3964
rect 25774 3952 25780 3964
rect 25832 3952 25838 4004
rect 2498 3924 2504 3936
rect 2459 3896 2504 3924
rect 2498 3884 2504 3896
rect 2556 3884 2562 3936
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 3789 3927 3847 3933
rect 3789 3924 3801 3927
rect 3752 3896 3801 3924
rect 3752 3884 3758 3896
rect 3789 3893 3801 3896
rect 3835 3893 3847 3927
rect 3789 3887 3847 3893
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 18840 3896 20453 3924
rect 18840 3884 18846 3896
rect 20441 3893 20453 3896
rect 20487 3893 20499 3927
rect 20441 3887 20499 3893
rect 22833 3927 22891 3933
rect 22833 3893 22845 3927
rect 22879 3924 22891 3927
rect 23842 3924 23848 3936
rect 22879 3896 23848 3924
rect 22879 3893 22891 3896
rect 22833 3887 22891 3893
rect 23842 3884 23848 3896
rect 23900 3884 23906 3936
rect 25130 3884 25136 3936
rect 25188 3924 25194 3936
rect 25225 3927 25283 3933
rect 25225 3924 25237 3927
rect 25188 3896 25237 3924
rect 25188 3884 25194 3896
rect 25225 3893 25237 3896
rect 25271 3893 25283 3927
rect 27246 3924 27252 3936
rect 27207 3896 27252 3924
rect 25225 3887 25283 3893
rect 27246 3884 27252 3896
rect 27304 3884 27310 3936
rect 1104 3834 28888 3856
rect 1104 3782 3350 3834
rect 3402 3782 3414 3834
rect 3466 3782 3478 3834
rect 3530 3782 3542 3834
rect 3594 3782 3606 3834
rect 3658 3782 8150 3834
rect 8202 3782 8214 3834
rect 8266 3782 8278 3834
rect 8330 3782 8342 3834
rect 8394 3782 8406 3834
rect 8458 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 17750 3834
rect 17802 3782 17814 3834
rect 17866 3782 17878 3834
rect 17930 3782 17942 3834
rect 17994 3782 18006 3834
rect 18058 3782 22550 3834
rect 22602 3782 22614 3834
rect 22666 3782 22678 3834
rect 22730 3782 22742 3834
rect 22794 3782 22806 3834
rect 22858 3782 27350 3834
rect 27402 3782 27414 3834
rect 27466 3782 27478 3834
rect 27530 3782 27542 3834
rect 27594 3782 27606 3834
rect 27658 3782 28888 3834
rect 1104 3760 28888 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3016 3692 3433 3720
rect 3016 3680 3022 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 21082 3720 21088 3732
rect 21043 3692 21088 3720
rect 3421 3683 3479 3689
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 23014 3680 23020 3732
rect 23072 3720 23078 3732
rect 23109 3723 23167 3729
rect 23109 3720 23121 3723
rect 23072 3692 23121 3720
rect 23072 3680 23078 3692
rect 23109 3689 23121 3692
rect 23155 3689 23167 3723
rect 23109 3683 23167 3689
rect 26970 3680 26976 3732
rect 27028 3720 27034 3732
rect 27065 3723 27123 3729
rect 27065 3720 27077 3723
rect 27028 3692 27077 3720
rect 27028 3680 27034 3692
rect 27065 3689 27077 3692
rect 27111 3689 27123 3723
rect 28350 3720 28356 3732
rect 28311 3692 28356 3720
rect 27065 3683 27123 3689
rect 28350 3680 28356 3692
rect 28408 3680 28414 3732
rect 26234 3652 26240 3664
rect 26206 3612 26240 3652
rect 26292 3612 26298 3664
rect 1670 3584 1676 3596
rect 1631 3556 1676 3584
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 3786 3544 3792 3596
rect 3844 3584 3850 3596
rect 13814 3584 13820 3596
rect 3844 3556 13820 3584
rect 3844 3544 3850 3556
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3584 18751 3587
rect 19334 3584 19340 3596
rect 18739 3556 19104 3584
rect 19247 3556 19340 3584
rect 18739 3553 18751 3556
rect 18693 3547 18751 3553
rect 3050 3476 3056 3528
rect 3108 3516 3114 3528
rect 3878 3516 3884 3528
rect 3108 3488 3884 3516
rect 3108 3476 3114 3488
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 18506 3516 18512 3528
rect 18467 3488 18512 3516
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 18782 3516 18788 3528
rect 18743 3488 18788 3516
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 18874 3476 18880 3528
rect 18932 3525 18938 3528
rect 18932 3516 18940 3525
rect 18932 3488 18977 3516
rect 18932 3479 18940 3488
rect 18932 3476 18938 3479
rect 1949 3451 2007 3457
rect 1949 3417 1961 3451
rect 1995 3448 2007 3451
rect 2222 3448 2228 3460
rect 1995 3420 2228 3448
rect 1995 3417 2007 3420
rect 1949 3411 2007 3417
rect 2222 3408 2228 3420
rect 2280 3408 2286 3460
rect 18230 3448 18236 3460
rect 18143 3420 18236 3448
rect 18230 3408 18236 3420
rect 18288 3448 18294 3460
rect 18693 3451 18751 3457
rect 18693 3448 18705 3451
rect 18288 3420 18705 3448
rect 18288 3408 18294 3420
rect 18693 3417 18705 3420
rect 18739 3417 18751 3451
rect 19076 3448 19104 3556
rect 19334 3544 19340 3556
rect 19392 3584 19398 3596
rect 21361 3587 21419 3593
rect 21361 3584 21373 3587
rect 19392 3556 21373 3584
rect 19392 3544 19398 3556
rect 21361 3553 21373 3556
rect 21407 3553 21419 3587
rect 21634 3584 21640 3596
rect 21595 3556 21640 3584
rect 21361 3547 21419 3553
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 22278 3544 22284 3596
rect 22336 3584 22342 3596
rect 24857 3587 24915 3593
rect 24857 3584 24869 3587
rect 22336 3556 24869 3584
rect 22336 3544 22342 3556
rect 24857 3553 24869 3556
rect 24903 3584 24915 3587
rect 26206 3584 26234 3612
rect 24903 3556 26234 3584
rect 24903 3553 24915 3556
rect 24857 3547 24915 3553
rect 27246 3516 27252 3528
rect 27207 3488 27252 3516
rect 27246 3476 27252 3488
rect 27304 3476 27310 3528
rect 28169 3519 28227 3525
rect 28169 3485 28181 3519
rect 28215 3516 28227 3519
rect 28442 3516 28448 3528
rect 28215 3488 28448 3516
rect 28215 3485 28227 3488
rect 28169 3479 28227 3485
rect 28442 3476 28448 3488
rect 28500 3476 28506 3528
rect 19613 3451 19671 3457
rect 19613 3448 19625 3451
rect 19076 3420 19625 3448
rect 18693 3411 18751 3417
rect 19613 3417 19625 3420
rect 19659 3417 19671 3451
rect 19613 3411 19671 3417
rect 20070 3408 20076 3460
rect 20128 3408 20134 3460
rect 23842 3448 23848 3460
rect 22862 3420 23848 3448
rect 23842 3408 23848 3420
rect 23900 3408 23906 3460
rect 25130 3448 25136 3460
rect 25091 3420 25136 3448
rect 25130 3408 25136 3420
rect 25188 3408 25194 3460
rect 26418 3448 26424 3460
rect 26331 3420 26424 3448
rect 26418 3408 26424 3420
rect 26476 3448 26482 3460
rect 27890 3448 27896 3460
rect 26476 3420 27896 3448
rect 26476 3408 26482 3420
rect 27890 3408 27896 3420
rect 27948 3408 27954 3460
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 2958 3380 2964 3392
rect 1820 3352 2964 3380
rect 1820 3340 1826 3352
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 21082 3340 21088 3392
rect 21140 3380 21146 3392
rect 26142 3380 26148 3392
rect 21140 3352 26148 3380
rect 21140 3340 21146 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 26602 3380 26608 3392
rect 26563 3352 26608 3380
rect 26602 3340 26608 3352
rect 26660 3340 26666 3392
rect 1104 3290 28888 3312
rect 1104 3238 5750 3290
rect 5802 3238 5814 3290
rect 5866 3238 5878 3290
rect 5930 3238 5942 3290
rect 5994 3238 6006 3290
rect 6058 3238 10550 3290
rect 10602 3238 10614 3290
rect 10666 3238 10678 3290
rect 10730 3238 10742 3290
rect 10794 3238 10806 3290
rect 10858 3238 15350 3290
rect 15402 3238 15414 3290
rect 15466 3238 15478 3290
rect 15530 3238 15542 3290
rect 15594 3238 15606 3290
rect 15658 3238 20150 3290
rect 20202 3238 20214 3290
rect 20266 3238 20278 3290
rect 20330 3238 20342 3290
rect 20394 3238 20406 3290
rect 20458 3238 24950 3290
rect 25002 3238 25014 3290
rect 25066 3238 25078 3290
rect 25130 3238 25142 3290
rect 25194 3238 25206 3290
rect 25258 3238 28888 3290
rect 1104 3216 28888 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3050 3176 3056 3188
rect 3007 3148 3056 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 19702 3176 19708 3188
rect 19663 3148 19708 3176
rect 19702 3136 19708 3148
rect 19760 3176 19766 3188
rect 23382 3176 23388 3188
rect 19760 3148 20484 3176
rect 19760 3136 19766 3148
rect 20070 3108 20076 3120
rect 20031 3080 20076 3108
rect 20070 3068 20076 3080
rect 20128 3068 20134 3120
rect 20456 3117 20484 3148
rect 22572 3148 23388 3176
rect 22572 3117 22600 3148
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 23566 3136 23572 3188
rect 23624 3176 23630 3188
rect 24029 3179 24087 3185
rect 24029 3176 24041 3179
rect 23624 3148 24041 3176
rect 23624 3136 23630 3148
rect 24029 3145 24041 3148
rect 24075 3145 24087 3179
rect 25406 3176 25412 3188
rect 25367 3148 25412 3176
rect 24029 3139 24087 3145
rect 25406 3136 25412 3148
rect 25464 3136 25470 3188
rect 25774 3176 25780 3188
rect 25735 3148 25780 3176
rect 25774 3136 25780 3148
rect 25832 3136 25838 3188
rect 20441 3111 20499 3117
rect 20441 3077 20453 3111
rect 20487 3077 20499 3111
rect 20441 3071 20499 3077
rect 22557 3111 22615 3117
rect 22557 3077 22569 3111
rect 22603 3077 22615 3111
rect 23842 3108 23848 3120
rect 23755 3080 23848 3108
rect 22557 3071 22615 3077
rect 23842 3068 23848 3080
rect 23900 3108 23906 3120
rect 26418 3108 26424 3120
rect 23900 3080 26424 3108
rect 23900 3068 23906 3080
rect 26418 3068 26424 3080
rect 26476 3068 26482 3120
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2498 3040 2504 3052
rect 2455 3012 2504 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 3694 3040 3700 3052
rect 3283 3012 3700 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 22278 3040 22284 3052
rect 22239 3012 22284 3040
rect 22278 3000 22284 3012
rect 22336 3000 22342 3052
rect 25869 3043 25927 3049
rect 25869 3009 25881 3043
rect 25915 3040 25927 3043
rect 26602 3040 26608 3052
rect 25915 3012 26608 3040
rect 25915 3009 25927 3012
rect 25869 3003 25927 3009
rect 26602 3000 26608 3012
rect 26660 3000 26666 3052
rect 3712 2913 3740 3000
rect 18417 2975 18475 2981
rect 18417 2941 18429 2975
rect 18463 2972 18475 2975
rect 18874 2972 18880 2984
rect 18463 2944 18880 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 18874 2932 18880 2944
rect 18932 2972 18938 2984
rect 25133 2975 25191 2981
rect 25133 2972 25145 2975
rect 18932 2944 25145 2972
rect 18932 2932 18938 2944
rect 25133 2941 25145 2944
rect 25179 2972 25191 2975
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 25179 2944 25973 2972
rect 25179 2941 25191 2944
rect 25133 2935 25191 2941
rect 25961 2941 25973 2944
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 3697 2907 3755 2913
rect 3697 2873 3709 2907
rect 3743 2904 3755 2907
rect 19702 2904 19708 2916
rect 3743 2876 19708 2904
rect 3743 2873 3755 2876
rect 3697 2867 3755 2873
rect 19702 2864 19708 2876
rect 19760 2864 19766 2916
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 1104 2746 28888 2768
rect 1104 2694 3350 2746
rect 3402 2694 3414 2746
rect 3466 2694 3478 2746
rect 3530 2694 3542 2746
rect 3594 2694 3606 2746
rect 3658 2694 8150 2746
rect 8202 2694 8214 2746
rect 8266 2694 8278 2746
rect 8330 2694 8342 2746
rect 8394 2694 8406 2746
rect 8458 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 17750 2746
rect 17802 2694 17814 2746
rect 17866 2694 17878 2746
rect 17930 2694 17942 2746
rect 17994 2694 18006 2746
rect 18058 2694 22550 2746
rect 22602 2694 22614 2746
rect 22666 2694 22678 2746
rect 22730 2694 22742 2746
rect 22794 2694 22806 2746
rect 22858 2694 27350 2746
rect 27402 2694 27414 2746
rect 27466 2694 27478 2746
rect 27530 2694 27542 2746
rect 27594 2694 27606 2746
rect 27658 2694 28888 2746
rect 1104 2672 28888 2694
rect 11606 2632 11612 2644
rect 11567 2604 11612 2632
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 18506 2592 18512 2644
rect 18564 2632 18570 2644
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 18564 2604 18797 2632
rect 18564 2592 18570 2604
rect 18785 2601 18797 2604
rect 18831 2601 18843 2635
rect 18785 2595 18843 2601
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11296 2400 11805 2428
rect 11296 2388 11302 2400
rect 11793 2397 11805 2400
rect 11839 2428 11851 2431
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 11839 2400 12081 2428
rect 11839 2397 11851 2400
rect 11793 2391 11851 2397
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 18969 2431 19027 2437
rect 18969 2428 18981 2431
rect 18748 2400 18981 2428
rect 18748 2388 18754 2400
rect 18969 2397 18981 2400
rect 19015 2428 19027 2431
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 19015 2400 19349 2428
rect 19015 2397 19027 2400
rect 18969 2391 19027 2397
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 19337 2391 19395 2397
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 26292 2400 26337 2428
rect 26292 2388 26298 2400
rect 26602 2388 26608 2440
rect 26660 2428 26666 2440
rect 28169 2431 28227 2437
rect 28169 2428 28181 2431
rect 26660 2400 28181 2428
rect 26660 2388 26666 2400
rect 28169 2397 28181 2400
rect 28215 2397 28227 2431
rect 28169 2391 28227 2397
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 26421 2295 26479 2301
rect 26421 2292 26433 2295
rect 26200 2264 26433 2292
rect 26200 2252 26206 2264
rect 26421 2261 26433 2264
rect 26467 2261 26479 2295
rect 28350 2292 28356 2304
rect 28311 2264 28356 2292
rect 26421 2255 26479 2261
rect 28350 2252 28356 2264
rect 28408 2252 28414 2304
rect 1104 2202 28888 2224
rect 1104 2150 5750 2202
rect 5802 2150 5814 2202
rect 5866 2150 5878 2202
rect 5930 2150 5942 2202
rect 5994 2150 6006 2202
rect 6058 2150 10550 2202
rect 10602 2150 10614 2202
rect 10666 2150 10678 2202
rect 10730 2150 10742 2202
rect 10794 2150 10806 2202
rect 10858 2150 15350 2202
rect 15402 2150 15414 2202
rect 15466 2150 15478 2202
rect 15530 2150 15542 2202
rect 15594 2150 15606 2202
rect 15658 2150 20150 2202
rect 20202 2150 20214 2202
rect 20266 2150 20278 2202
rect 20330 2150 20342 2202
rect 20394 2150 20406 2202
rect 20458 2150 24950 2202
rect 25002 2150 25014 2202
rect 25066 2150 25078 2202
rect 25130 2150 25142 2202
rect 25194 2150 25206 2202
rect 25258 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3350 27718 3402 27770
rect 3414 27718 3466 27770
rect 3478 27718 3530 27770
rect 3542 27718 3594 27770
rect 3606 27718 3658 27770
rect 8150 27718 8202 27770
rect 8214 27718 8266 27770
rect 8278 27718 8330 27770
rect 8342 27718 8394 27770
rect 8406 27718 8458 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 17750 27718 17802 27770
rect 17814 27718 17866 27770
rect 17878 27718 17930 27770
rect 17942 27718 17994 27770
rect 18006 27718 18058 27770
rect 22550 27718 22602 27770
rect 22614 27718 22666 27770
rect 22678 27718 22730 27770
rect 22742 27718 22794 27770
rect 22806 27718 22858 27770
rect 27350 27718 27402 27770
rect 27414 27718 27466 27770
rect 27478 27718 27530 27770
rect 27542 27718 27594 27770
rect 27606 27718 27658 27770
rect 28356 27591 28408 27600
rect 28356 27557 28365 27591
rect 28365 27557 28399 27591
rect 28399 27557 28408 27591
rect 28356 27548 28408 27557
rect 3056 27412 3108 27464
rect 27804 27412 27856 27464
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 5750 27174 5802 27226
rect 5814 27174 5866 27226
rect 5878 27174 5930 27226
rect 5942 27174 5994 27226
rect 6006 27174 6058 27226
rect 10550 27174 10602 27226
rect 10614 27174 10666 27226
rect 10678 27174 10730 27226
rect 10742 27174 10794 27226
rect 10806 27174 10858 27226
rect 15350 27174 15402 27226
rect 15414 27174 15466 27226
rect 15478 27174 15530 27226
rect 15542 27174 15594 27226
rect 15606 27174 15658 27226
rect 20150 27174 20202 27226
rect 20214 27174 20266 27226
rect 20278 27174 20330 27226
rect 20342 27174 20394 27226
rect 20406 27174 20458 27226
rect 24950 27174 25002 27226
rect 25014 27174 25066 27226
rect 25078 27174 25130 27226
rect 25142 27174 25194 27226
rect 25206 27174 25258 27226
rect 3350 26630 3402 26682
rect 3414 26630 3466 26682
rect 3478 26630 3530 26682
rect 3542 26630 3594 26682
rect 3606 26630 3658 26682
rect 8150 26630 8202 26682
rect 8214 26630 8266 26682
rect 8278 26630 8330 26682
rect 8342 26630 8394 26682
rect 8406 26630 8458 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 17750 26630 17802 26682
rect 17814 26630 17866 26682
rect 17878 26630 17930 26682
rect 17942 26630 17994 26682
rect 18006 26630 18058 26682
rect 22550 26630 22602 26682
rect 22614 26630 22666 26682
rect 22678 26630 22730 26682
rect 22742 26630 22794 26682
rect 22806 26630 22858 26682
rect 27350 26630 27402 26682
rect 27414 26630 27466 26682
rect 27478 26630 27530 26682
rect 27542 26630 27594 26682
rect 27606 26630 27658 26682
rect 28356 26503 28408 26512
rect 28356 26469 28365 26503
rect 28365 26469 28399 26503
rect 28399 26469 28408 26503
rect 28356 26460 28408 26469
rect 27712 26324 27764 26376
rect 5750 26086 5802 26138
rect 5814 26086 5866 26138
rect 5878 26086 5930 26138
rect 5942 26086 5994 26138
rect 6006 26086 6058 26138
rect 10550 26086 10602 26138
rect 10614 26086 10666 26138
rect 10678 26086 10730 26138
rect 10742 26086 10794 26138
rect 10806 26086 10858 26138
rect 15350 26086 15402 26138
rect 15414 26086 15466 26138
rect 15478 26086 15530 26138
rect 15542 26086 15594 26138
rect 15606 26086 15658 26138
rect 20150 26086 20202 26138
rect 20214 26086 20266 26138
rect 20278 26086 20330 26138
rect 20342 26086 20394 26138
rect 20406 26086 20458 26138
rect 24950 26086 25002 26138
rect 25014 26086 25066 26138
rect 25078 26086 25130 26138
rect 25142 26086 25194 26138
rect 25206 26086 25258 26138
rect 3350 25542 3402 25594
rect 3414 25542 3466 25594
rect 3478 25542 3530 25594
rect 3542 25542 3594 25594
rect 3606 25542 3658 25594
rect 8150 25542 8202 25594
rect 8214 25542 8266 25594
rect 8278 25542 8330 25594
rect 8342 25542 8394 25594
rect 8406 25542 8458 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 17750 25542 17802 25594
rect 17814 25542 17866 25594
rect 17878 25542 17930 25594
rect 17942 25542 17994 25594
rect 18006 25542 18058 25594
rect 22550 25542 22602 25594
rect 22614 25542 22666 25594
rect 22678 25542 22730 25594
rect 22742 25542 22794 25594
rect 22806 25542 22858 25594
rect 27350 25542 27402 25594
rect 27414 25542 27466 25594
rect 27478 25542 27530 25594
rect 27542 25542 27594 25594
rect 27606 25542 27658 25594
rect 5750 24998 5802 25050
rect 5814 24998 5866 25050
rect 5878 24998 5930 25050
rect 5942 24998 5994 25050
rect 6006 24998 6058 25050
rect 10550 24998 10602 25050
rect 10614 24998 10666 25050
rect 10678 24998 10730 25050
rect 10742 24998 10794 25050
rect 10806 24998 10858 25050
rect 15350 24998 15402 25050
rect 15414 24998 15466 25050
rect 15478 24998 15530 25050
rect 15542 24998 15594 25050
rect 15606 24998 15658 25050
rect 20150 24998 20202 25050
rect 20214 24998 20266 25050
rect 20278 24998 20330 25050
rect 20342 24998 20394 25050
rect 20406 24998 20458 25050
rect 24950 24998 25002 25050
rect 25014 24998 25066 25050
rect 25078 24998 25130 25050
rect 25142 24998 25194 25050
rect 25206 24998 25258 25050
rect 3350 24454 3402 24506
rect 3414 24454 3466 24506
rect 3478 24454 3530 24506
rect 3542 24454 3594 24506
rect 3606 24454 3658 24506
rect 8150 24454 8202 24506
rect 8214 24454 8266 24506
rect 8278 24454 8330 24506
rect 8342 24454 8394 24506
rect 8406 24454 8458 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 17750 24454 17802 24506
rect 17814 24454 17866 24506
rect 17878 24454 17930 24506
rect 17942 24454 17994 24506
rect 18006 24454 18058 24506
rect 22550 24454 22602 24506
rect 22614 24454 22666 24506
rect 22678 24454 22730 24506
rect 22742 24454 22794 24506
rect 22806 24454 22858 24506
rect 27350 24454 27402 24506
rect 27414 24454 27466 24506
rect 27478 24454 27530 24506
rect 27542 24454 27594 24506
rect 27606 24454 27658 24506
rect 5750 23910 5802 23962
rect 5814 23910 5866 23962
rect 5878 23910 5930 23962
rect 5942 23910 5994 23962
rect 6006 23910 6058 23962
rect 10550 23910 10602 23962
rect 10614 23910 10666 23962
rect 10678 23910 10730 23962
rect 10742 23910 10794 23962
rect 10806 23910 10858 23962
rect 15350 23910 15402 23962
rect 15414 23910 15466 23962
rect 15478 23910 15530 23962
rect 15542 23910 15594 23962
rect 15606 23910 15658 23962
rect 20150 23910 20202 23962
rect 20214 23910 20266 23962
rect 20278 23910 20330 23962
rect 20342 23910 20394 23962
rect 20406 23910 20458 23962
rect 24950 23910 25002 23962
rect 25014 23910 25066 23962
rect 25078 23910 25130 23962
rect 25142 23910 25194 23962
rect 25206 23910 25258 23962
rect 24216 23672 24268 23724
rect 28356 23511 28408 23520
rect 28356 23477 28365 23511
rect 28365 23477 28399 23511
rect 28399 23477 28408 23511
rect 28356 23468 28408 23477
rect 3350 23366 3402 23418
rect 3414 23366 3466 23418
rect 3478 23366 3530 23418
rect 3542 23366 3594 23418
rect 3606 23366 3658 23418
rect 8150 23366 8202 23418
rect 8214 23366 8266 23418
rect 8278 23366 8330 23418
rect 8342 23366 8394 23418
rect 8406 23366 8458 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 17750 23366 17802 23418
rect 17814 23366 17866 23418
rect 17878 23366 17930 23418
rect 17942 23366 17994 23418
rect 18006 23366 18058 23418
rect 22550 23366 22602 23418
rect 22614 23366 22666 23418
rect 22678 23366 22730 23418
rect 22742 23366 22794 23418
rect 22806 23366 22858 23418
rect 27350 23366 27402 23418
rect 27414 23366 27466 23418
rect 27478 23366 27530 23418
rect 27542 23366 27594 23418
rect 27606 23366 27658 23418
rect 5750 22822 5802 22874
rect 5814 22822 5866 22874
rect 5878 22822 5930 22874
rect 5942 22822 5994 22874
rect 6006 22822 6058 22874
rect 10550 22822 10602 22874
rect 10614 22822 10666 22874
rect 10678 22822 10730 22874
rect 10742 22822 10794 22874
rect 10806 22822 10858 22874
rect 15350 22822 15402 22874
rect 15414 22822 15466 22874
rect 15478 22822 15530 22874
rect 15542 22822 15594 22874
rect 15606 22822 15658 22874
rect 20150 22822 20202 22874
rect 20214 22822 20266 22874
rect 20278 22822 20330 22874
rect 20342 22822 20394 22874
rect 20406 22822 20458 22874
rect 24950 22822 25002 22874
rect 25014 22822 25066 22874
rect 25078 22822 25130 22874
rect 25142 22822 25194 22874
rect 25206 22822 25258 22874
rect 24216 22720 24268 22772
rect 23480 22652 23532 22704
rect 3148 22584 3200 22636
rect 25872 22627 25924 22636
rect 25872 22593 25881 22627
rect 25881 22593 25915 22627
rect 25915 22593 25924 22627
rect 25872 22584 25924 22593
rect 26608 22448 26660 22500
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 24124 22380 24176 22432
rect 25688 22423 25740 22432
rect 25688 22389 25697 22423
rect 25697 22389 25731 22423
rect 25731 22389 25740 22423
rect 25688 22380 25740 22389
rect 3350 22278 3402 22330
rect 3414 22278 3466 22330
rect 3478 22278 3530 22330
rect 3542 22278 3594 22330
rect 3606 22278 3658 22330
rect 8150 22278 8202 22330
rect 8214 22278 8266 22330
rect 8278 22278 8330 22330
rect 8342 22278 8394 22330
rect 8406 22278 8458 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 17750 22278 17802 22330
rect 17814 22278 17866 22330
rect 17878 22278 17930 22330
rect 17942 22278 17994 22330
rect 18006 22278 18058 22330
rect 22550 22278 22602 22330
rect 22614 22278 22666 22330
rect 22678 22278 22730 22330
rect 22742 22278 22794 22330
rect 22806 22278 22858 22330
rect 27350 22278 27402 22330
rect 27414 22278 27466 22330
rect 27478 22278 27530 22330
rect 27542 22278 27594 22330
rect 27606 22278 27658 22330
rect 23940 22176 23992 22228
rect 24216 22176 24268 22228
rect 25688 22176 25740 22228
rect 19156 22040 19208 22092
rect 23664 22040 23716 22092
rect 27620 22040 27672 22092
rect 27804 22083 27856 22092
rect 27804 22049 27813 22083
rect 27813 22049 27847 22083
rect 27847 22049 27856 22083
rect 27804 22040 27856 22049
rect 19984 21972 20036 22024
rect 25320 22015 25372 22024
rect 25320 21981 25329 22015
rect 25329 21981 25363 22015
rect 25363 21981 25372 22015
rect 25320 21972 25372 21981
rect 27344 21972 27396 22024
rect 26056 21904 26108 21956
rect 19432 21836 19484 21888
rect 26332 21836 26384 21888
rect 27252 21836 27304 21888
rect 27712 21879 27764 21888
rect 27712 21845 27721 21879
rect 27721 21845 27755 21879
rect 27755 21845 27764 21879
rect 27712 21836 27764 21845
rect 5750 21734 5802 21786
rect 5814 21734 5866 21786
rect 5878 21734 5930 21786
rect 5942 21734 5994 21786
rect 6006 21734 6058 21786
rect 10550 21734 10602 21786
rect 10614 21734 10666 21786
rect 10678 21734 10730 21786
rect 10742 21734 10794 21786
rect 10806 21734 10858 21786
rect 15350 21734 15402 21786
rect 15414 21734 15466 21786
rect 15478 21734 15530 21786
rect 15542 21734 15594 21786
rect 15606 21734 15658 21786
rect 20150 21734 20202 21786
rect 20214 21734 20266 21786
rect 20278 21734 20330 21786
rect 20342 21734 20394 21786
rect 20406 21734 20458 21786
rect 24950 21734 25002 21786
rect 25014 21734 25066 21786
rect 25078 21734 25130 21786
rect 25142 21734 25194 21786
rect 25206 21734 25258 21786
rect 3056 21632 3108 21684
rect 18236 21632 18288 21684
rect 23940 21675 23992 21684
rect 2780 21564 2832 21616
rect 19432 21607 19484 21616
rect 19432 21573 19441 21607
rect 19441 21573 19475 21607
rect 19475 21573 19484 21607
rect 19432 21564 19484 21573
rect 19524 21564 19576 21616
rect 23480 21564 23532 21616
rect 23940 21641 23949 21675
rect 23949 21641 23983 21675
rect 23983 21641 23992 21675
rect 23940 21632 23992 21641
rect 25872 21632 25924 21684
rect 26332 21675 26384 21684
rect 26332 21641 26341 21675
rect 26341 21641 26375 21675
rect 26375 21641 26384 21675
rect 26332 21632 26384 21641
rect 27620 21632 27672 21684
rect 27712 21564 27764 21616
rect 19156 21539 19208 21548
rect 19156 21505 19165 21539
rect 19165 21505 19199 21539
rect 19199 21505 19208 21539
rect 19156 21496 19208 21505
rect 24124 21539 24176 21548
rect 1768 21428 1820 21480
rect 2136 21471 2188 21480
rect 2136 21437 2145 21471
rect 2145 21437 2179 21471
rect 2179 21437 2188 21471
rect 2136 21428 2188 21437
rect 19524 21428 19576 21480
rect 24124 21505 24133 21539
rect 24133 21505 24167 21539
rect 24167 21505 24176 21539
rect 24124 21496 24176 21505
rect 27252 21539 27304 21548
rect 27252 21505 27261 21539
rect 27261 21505 27295 21539
rect 27295 21505 27304 21539
rect 27252 21496 27304 21505
rect 28172 21539 28224 21548
rect 28172 21505 28181 21539
rect 28181 21505 28215 21539
rect 28215 21505 28224 21539
rect 28172 21496 28224 21505
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 26608 21471 26660 21480
rect 23664 21428 23716 21437
rect 26608 21437 26617 21471
rect 26617 21437 26651 21471
rect 26651 21437 26660 21471
rect 26608 21428 26660 21437
rect 26332 21360 26384 21412
rect 27252 21360 27304 21412
rect 20444 21292 20496 21344
rect 22376 21292 22428 21344
rect 26608 21292 26660 21344
rect 28356 21335 28408 21344
rect 28356 21301 28365 21335
rect 28365 21301 28399 21335
rect 28399 21301 28408 21335
rect 28356 21292 28408 21301
rect 3350 21190 3402 21242
rect 3414 21190 3466 21242
rect 3478 21190 3530 21242
rect 3542 21190 3594 21242
rect 3606 21190 3658 21242
rect 8150 21190 8202 21242
rect 8214 21190 8266 21242
rect 8278 21190 8330 21242
rect 8342 21190 8394 21242
rect 8406 21190 8458 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 17750 21190 17802 21242
rect 17814 21190 17866 21242
rect 17878 21190 17930 21242
rect 17942 21190 17994 21242
rect 18006 21190 18058 21242
rect 22550 21190 22602 21242
rect 22614 21190 22666 21242
rect 22678 21190 22730 21242
rect 22742 21190 22794 21242
rect 22806 21190 22858 21242
rect 27350 21190 27402 21242
rect 27414 21190 27466 21242
rect 27478 21190 27530 21242
rect 27542 21190 27594 21242
rect 27606 21190 27658 21242
rect 3148 21088 3200 21140
rect 19984 21131 20036 21140
rect 1768 20995 1820 21004
rect 1768 20961 1777 20995
rect 1777 20961 1811 20995
rect 1811 20961 1820 20995
rect 1768 20952 1820 20961
rect 3240 20952 3292 21004
rect 19984 21097 19993 21131
rect 19993 21097 20027 21131
rect 20027 21097 20036 21131
rect 19984 21088 20036 21097
rect 23480 21088 23532 21140
rect 27804 21088 27856 21140
rect 4896 20952 4948 21004
rect 20444 20995 20496 21004
rect 20444 20961 20453 20995
rect 20453 20961 20487 20995
rect 20487 20961 20496 20995
rect 20444 20952 20496 20961
rect 20720 20952 20772 21004
rect 26608 20995 26660 21004
rect 26608 20961 26617 20995
rect 26617 20961 26651 20995
rect 26651 20961 26660 20995
rect 26608 20952 26660 20961
rect 16856 20927 16908 20936
rect 16856 20893 16865 20927
rect 16865 20893 16899 20927
rect 16899 20893 16908 20927
rect 16856 20884 16908 20893
rect 22008 20927 22060 20936
rect 22008 20893 22017 20927
rect 22017 20893 22051 20927
rect 22051 20893 22060 20927
rect 22008 20884 22060 20893
rect 26332 20927 26384 20936
rect 26332 20893 26341 20927
rect 26341 20893 26375 20927
rect 26375 20893 26384 20927
rect 26332 20884 26384 20893
rect 2044 20859 2096 20868
rect 2044 20825 2053 20859
rect 2053 20825 2087 20859
rect 2087 20825 2096 20859
rect 2044 20816 2096 20825
rect 2780 20816 2832 20868
rect 6736 20816 6788 20868
rect 26056 20859 26108 20868
rect 26056 20825 26065 20859
rect 26065 20825 26099 20859
rect 26099 20825 26108 20859
rect 26056 20816 26108 20825
rect 3884 20791 3936 20800
rect 3884 20757 3893 20791
rect 3893 20757 3927 20791
rect 3927 20757 3936 20791
rect 3884 20748 3936 20757
rect 4896 20791 4948 20800
rect 4896 20757 4905 20791
rect 4905 20757 4939 20791
rect 4939 20757 4948 20791
rect 4896 20748 4948 20757
rect 18236 20748 18288 20800
rect 19524 20748 19576 20800
rect 5750 20646 5802 20698
rect 5814 20646 5866 20698
rect 5878 20646 5930 20698
rect 5942 20646 5994 20698
rect 6006 20646 6058 20698
rect 10550 20646 10602 20698
rect 10614 20646 10666 20698
rect 10678 20646 10730 20698
rect 10742 20646 10794 20698
rect 10806 20646 10858 20698
rect 15350 20646 15402 20698
rect 15414 20646 15466 20698
rect 15478 20646 15530 20698
rect 15542 20646 15594 20698
rect 15606 20646 15658 20698
rect 20150 20646 20202 20698
rect 20214 20646 20266 20698
rect 20278 20646 20330 20698
rect 20342 20646 20394 20698
rect 20406 20646 20458 20698
rect 24950 20646 25002 20698
rect 25014 20646 25066 20698
rect 25078 20646 25130 20698
rect 25142 20646 25194 20698
rect 25206 20646 25258 20698
rect 2136 20544 2188 20596
rect 3056 20544 3108 20596
rect 22008 20544 22060 20596
rect 22376 20587 22428 20596
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 18236 20519 18288 20528
rect 18236 20485 18245 20519
rect 18245 20485 18279 20519
rect 18279 20485 18288 20519
rect 18236 20476 18288 20485
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 17132 20408 17184 20460
rect 19156 20408 19208 20460
rect 19800 20408 19852 20460
rect 21272 20408 21324 20460
rect 28172 20544 28224 20596
rect 4896 20340 4948 20392
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 24308 20340 24360 20392
rect 24860 20340 24912 20392
rect 27252 20272 27304 20324
rect 3792 20247 3844 20256
rect 3792 20213 3801 20247
rect 3801 20213 3835 20247
rect 3835 20213 3844 20247
rect 3792 20204 3844 20213
rect 16764 20247 16816 20256
rect 16764 20213 16773 20247
rect 16773 20213 16807 20247
rect 16807 20213 16816 20247
rect 16764 20204 16816 20213
rect 26424 20204 26476 20256
rect 3350 20102 3402 20154
rect 3414 20102 3466 20154
rect 3478 20102 3530 20154
rect 3542 20102 3594 20154
rect 3606 20102 3658 20154
rect 8150 20102 8202 20154
rect 8214 20102 8266 20154
rect 8278 20102 8330 20154
rect 8342 20102 8394 20154
rect 8406 20102 8458 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 17750 20102 17802 20154
rect 17814 20102 17866 20154
rect 17878 20102 17930 20154
rect 17942 20102 17994 20154
rect 18006 20102 18058 20154
rect 22550 20102 22602 20154
rect 22614 20102 22666 20154
rect 22678 20102 22730 20154
rect 22742 20102 22794 20154
rect 22806 20102 22858 20154
rect 27350 20102 27402 20154
rect 27414 20102 27466 20154
rect 27478 20102 27530 20154
rect 27542 20102 27594 20154
rect 27606 20102 27658 20154
rect 2044 20000 2096 20052
rect 16856 20043 16908 20052
rect 16856 20009 16865 20043
rect 16865 20009 16899 20043
rect 16899 20009 16908 20043
rect 16856 20000 16908 20009
rect 22468 20000 22520 20052
rect 28172 20000 28224 20052
rect 16764 19864 16816 19916
rect 17408 19907 17460 19916
rect 17408 19873 17417 19907
rect 17417 19873 17451 19907
rect 17451 19873 17460 19907
rect 17408 19864 17460 19873
rect 20720 19864 20772 19916
rect 3884 19796 3936 19848
rect 23296 19864 23348 19916
rect 25320 19864 25372 19916
rect 26424 19907 26476 19916
rect 26424 19873 26433 19907
rect 26433 19873 26467 19907
rect 26467 19873 26476 19907
rect 26424 19864 26476 19873
rect 17500 19660 17552 19712
rect 26240 19660 26292 19712
rect 27712 19660 27764 19712
rect 5750 19558 5802 19610
rect 5814 19558 5866 19610
rect 5878 19558 5930 19610
rect 5942 19558 5994 19610
rect 6006 19558 6058 19610
rect 10550 19558 10602 19610
rect 10614 19558 10666 19610
rect 10678 19558 10730 19610
rect 10742 19558 10794 19610
rect 10806 19558 10858 19610
rect 15350 19558 15402 19610
rect 15414 19558 15466 19610
rect 15478 19558 15530 19610
rect 15542 19558 15594 19610
rect 15606 19558 15658 19610
rect 20150 19558 20202 19610
rect 20214 19558 20266 19610
rect 20278 19558 20330 19610
rect 20342 19558 20394 19610
rect 20406 19558 20458 19610
rect 24950 19558 25002 19610
rect 25014 19558 25066 19610
rect 25078 19558 25130 19610
rect 25142 19558 25194 19610
rect 25206 19558 25258 19610
rect 16580 19388 16632 19440
rect 17132 19388 17184 19440
rect 19340 19456 19392 19508
rect 19524 19499 19576 19508
rect 19524 19465 19533 19499
rect 19533 19465 19567 19499
rect 19567 19465 19576 19499
rect 19524 19456 19576 19465
rect 17224 19320 17276 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 18144 19252 18196 19304
rect 24860 19252 24912 19304
rect 24952 19116 25004 19168
rect 3350 19014 3402 19066
rect 3414 19014 3466 19066
rect 3478 19014 3530 19066
rect 3542 19014 3594 19066
rect 3606 19014 3658 19066
rect 8150 19014 8202 19066
rect 8214 19014 8266 19066
rect 8278 19014 8330 19066
rect 8342 19014 8394 19066
rect 8406 19014 8458 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 17750 19014 17802 19066
rect 17814 19014 17866 19066
rect 17878 19014 17930 19066
rect 17942 19014 17994 19066
rect 18006 19014 18058 19066
rect 22550 19014 22602 19066
rect 22614 19014 22666 19066
rect 22678 19014 22730 19066
rect 22742 19014 22794 19066
rect 22806 19014 22858 19066
rect 27350 19014 27402 19066
rect 27414 19014 27466 19066
rect 27478 19014 27530 19066
rect 27542 19014 27594 19066
rect 27606 19014 27658 19066
rect 6736 18955 6788 18964
rect 6736 18921 6745 18955
rect 6745 18921 6779 18955
rect 6779 18921 6788 18955
rect 6736 18912 6788 18921
rect 18144 18912 18196 18964
rect 24860 18912 24912 18964
rect 21272 18819 21324 18828
rect 21272 18785 21281 18819
rect 21281 18785 21315 18819
rect 21315 18785 21324 18819
rect 21272 18776 21324 18785
rect 3240 18708 3292 18760
rect 18788 18708 18840 18760
rect 24952 18819 25004 18828
rect 24952 18785 24961 18819
rect 24961 18785 24995 18819
rect 24995 18785 25004 18819
rect 24952 18776 25004 18785
rect 5264 18683 5316 18692
rect 5264 18649 5273 18683
rect 5273 18649 5307 18683
rect 5307 18649 5316 18683
rect 5264 18640 5316 18649
rect 2780 18572 2832 18624
rect 3976 18572 4028 18624
rect 21548 18640 21600 18692
rect 28172 18751 28224 18760
rect 28172 18717 28181 18751
rect 28181 18717 28215 18751
rect 28215 18717 28224 18751
rect 28172 18708 28224 18717
rect 8300 18572 8352 18624
rect 20904 18615 20956 18624
rect 20904 18581 20913 18615
rect 20913 18581 20947 18615
rect 20947 18581 20956 18615
rect 20904 18572 20956 18581
rect 24308 18572 24360 18624
rect 28356 18615 28408 18624
rect 28356 18581 28365 18615
rect 28365 18581 28399 18615
rect 28399 18581 28408 18615
rect 28356 18572 28408 18581
rect 5750 18470 5802 18522
rect 5814 18470 5866 18522
rect 5878 18470 5930 18522
rect 5942 18470 5994 18522
rect 6006 18470 6058 18522
rect 10550 18470 10602 18522
rect 10614 18470 10666 18522
rect 10678 18470 10730 18522
rect 10742 18470 10794 18522
rect 10806 18470 10858 18522
rect 15350 18470 15402 18522
rect 15414 18470 15466 18522
rect 15478 18470 15530 18522
rect 15542 18470 15594 18522
rect 15606 18470 15658 18522
rect 20150 18470 20202 18522
rect 20214 18470 20266 18522
rect 20278 18470 20330 18522
rect 20342 18470 20394 18522
rect 20406 18470 20458 18522
rect 24950 18470 25002 18522
rect 25014 18470 25066 18522
rect 25078 18470 25130 18522
rect 25142 18470 25194 18522
rect 25206 18470 25258 18522
rect 3148 18368 3200 18420
rect 4068 18368 4120 18420
rect 21364 18368 21416 18420
rect 24308 18411 24360 18420
rect 24308 18377 24317 18411
rect 24317 18377 24351 18411
rect 24351 18377 24360 18411
rect 24308 18368 24360 18377
rect 2780 18300 2832 18352
rect 7380 18300 7432 18352
rect 8300 18300 8352 18352
rect 19340 18300 19392 18352
rect 20536 18300 20588 18352
rect 2228 18275 2280 18284
rect 2228 18241 2237 18275
rect 2237 18241 2271 18275
rect 2271 18241 2280 18275
rect 2228 18232 2280 18241
rect 19800 18275 19852 18284
rect 19800 18241 19809 18275
rect 19809 18241 19843 18275
rect 19843 18241 19852 18275
rect 19800 18232 19852 18241
rect 4436 18207 4488 18216
rect 4436 18173 4445 18207
rect 4445 18173 4479 18207
rect 4479 18173 4488 18207
rect 4436 18164 4488 18173
rect 2872 18028 2924 18080
rect 3240 18028 3292 18080
rect 20628 18164 20680 18216
rect 24860 18164 24912 18216
rect 28172 18232 28224 18284
rect 27252 18096 27304 18148
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 5080 18028 5132 18037
rect 9128 18071 9180 18080
rect 9128 18037 9137 18071
rect 9137 18037 9171 18071
rect 9171 18037 9180 18071
rect 9128 18028 9180 18037
rect 20536 18028 20588 18080
rect 21180 18028 21232 18080
rect 26608 18028 26660 18080
rect 3350 17926 3402 17978
rect 3414 17926 3466 17978
rect 3478 17926 3530 17978
rect 3542 17926 3594 17978
rect 3606 17926 3658 17978
rect 8150 17926 8202 17978
rect 8214 17926 8266 17978
rect 8278 17926 8330 17978
rect 8342 17926 8394 17978
rect 8406 17926 8458 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 17750 17926 17802 17978
rect 17814 17926 17866 17978
rect 17878 17926 17930 17978
rect 17942 17926 17994 17978
rect 18006 17926 18058 17978
rect 22550 17926 22602 17978
rect 22614 17926 22666 17978
rect 22678 17926 22730 17978
rect 22742 17926 22794 17978
rect 22806 17926 22858 17978
rect 27350 17926 27402 17978
rect 27414 17926 27466 17978
rect 27478 17926 27530 17978
rect 27542 17926 27594 17978
rect 27606 17926 27658 17978
rect 4436 17824 4488 17876
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 24860 17824 24912 17876
rect 28172 17824 28224 17876
rect 4344 17756 4396 17808
rect 18144 17799 18196 17808
rect 18144 17765 18153 17799
rect 18153 17765 18187 17799
rect 18187 17765 18196 17799
rect 18144 17756 18196 17765
rect 19524 17756 19576 17808
rect 19984 17756 20036 17808
rect 20812 17756 20864 17808
rect 2872 17688 2924 17740
rect 3240 17731 3292 17740
rect 3240 17697 3249 17731
rect 3249 17697 3283 17731
rect 3283 17697 3292 17731
rect 3240 17688 3292 17697
rect 21364 17731 21416 17740
rect 4068 17620 4120 17672
rect 4528 17663 4580 17672
rect 4528 17629 4537 17663
rect 4537 17629 4571 17663
rect 4571 17629 4580 17663
rect 4528 17620 4580 17629
rect 5080 17620 5132 17672
rect 5264 17620 5316 17672
rect 2688 17552 2740 17604
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 4344 17484 4396 17536
rect 5724 17663 5776 17672
rect 5724 17629 5733 17663
rect 5733 17629 5767 17663
rect 5767 17629 5776 17663
rect 21364 17697 21373 17731
rect 21373 17697 21407 17731
rect 21407 17697 21416 17731
rect 21364 17688 21416 17697
rect 26608 17731 26660 17740
rect 26608 17697 26617 17731
rect 26617 17697 26651 17731
rect 26651 17697 26660 17731
rect 26608 17688 26660 17697
rect 5724 17620 5776 17629
rect 6736 17620 6788 17672
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 8024 17663 8076 17672
rect 8024 17629 8033 17663
rect 8033 17629 8067 17663
rect 8067 17629 8076 17663
rect 8024 17620 8076 17629
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 17500 17663 17552 17672
rect 17500 17629 17509 17663
rect 17509 17629 17543 17663
rect 17543 17629 17552 17663
rect 17500 17620 17552 17629
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 20720 17620 20772 17672
rect 20904 17620 20956 17672
rect 7748 17595 7800 17604
rect 6276 17527 6328 17536
rect 6276 17493 6285 17527
rect 6285 17493 6319 17527
rect 6319 17493 6328 17527
rect 6276 17484 6328 17493
rect 7472 17527 7524 17536
rect 7472 17493 7481 17527
rect 7481 17493 7515 17527
rect 7515 17493 7524 17527
rect 7472 17484 7524 17493
rect 7748 17561 7757 17595
rect 7757 17561 7791 17595
rect 7791 17561 7800 17595
rect 7748 17552 7800 17561
rect 8484 17552 8536 17604
rect 9128 17552 9180 17604
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 21548 17620 21600 17672
rect 24492 17663 24544 17672
rect 24492 17629 24501 17663
rect 24501 17629 24535 17663
rect 24535 17629 24544 17663
rect 24492 17620 24544 17629
rect 26332 17663 26384 17672
rect 26332 17629 26341 17663
rect 26341 17629 26375 17663
rect 26375 17629 26384 17663
rect 26332 17620 26384 17629
rect 27712 17620 27764 17672
rect 15844 17484 15896 17536
rect 19800 17484 19852 17536
rect 20536 17484 20588 17536
rect 21456 17552 21508 17604
rect 5750 17382 5802 17434
rect 5814 17382 5866 17434
rect 5878 17382 5930 17434
rect 5942 17382 5994 17434
rect 6006 17382 6058 17434
rect 10550 17382 10602 17434
rect 10614 17382 10666 17434
rect 10678 17382 10730 17434
rect 10742 17382 10794 17434
rect 10806 17382 10858 17434
rect 15350 17382 15402 17434
rect 15414 17382 15466 17434
rect 15478 17382 15530 17434
rect 15542 17382 15594 17434
rect 15606 17382 15658 17434
rect 20150 17382 20202 17434
rect 20214 17382 20266 17434
rect 20278 17382 20330 17434
rect 20342 17382 20394 17434
rect 20406 17382 20458 17434
rect 24950 17382 25002 17434
rect 25014 17382 25066 17434
rect 25078 17382 25130 17434
rect 25142 17382 25194 17434
rect 25206 17382 25258 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 2228 17323 2280 17332
rect 2228 17289 2237 17323
rect 2237 17289 2271 17323
rect 2271 17289 2280 17323
rect 2228 17280 2280 17289
rect 1492 17144 1544 17196
rect 4068 17212 4120 17264
rect 7932 17280 7984 17332
rect 7472 17212 7524 17264
rect 8576 17212 8628 17264
rect 2596 17187 2648 17196
rect 2596 17153 2605 17187
rect 2605 17153 2639 17187
rect 2639 17153 2648 17187
rect 2596 17144 2648 17153
rect 3792 17076 3844 17128
rect 4068 17076 4120 17128
rect 7564 17119 7616 17128
rect 5264 17008 5316 17060
rect 5540 17008 5592 17060
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 10048 17076 10100 17128
rect 15108 17212 15160 17264
rect 17224 17212 17276 17264
rect 17500 17212 17552 17264
rect 20536 17280 20588 17332
rect 18236 17187 18288 17196
rect 14556 17119 14608 17128
rect 14556 17085 14565 17119
rect 14565 17085 14599 17119
rect 14599 17085 14608 17119
rect 14556 17076 14608 17085
rect 15752 17076 15804 17128
rect 16948 17076 17000 17128
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 19800 17187 19852 17196
rect 19800 17153 19809 17187
rect 19809 17153 19843 17187
rect 19843 17153 19852 17187
rect 19800 17144 19852 17153
rect 20076 17212 20128 17264
rect 24768 17280 24820 17332
rect 20168 17144 20220 17196
rect 15200 17008 15252 17060
rect 4528 16940 4580 16992
rect 5632 16940 5684 16992
rect 9312 16983 9364 16992
rect 9312 16949 9321 16983
rect 9321 16949 9355 16983
rect 9355 16949 9364 16983
rect 9312 16940 9364 16949
rect 9772 16940 9824 16992
rect 10876 16940 10928 16992
rect 12348 16940 12400 16992
rect 12808 16940 12860 16992
rect 17592 16940 17644 16992
rect 19340 17008 19392 17060
rect 20720 17144 20772 17196
rect 20812 17144 20864 17196
rect 20996 17144 21048 17196
rect 23296 17144 23348 17196
rect 23112 17076 23164 17128
rect 26056 17212 26108 17264
rect 20628 17051 20680 17060
rect 20628 17017 20637 17051
rect 20637 17017 20671 17051
rect 20671 17017 20680 17051
rect 20628 17008 20680 17017
rect 18788 16983 18840 16992
rect 18788 16949 18797 16983
rect 18797 16949 18831 16983
rect 18831 16949 18840 16983
rect 18788 16940 18840 16949
rect 19984 16940 20036 16992
rect 20168 16940 20220 16992
rect 24952 16940 25004 16992
rect 3350 16838 3402 16890
rect 3414 16838 3466 16890
rect 3478 16838 3530 16890
rect 3542 16838 3594 16890
rect 3606 16838 3658 16890
rect 8150 16838 8202 16890
rect 8214 16838 8266 16890
rect 8278 16838 8330 16890
rect 8342 16838 8394 16890
rect 8406 16838 8458 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 17750 16838 17802 16890
rect 17814 16838 17866 16890
rect 17878 16838 17930 16890
rect 17942 16838 17994 16890
rect 18006 16838 18058 16890
rect 22550 16838 22602 16890
rect 22614 16838 22666 16890
rect 22678 16838 22730 16890
rect 22742 16838 22794 16890
rect 22806 16838 22858 16890
rect 27350 16838 27402 16890
rect 27414 16838 27466 16890
rect 27478 16838 27530 16890
rect 27542 16838 27594 16890
rect 27606 16838 27658 16890
rect 14556 16736 14608 16788
rect 16488 16736 16540 16788
rect 19156 16736 19208 16788
rect 24124 16779 24176 16788
rect 24124 16745 24133 16779
rect 24133 16745 24167 16779
rect 24167 16745 24176 16779
rect 24124 16736 24176 16745
rect 24308 16736 24360 16788
rect 24492 16779 24544 16788
rect 24492 16745 24501 16779
rect 24501 16745 24535 16779
rect 24535 16745 24544 16779
rect 24492 16736 24544 16745
rect 24584 16668 24636 16720
rect 8484 16600 8536 16652
rect 12256 16600 12308 16652
rect 12808 16600 12860 16652
rect 7932 16575 7984 16584
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 8208 16532 8260 16584
rect 9680 16575 9732 16584
rect 7380 16439 7432 16448
rect 7380 16405 7389 16439
rect 7389 16405 7423 16439
rect 7423 16405 7432 16439
rect 7380 16396 7432 16405
rect 8024 16464 8076 16516
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 10416 16532 10468 16584
rect 12072 16532 12124 16584
rect 15108 16600 15160 16652
rect 15844 16600 15896 16652
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 17500 16600 17552 16652
rect 19156 16600 19208 16652
rect 14832 16575 14884 16584
rect 9128 16464 9180 16516
rect 9956 16507 10008 16516
rect 9956 16473 9965 16507
rect 9965 16473 9999 16507
rect 9999 16473 10008 16507
rect 9956 16464 10008 16473
rect 7840 16396 7892 16448
rect 10876 16464 10928 16516
rect 14832 16541 14841 16575
rect 14841 16541 14875 16575
rect 14875 16541 14884 16575
rect 14832 16532 14884 16541
rect 16580 16532 16632 16584
rect 19432 16532 19484 16584
rect 15200 16464 15252 16516
rect 17684 16507 17736 16516
rect 17684 16473 17711 16507
rect 17711 16473 17736 16507
rect 17684 16464 17736 16473
rect 12164 16396 12216 16448
rect 18144 16464 18196 16516
rect 18696 16507 18748 16516
rect 18696 16473 18705 16507
rect 18705 16473 18739 16507
rect 18739 16473 18748 16507
rect 18696 16464 18748 16473
rect 18236 16396 18288 16448
rect 22008 16600 22060 16652
rect 23296 16600 23348 16652
rect 24860 16532 24912 16584
rect 26608 16532 26660 16584
rect 28172 16575 28224 16584
rect 28172 16541 28181 16575
rect 28181 16541 28215 16575
rect 28215 16541 28224 16575
rect 28172 16532 28224 16541
rect 22100 16464 22152 16516
rect 24952 16507 25004 16516
rect 24952 16473 24961 16507
rect 24961 16473 24995 16507
rect 24995 16473 25004 16507
rect 24952 16464 25004 16473
rect 22192 16396 22244 16448
rect 28356 16439 28408 16448
rect 28356 16405 28365 16439
rect 28365 16405 28399 16439
rect 28399 16405 28408 16439
rect 28356 16396 28408 16405
rect 5750 16294 5802 16346
rect 5814 16294 5866 16346
rect 5878 16294 5930 16346
rect 5942 16294 5994 16346
rect 6006 16294 6058 16346
rect 10550 16294 10602 16346
rect 10614 16294 10666 16346
rect 10678 16294 10730 16346
rect 10742 16294 10794 16346
rect 10806 16294 10858 16346
rect 15350 16294 15402 16346
rect 15414 16294 15466 16346
rect 15478 16294 15530 16346
rect 15542 16294 15594 16346
rect 15606 16294 15658 16346
rect 20150 16294 20202 16346
rect 20214 16294 20266 16346
rect 20278 16294 20330 16346
rect 20342 16294 20394 16346
rect 20406 16294 20458 16346
rect 24950 16294 25002 16346
rect 25014 16294 25066 16346
rect 25078 16294 25130 16346
rect 25142 16294 25194 16346
rect 25206 16294 25258 16346
rect 7748 16192 7800 16244
rect 2596 16056 2648 16108
rect 4160 16099 4212 16108
rect 4160 16065 4169 16099
rect 4169 16065 4203 16099
rect 4203 16065 4212 16099
rect 4160 16056 4212 16065
rect 4344 15920 4396 15972
rect 3700 15895 3752 15904
rect 3700 15861 3709 15895
rect 3709 15861 3743 15895
rect 3743 15861 3752 15895
rect 3700 15852 3752 15861
rect 7472 16056 7524 16108
rect 8024 16124 8076 16176
rect 8484 16124 8536 16176
rect 7656 15920 7708 15972
rect 9312 16056 9364 16108
rect 8208 15988 8260 16040
rect 12808 16192 12860 16244
rect 19156 16192 19208 16244
rect 20996 16192 21048 16244
rect 22100 16235 22152 16244
rect 22100 16201 22109 16235
rect 22109 16201 22143 16235
rect 22143 16201 22152 16235
rect 22100 16192 22152 16201
rect 25964 16192 26016 16244
rect 9680 16124 9732 16176
rect 11980 16124 12032 16176
rect 12348 16124 12400 16176
rect 15752 16124 15804 16176
rect 18696 16124 18748 16176
rect 27252 16124 27304 16176
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 14832 16056 14884 16108
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 20536 16056 20588 16108
rect 25504 16056 25556 16108
rect 9956 15988 10008 16040
rect 11060 15988 11112 16040
rect 11612 16031 11664 16040
rect 11612 15997 11621 16031
rect 11621 15997 11655 16031
rect 11655 15997 11664 16031
rect 11612 15988 11664 15997
rect 11888 16031 11940 16040
rect 11888 15997 11897 16031
rect 11897 15997 11931 16031
rect 11931 15997 11940 16031
rect 11888 15988 11940 15997
rect 12348 15988 12400 16040
rect 5172 15852 5224 15904
rect 5264 15895 5316 15904
rect 5264 15861 5273 15895
rect 5273 15861 5307 15895
rect 5307 15861 5316 15895
rect 5264 15852 5316 15861
rect 7840 15852 7892 15904
rect 9128 15895 9180 15904
rect 9128 15861 9137 15895
rect 9137 15861 9171 15895
rect 9171 15861 9180 15895
rect 9128 15852 9180 15861
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 11244 15920 11296 15972
rect 28172 16056 28224 16108
rect 27252 15988 27304 16040
rect 12440 15852 12492 15904
rect 18144 15852 18196 15904
rect 26884 15852 26936 15904
rect 3350 15750 3402 15802
rect 3414 15750 3466 15802
rect 3478 15750 3530 15802
rect 3542 15750 3594 15802
rect 3606 15750 3658 15802
rect 8150 15750 8202 15802
rect 8214 15750 8266 15802
rect 8278 15750 8330 15802
rect 8342 15750 8394 15802
rect 8406 15750 8458 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 17750 15750 17802 15802
rect 17814 15750 17866 15802
rect 17878 15750 17930 15802
rect 17942 15750 17994 15802
rect 18006 15750 18058 15802
rect 22550 15750 22602 15802
rect 22614 15750 22666 15802
rect 22678 15750 22730 15802
rect 22742 15750 22794 15802
rect 22806 15750 22858 15802
rect 27350 15750 27402 15802
rect 27414 15750 27466 15802
rect 27478 15750 27530 15802
rect 27542 15750 27594 15802
rect 27606 15750 27658 15802
rect 2596 15648 2648 15700
rect 3700 15648 3752 15700
rect 4160 15648 4212 15700
rect 5264 15648 5316 15700
rect 8576 15648 8628 15700
rect 10600 15648 10652 15700
rect 11152 15648 11204 15700
rect 11612 15648 11664 15700
rect 3240 15512 3292 15564
rect 19432 15648 19484 15700
rect 20536 15691 20588 15700
rect 20536 15657 20545 15691
rect 20545 15657 20579 15691
rect 20579 15657 20588 15691
rect 20536 15648 20588 15657
rect 28172 15648 28224 15700
rect 19340 15623 19392 15632
rect 19340 15589 19349 15623
rect 19349 15589 19383 15623
rect 19383 15589 19392 15623
rect 19340 15580 19392 15589
rect 20076 15580 20128 15632
rect 24860 15580 24912 15632
rect 15108 15512 15160 15564
rect 2688 15376 2740 15428
rect 11060 15444 11112 15496
rect 19800 15512 19852 15564
rect 21548 15512 21600 15564
rect 26332 15512 26384 15564
rect 26884 15555 26936 15564
rect 26884 15521 26893 15555
rect 26893 15521 26927 15555
rect 26927 15521 26936 15555
rect 26884 15512 26936 15521
rect 21456 15444 21508 15496
rect 9772 15308 9824 15360
rect 12072 15376 12124 15428
rect 15752 15376 15804 15428
rect 20812 15419 20864 15428
rect 20812 15385 20821 15419
rect 20821 15385 20855 15419
rect 20855 15385 20864 15419
rect 20812 15376 20864 15385
rect 15936 15308 15988 15360
rect 21916 15308 21968 15360
rect 24952 15444 25004 15496
rect 26608 15487 26660 15496
rect 26608 15453 26617 15487
rect 26617 15453 26651 15487
rect 26651 15453 26660 15487
rect 26608 15444 26660 15453
rect 27896 15444 27948 15496
rect 25964 15419 26016 15428
rect 25964 15385 25973 15419
rect 25973 15385 26007 15419
rect 26007 15385 26016 15419
rect 25964 15376 26016 15385
rect 25320 15308 25372 15360
rect 5750 15206 5802 15258
rect 5814 15206 5866 15258
rect 5878 15206 5930 15258
rect 5942 15206 5994 15258
rect 6006 15206 6058 15258
rect 10550 15206 10602 15258
rect 10614 15206 10666 15258
rect 10678 15206 10730 15258
rect 10742 15206 10794 15258
rect 10806 15206 10858 15258
rect 15350 15206 15402 15258
rect 15414 15206 15466 15258
rect 15478 15206 15530 15258
rect 15542 15206 15594 15258
rect 15606 15206 15658 15258
rect 20150 15206 20202 15258
rect 20214 15206 20266 15258
rect 20278 15206 20330 15258
rect 20342 15206 20394 15258
rect 20406 15206 20458 15258
rect 24950 15206 25002 15258
rect 25014 15206 25066 15258
rect 25078 15206 25130 15258
rect 25142 15206 25194 15258
rect 25206 15206 25258 15258
rect 7564 15104 7616 15156
rect 11612 15104 11664 15156
rect 3976 15036 4028 15088
rect 5632 15079 5684 15088
rect 5632 15045 5641 15079
rect 5641 15045 5675 15079
rect 5675 15045 5684 15079
rect 5632 15036 5684 15045
rect 7840 15079 7892 15088
rect 7840 15045 7849 15079
rect 7849 15045 7883 15079
rect 7883 15045 7892 15079
rect 7840 15036 7892 15045
rect 8576 15036 8628 15088
rect 11152 15036 11204 15088
rect 12164 15104 12216 15156
rect 17592 15104 17644 15156
rect 12072 15036 12124 15088
rect 3148 15011 3200 15020
rect 3148 14977 3157 15011
rect 3157 14977 3191 15011
rect 3191 14977 3200 15011
rect 3148 14968 3200 14977
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 7564 15011 7616 15020
rect 3884 14900 3936 14952
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 11244 14968 11296 15020
rect 11980 15011 12032 15020
rect 2596 14764 2648 14816
rect 4160 14764 4212 14816
rect 7472 14900 7524 14952
rect 9128 14900 9180 14952
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 19340 15011 19392 15020
rect 19340 14977 19349 15011
rect 19349 14977 19383 15011
rect 19383 14977 19392 15011
rect 19340 14968 19392 14977
rect 20812 15104 20864 15156
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 24860 15104 24912 15156
rect 25504 15147 25556 15156
rect 25504 15113 25513 15147
rect 25513 15113 25547 15147
rect 25547 15113 25556 15147
rect 25504 15104 25556 15113
rect 22284 15079 22336 15088
rect 22284 15045 22293 15079
rect 22293 15045 22327 15079
rect 22327 15045 22336 15079
rect 22284 15036 22336 15045
rect 20720 14968 20772 15020
rect 21272 14968 21324 15020
rect 22192 14968 22244 15020
rect 11888 14832 11940 14884
rect 6552 14764 6604 14816
rect 8484 14764 8536 14816
rect 19156 14943 19208 14952
rect 19156 14909 19165 14943
rect 19165 14909 19199 14943
rect 19199 14909 19208 14943
rect 19156 14900 19208 14909
rect 21916 14900 21968 14952
rect 24216 14968 24268 15020
rect 24124 14900 24176 14952
rect 17224 14832 17276 14884
rect 19708 14832 19760 14884
rect 23112 14832 23164 14884
rect 12348 14764 12400 14816
rect 15752 14764 15804 14816
rect 18420 14764 18472 14816
rect 24400 14807 24452 14816
rect 24400 14773 24409 14807
rect 24409 14773 24443 14807
rect 24443 14773 24452 14807
rect 24400 14764 24452 14773
rect 3350 14662 3402 14714
rect 3414 14662 3466 14714
rect 3478 14662 3530 14714
rect 3542 14662 3594 14714
rect 3606 14662 3658 14714
rect 8150 14662 8202 14714
rect 8214 14662 8266 14714
rect 8278 14662 8330 14714
rect 8342 14662 8394 14714
rect 8406 14662 8458 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 17750 14662 17802 14714
rect 17814 14662 17866 14714
rect 17878 14662 17930 14714
rect 17942 14662 17994 14714
rect 18006 14662 18058 14714
rect 22550 14662 22602 14714
rect 22614 14662 22666 14714
rect 22678 14662 22730 14714
rect 22742 14662 22794 14714
rect 22806 14662 22858 14714
rect 27350 14662 27402 14714
rect 27414 14662 27466 14714
rect 27478 14662 27530 14714
rect 27542 14662 27594 14714
rect 27606 14662 27658 14714
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 19432 14560 19484 14612
rect 21548 14603 21600 14612
rect 21548 14569 21557 14603
rect 21557 14569 21591 14603
rect 21591 14569 21600 14603
rect 21548 14560 21600 14569
rect 4344 14492 4396 14544
rect 21272 14492 21324 14544
rect 21916 14492 21968 14544
rect 4160 14399 4212 14408
rect 4160 14365 4183 14399
rect 4183 14365 4212 14399
rect 4160 14356 4212 14365
rect 8484 14424 8536 14476
rect 12256 14424 12308 14476
rect 16212 14424 16264 14476
rect 5172 14399 5224 14408
rect 5172 14365 5181 14399
rect 5181 14365 5215 14399
rect 5215 14365 5224 14399
rect 5172 14356 5224 14365
rect 6276 14356 6328 14408
rect 5264 14288 5316 14340
rect 5816 14288 5868 14340
rect 6644 14331 6696 14340
rect 6644 14297 6653 14331
rect 6653 14297 6687 14331
rect 6687 14297 6696 14331
rect 6644 14288 6696 14297
rect 7104 14288 7156 14340
rect 15108 14288 15160 14340
rect 16580 14288 16632 14340
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17500 14356 17552 14408
rect 22284 14424 22336 14476
rect 22192 14356 22244 14408
rect 16948 14331 17000 14340
rect 16948 14297 16957 14331
rect 16957 14297 16991 14331
rect 16991 14297 17000 14331
rect 16948 14288 17000 14297
rect 22100 14331 22152 14340
rect 4804 14263 4856 14272
rect 4804 14229 4813 14263
rect 4813 14229 4847 14263
rect 4847 14229 4856 14263
rect 4804 14220 4856 14229
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 16672 14220 16724 14272
rect 22100 14297 22109 14331
rect 22109 14297 22143 14331
rect 22143 14297 22152 14331
rect 22100 14288 22152 14297
rect 21824 14220 21876 14272
rect 5750 14118 5802 14170
rect 5814 14118 5866 14170
rect 5878 14118 5930 14170
rect 5942 14118 5994 14170
rect 6006 14118 6058 14170
rect 10550 14118 10602 14170
rect 10614 14118 10666 14170
rect 10678 14118 10730 14170
rect 10742 14118 10794 14170
rect 10806 14118 10858 14170
rect 15350 14118 15402 14170
rect 15414 14118 15466 14170
rect 15478 14118 15530 14170
rect 15542 14118 15594 14170
rect 15606 14118 15658 14170
rect 20150 14118 20202 14170
rect 20214 14118 20266 14170
rect 20278 14118 20330 14170
rect 20342 14118 20394 14170
rect 20406 14118 20458 14170
rect 24950 14118 25002 14170
rect 25014 14118 25066 14170
rect 25078 14118 25130 14170
rect 25142 14118 25194 14170
rect 25206 14118 25258 14170
rect 6552 13991 6604 14000
rect 6552 13957 6561 13991
rect 6561 13957 6595 13991
rect 6595 13957 6604 13991
rect 6552 13948 6604 13957
rect 15752 14016 15804 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 24216 14059 24268 14068
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 16672 13948 16724 14000
rect 18420 13991 18472 14000
rect 18420 13957 18429 13991
rect 18429 13957 18463 13991
rect 18463 13957 18472 13991
rect 18420 13948 18472 13957
rect 24216 14025 24225 14059
rect 24225 14025 24259 14059
rect 24259 14025 24268 14059
rect 24216 14016 24268 14025
rect 25320 13948 25372 14000
rect 15384 13880 15436 13889
rect 12440 13812 12492 13864
rect 6736 13787 6788 13796
rect 6736 13753 6745 13787
rect 6745 13753 6779 13787
rect 6779 13753 6788 13787
rect 6736 13744 6788 13753
rect 14188 13744 14240 13796
rect 15752 13812 15804 13864
rect 15108 13787 15160 13796
rect 15108 13753 15117 13787
rect 15117 13753 15151 13787
rect 15151 13753 15160 13787
rect 15108 13744 15160 13753
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 16212 13812 16264 13864
rect 20720 13880 20772 13932
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 22284 13880 22336 13932
rect 27252 13923 27304 13932
rect 12532 13719 12584 13728
rect 12532 13685 12541 13719
rect 12541 13685 12575 13719
rect 12575 13685 12584 13719
rect 12532 13676 12584 13685
rect 14832 13676 14884 13728
rect 20996 13812 21048 13864
rect 22008 13812 22060 13864
rect 27252 13889 27261 13923
rect 27261 13889 27295 13923
rect 27295 13889 27304 13923
rect 27252 13880 27304 13889
rect 28172 13923 28224 13932
rect 28172 13889 28181 13923
rect 28181 13889 28215 13923
rect 28215 13889 28224 13923
rect 28172 13880 28224 13889
rect 21180 13676 21232 13728
rect 21916 13676 21968 13728
rect 26884 13676 26936 13728
rect 28356 13719 28408 13728
rect 28356 13685 28365 13719
rect 28365 13685 28399 13719
rect 28399 13685 28408 13719
rect 28356 13676 28408 13685
rect 3350 13574 3402 13626
rect 3414 13574 3466 13626
rect 3478 13574 3530 13626
rect 3542 13574 3594 13626
rect 3606 13574 3658 13626
rect 8150 13574 8202 13626
rect 8214 13574 8266 13626
rect 8278 13574 8330 13626
rect 8342 13574 8394 13626
rect 8406 13574 8458 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 17750 13574 17802 13626
rect 17814 13574 17866 13626
rect 17878 13574 17930 13626
rect 17942 13574 17994 13626
rect 18006 13574 18058 13626
rect 22550 13574 22602 13626
rect 22614 13574 22666 13626
rect 22678 13574 22730 13626
rect 22742 13574 22794 13626
rect 22806 13574 22858 13626
rect 27350 13574 27402 13626
rect 27414 13574 27466 13626
rect 27478 13574 27530 13626
rect 27542 13574 27594 13626
rect 27606 13574 27658 13626
rect 2412 13311 2464 13320
rect 2412 13277 2421 13311
rect 2421 13277 2455 13311
rect 2455 13277 2464 13311
rect 2412 13268 2464 13277
rect 4988 13268 5040 13320
rect 9772 13472 9824 13524
rect 10968 13472 11020 13524
rect 13544 13472 13596 13524
rect 14096 13472 14148 13524
rect 14832 13515 14884 13524
rect 14832 13481 14841 13515
rect 14841 13481 14875 13515
rect 14875 13481 14884 13515
rect 15384 13515 15436 13524
rect 14832 13472 14884 13481
rect 15384 13481 15393 13515
rect 15393 13481 15427 13515
rect 15427 13481 15436 13515
rect 15384 13472 15436 13481
rect 20536 13515 20588 13524
rect 20536 13481 20545 13515
rect 20545 13481 20579 13515
rect 20579 13481 20588 13515
rect 20536 13472 20588 13481
rect 20812 13472 20864 13524
rect 22008 13472 22060 13524
rect 12532 13404 12584 13456
rect 8576 13336 8628 13388
rect 9036 13311 9088 13320
rect 9036 13277 9045 13311
rect 9045 13277 9079 13311
rect 9079 13277 9088 13311
rect 9036 13268 9088 13277
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 2964 13200 3016 13252
rect 3976 13200 4028 13252
rect 1768 13132 1820 13184
rect 5080 13175 5132 13184
rect 5080 13141 5089 13175
rect 5089 13141 5123 13175
rect 5123 13141 5132 13175
rect 5080 13132 5132 13141
rect 9588 13200 9640 13252
rect 9772 13200 9824 13252
rect 11152 13132 11204 13184
rect 12256 13132 12308 13184
rect 12808 13132 12860 13184
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 15200 13336 15252 13388
rect 17592 13404 17644 13456
rect 16948 13336 17000 13388
rect 17316 13336 17368 13388
rect 26884 13379 26936 13388
rect 26884 13345 26893 13379
rect 26893 13345 26927 13379
rect 26927 13345 26936 13379
rect 26884 13336 26936 13345
rect 16672 13311 16724 13320
rect 15844 13200 15896 13252
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 17224 13268 17276 13320
rect 20812 13311 20864 13320
rect 20812 13277 20821 13311
rect 20821 13277 20855 13311
rect 20855 13277 20864 13311
rect 20812 13268 20864 13277
rect 21916 13268 21968 13320
rect 25412 13268 25464 13320
rect 26608 13311 26660 13320
rect 26608 13277 26617 13311
rect 26617 13277 26651 13311
rect 26651 13277 26660 13311
rect 26608 13268 26660 13277
rect 16764 13200 16816 13252
rect 17040 13200 17092 13252
rect 25320 13200 25372 13252
rect 15200 13132 15252 13184
rect 16580 13132 16632 13184
rect 16948 13175 17000 13184
rect 16948 13141 16957 13175
rect 16957 13141 16991 13175
rect 16991 13141 17000 13175
rect 23020 13175 23072 13184
rect 16948 13132 17000 13141
rect 23020 13141 23029 13175
rect 23029 13141 23063 13175
rect 23063 13141 23072 13175
rect 23020 13132 23072 13141
rect 25872 13132 25924 13184
rect 27712 13132 27764 13184
rect 28172 13132 28224 13184
rect 5750 13030 5802 13082
rect 5814 13030 5866 13082
rect 5878 13030 5930 13082
rect 5942 13030 5994 13082
rect 6006 13030 6058 13082
rect 10550 13030 10602 13082
rect 10614 13030 10666 13082
rect 10678 13030 10730 13082
rect 10742 13030 10794 13082
rect 10806 13030 10858 13082
rect 15350 13030 15402 13082
rect 15414 13030 15466 13082
rect 15478 13030 15530 13082
rect 15542 13030 15594 13082
rect 15606 13030 15658 13082
rect 20150 13030 20202 13082
rect 20214 13030 20266 13082
rect 20278 13030 20330 13082
rect 20342 13030 20394 13082
rect 20406 13030 20458 13082
rect 24950 13030 25002 13082
rect 25014 13030 25066 13082
rect 25078 13030 25130 13082
rect 25142 13030 25194 13082
rect 25206 13030 25258 13082
rect 1768 12903 1820 12912
rect 1768 12869 1777 12903
rect 1777 12869 1811 12903
rect 1811 12869 1820 12903
rect 1768 12860 1820 12869
rect 3148 12860 3200 12912
rect 3976 12860 4028 12912
rect 4804 12860 4856 12912
rect 6644 12860 6696 12912
rect 8484 12928 8536 12980
rect 9588 12971 9640 12980
rect 9588 12937 9597 12971
rect 9597 12937 9631 12971
rect 9631 12937 9640 12971
rect 9588 12928 9640 12937
rect 11244 12928 11296 12980
rect 11336 12928 11388 12980
rect 12440 12928 12492 12980
rect 16764 12971 16816 12980
rect 16764 12937 16773 12971
rect 16773 12937 16807 12971
rect 16807 12937 16816 12971
rect 16764 12928 16816 12937
rect 23020 12928 23072 12980
rect 27252 12971 27304 12980
rect 27252 12937 27261 12971
rect 27261 12937 27295 12971
rect 27295 12937 27304 12971
rect 27252 12928 27304 12937
rect 27712 12971 27764 12980
rect 27712 12937 27721 12971
rect 27721 12937 27755 12971
rect 27755 12937 27764 12971
rect 27712 12928 27764 12937
rect 1768 12724 1820 12776
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 3976 12588 4028 12640
rect 5080 12792 5132 12844
rect 12532 12860 12584 12912
rect 20996 12860 21048 12912
rect 21824 12860 21876 12912
rect 8576 12792 8628 12844
rect 9680 12835 9732 12844
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6736 12724 6788 12733
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 10968 12835 11020 12844
rect 9864 12724 9916 12776
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 12256 12835 12308 12844
rect 12256 12801 12265 12835
rect 12265 12801 12299 12835
rect 12299 12801 12308 12835
rect 12256 12792 12308 12801
rect 13820 12792 13872 12844
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 21456 12835 21508 12844
rect 15936 12767 15988 12776
rect 4344 12656 4396 12708
rect 15936 12733 15945 12767
rect 15945 12733 15979 12767
rect 15979 12733 15988 12767
rect 15936 12724 15988 12733
rect 16488 12724 16540 12776
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 22284 12903 22336 12912
rect 22284 12869 22293 12903
rect 22293 12869 22327 12903
rect 22327 12869 22336 12903
rect 22284 12860 22336 12869
rect 25320 12860 25372 12912
rect 25872 12903 25924 12912
rect 25872 12869 25881 12903
rect 25881 12869 25915 12903
rect 25915 12869 25924 12903
rect 25872 12860 25924 12869
rect 21456 12792 21508 12801
rect 26608 12792 26660 12844
rect 22100 12724 22152 12776
rect 22284 12724 22336 12776
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 6368 12588 6420 12640
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 8668 12631 8720 12640
rect 8668 12597 8677 12631
rect 8677 12597 8711 12631
rect 8711 12597 8720 12631
rect 8668 12588 8720 12597
rect 9680 12588 9732 12640
rect 11336 12656 11388 12708
rect 10416 12588 10468 12640
rect 12348 12631 12400 12640
rect 12348 12597 12357 12631
rect 12357 12597 12391 12631
rect 12391 12597 12400 12631
rect 12348 12588 12400 12597
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 16948 12631 17000 12640
rect 16948 12597 16957 12631
rect 16957 12597 16991 12631
rect 16991 12597 17000 12631
rect 16948 12588 17000 12597
rect 21916 12699 21968 12708
rect 21916 12665 21925 12699
rect 21925 12665 21959 12699
rect 21959 12665 21968 12699
rect 21916 12656 21968 12665
rect 20812 12588 20864 12640
rect 21824 12588 21876 12640
rect 24860 12588 24912 12640
rect 26700 12631 26752 12640
rect 26700 12597 26709 12631
rect 26709 12597 26743 12631
rect 26743 12597 26752 12631
rect 26700 12588 26752 12597
rect 3350 12486 3402 12538
rect 3414 12486 3466 12538
rect 3478 12486 3530 12538
rect 3542 12486 3594 12538
rect 3606 12486 3658 12538
rect 8150 12486 8202 12538
rect 8214 12486 8266 12538
rect 8278 12486 8330 12538
rect 8342 12486 8394 12538
rect 8406 12486 8458 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 17750 12486 17802 12538
rect 17814 12486 17866 12538
rect 17878 12486 17930 12538
rect 17942 12486 17994 12538
rect 18006 12486 18058 12538
rect 22550 12486 22602 12538
rect 22614 12486 22666 12538
rect 22678 12486 22730 12538
rect 22742 12486 22794 12538
rect 22806 12486 22858 12538
rect 27350 12486 27402 12538
rect 27414 12486 27466 12538
rect 27478 12486 27530 12538
rect 27542 12486 27594 12538
rect 27606 12486 27658 12538
rect 1492 12384 1544 12436
rect 2412 12384 2464 12436
rect 15200 12384 15252 12436
rect 25412 12427 25464 12436
rect 6736 12316 6788 12368
rect 12348 12359 12400 12368
rect 12348 12325 12357 12359
rect 12357 12325 12391 12359
rect 12391 12325 12400 12359
rect 12348 12316 12400 12325
rect 3884 12248 3936 12300
rect 7380 12248 7432 12300
rect 9588 12248 9640 12300
rect 3240 12180 3292 12232
rect 6368 12223 6420 12232
rect 2596 12155 2648 12164
rect 2596 12121 2605 12155
rect 2605 12121 2639 12155
rect 2639 12121 2648 12155
rect 2596 12112 2648 12121
rect 3148 12044 3200 12096
rect 3700 12044 3752 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 12256 12180 12308 12232
rect 25412 12393 25421 12427
rect 25421 12393 25455 12427
rect 25455 12393 25464 12427
rect 25412 12384 25464 12393
rect 17040 12316 17092 12368
rect 16948 12248 17000 12300
rect 19984 12291 20036 12300
rect 19984 12257 19993 12291
rect 19993 12257 20027 12291
rect 20027 12257 20036 12291
rect 19984 12248 20036 12257
rect 12900 12180 12952 12232
rect 9864 12155 9916 12164
rect 9864 12121 9873 12155
rect 9873 12121 9907 12155
rect 9907 12121 9916 12155
rect 9864 12112 9916 12121
rect 10968 12112 11020 12164
rect 16764 12180 16816 12232
rect 17040 12180 17092 12232
rect 17316 12180 17368 12232
rect 24216 12248 24268 12300
rect 24400 12248 24452 12300
rect 24860 12248 24912 12300
rect 22284 12180 22336 12232
rect 6828 12044 6880 12096
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 10140 12044 10192 12096
rect 12808 12044 12860 12096
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 17500 12044 17552 12096
rect 17776 12044 17828 12096
rect 23388 12112 23440 12164
rect 20628 12044 20680 12096
rect 24216 12044 24268 12096
rect 5750 11942 5802 11994
rect 5814 11942 5866 11994
rect 5878 11942 5930 11994
rect 5942 11942 5994 11994
rect 6006 11942 6058 11994
rect 10550 11942 10602 11994
rect 10614 11942 10666 11994
rect 10678 11942 10730 11994
rect 10742 11942 10794 11994
rect 10806 11942 10858 11994
rect 15350 11942 15402 11994
rect 15414 11942 15466 11994
rect 15478 11942 15530 11994
rect 15542 11942 15594 11994
rect 15606 11942 15658 11994
rect 20150 11942 20202 11994
rect 20214 11942 20266 11994
rect 20278 11942 20330 11994
rect 20342 11942 20394 11994
rect 20406 11942 20458 11994
rect 24950 11942 25002 11994
rect 25014 11942 25066 11994
rect 25078 11942 25130 11994
rect 25142 11942 25194 11994
rect 25206 11942 25258 11994
rect 4988 11840 5040 11892
rect 16672 11840 16724 11892
rect 17132 11840 17184 11892
rect 20628 11840 20680 11892
rect 3700 11772 3752 11824
rect 3976 11815 4028 11824
rect 3976 11781 3985 11815
rect 3985 11781 4019 11815
rect 4019 11781 4028 11815
rect 3976 11772 4028 11781
rect 13544 11772 13596 11824
rect 18236 11772 18288 11824
rect 6368 11704 6420 11756
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 17776 11747 17828 11756
rect 17776 11713 17785 11747
rect 17785 11713 17819 11747
rect 17819 11713 17828 11747
rect 17776 11704 17828 11713
rect 20812 11704 20864 11756
rect 23940 11704 23992 11756
rect 27160 11704 27212 11756
rect 28172 11747 28224 11756
rect 28172 11713 28181 11747
rect 28181 11713 28215 11747
rect 28215 11713 28224 11747
rect 28172 11704 28224 11713
rect 1768 11636 1820 11688
rect 4804 11636 4856 11688
rect 8760 11636 8812 11688
rect 9036 11568 9088 11620
rect 2964 11500 3016 11552
rect 7564 11500 7616 11552
rect 13360 11500 13412 11552
rect 13912 11543 13964 11552
rect 13912 11509 13921 11543
rect 13921 11509 13955 11543
rect 13955 11509 13964 11543
rect 13912 11500 13964 11509
rect 19248 11568 19300 11620
rect 18144 11500 18196 11552
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 26700 11636 26752 11688
rect 18420 11500 18472 11509
rect 23848 11500 23900 11552
rect 26792 11500 26844 11552
rect 28356 11543 28408 11552
rect 28356 11509 28365 11543
rect 28365 11509 28399 11543
rect 28399 11509 28408 11543
rect 28356 11500 28408 11509
rect 3350 11398 3402 11450
rect 3414 11398 3466 11450
rect 3478 11398 3530 11450
rect 3542 11398 3594 11450
rect 3606 11398 3658 11450
rect 8150 11398 8202 11450
rect 8214 11398 8266 11450
rect 8278 11398 8330 11450
rect 8342 11398 8394 11450
rect 8406 11398 8458 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 17750 11398 17802 11450
rect 17814 11398 17866 11450
rect 17878 11398 17930 11450
rect 17942 11398 17994 11450
rect 18006 11398 18058 11450
rect 22550 11398 22602 11450
rect 22614 11398 22666 11450
rect 22678 11398 22730 11450
rect 22742 11398 22794 11450
rect 22806 11398 22858 11450
rect 27350 11398 27402 11450
rect 27414 11398 27466 11450
rect 27478 11398 27530 11450
rect 27542 11398 27594 11450
rect 27606 11398 27658 11450
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 4528 10956 4580 11008
rect 7012 11092 7064 11144
rect 10968 11296 11020 11348
rect 12808 11296 12860 11348
rect 9588 11203 9640 11212
rect 9588 11169 9597 11203
rect 9597 11169 9631 11203
rect 9631 11169 9640 11203
rect 9588 11160 9640 11169
rect 11060 11160 11112 11212
rect 13360 11203 13412 11212
rect 13360 11169 13369 11203
rect 13369 11169 13403 11203
rect 13403 11169 13412 11203
rect 13360 11160 13412 11169
rect 8668 11092 8720 11144
rect 16304 11160 16356 11212
rect 16764 11092 16816 11144
rect 23480 11160 23532 11212
rect 26792 11203 26844 11212
rect 26792 11169 26801 11203
rect 26801 11169 26835 11203
rect 26835 11169 26844 11203
rect 26792 11160 26844 11169
rect 17316 11092 17368 11144
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 10416 10956 10468 11008
rect 15752 10956 15804 11008
rect 16672 10956 16724 11008
rect 16764 10956 16816 11008
rect 16948 10956 17000 11008
rect 17592 10956 17644 11008
rect 18236 11024 18288 11076
rect 23388 11024 23440 11076
rect 23848 11067 23900 11076
rect 23848 11033 23857 11067
rect 23857 11033 23891 11067
rect 23891 11033 23900 11067
rect 23848 11024 23900 11033
rect 27804 11024 27856 11076
rect 27620 10956 27672 11008
rect 27712 10956 27764 11008
rect 28172 10956 28224 11008
rect 5750 10854 5802 10906
rect 5814 10854 5866 10906
rect 5878 10854 5930 10906
rect 5942 10854 5994 10906
rect 6006 10854 6058 10906
rect 10550 10854 10602 10906
rect 10614 10854 10666 10906
rect 10678 10854 10730 10906
rect 10742 10854 10794 10906
rect 10806 10854 10858 10906
rect 15350 10854 15402 10906
rect 15414 10854 15466 10906
rect 15478 10854 15530 10906
rect 15542 10854 15594 10906
rect 15606 10854 15658 10906
rect 20150 10854 20202 10906
rect 20214 10854 20266 10906
rect 20278 10854 20330 10906
rect 20342 10854 20394 10906
rect 20406 10854 20458 10906
rect 24950 10854 25002 10906
rect 25014 10854 25066 10906
rect 25078 10854 25130 10906
rect 25142 10854 25194 10906
rect 25206 10854 25258 10906
rect 4528 10752 4580 10804
rect 9036 10752 9088 10804
rect 12808 10752 12860 10804
rect 9496 10684 9548 10736
rect 10968 10684 11020 10736
rect 4620 10659 4672 10668
rect 4620 10625 4629 10659
rect 4629 10625 4663 10659
rect 4663 10625 4672 10659
rect 4620 10616 4672 10625
rect 4252 10591 4304 10600
rect 4252 10557 4261 10591
rect 4261 10557 4295 10591
rect 4295 10557 4304 10591
rect 4252 10548 4304 10557
rect 4988 10548 5040 10600
rect 5540 10616 5592 10668
rect 10324 10616 10376 10668
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 11060 10659 11112 10668
rect 10416 10616 10468 10625
rect 11060 10625 11069 10659
rect 11069 10625 11103 10659
rect 11103 10625 11112 10659
rect 11060 10616 11112 10625
rect 11980 10616 12032 10668
rect 16212 10752 16264 10804
rect 19984 10752 20036 10804
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 23940 10795 23992 10804
rect 23940 10761 23949 10795
rect 23949 10761 23983 10795
rect 23983 10761 23992 10795
rect 23940 10752 23992 10761
rect 27160 10752 27212 10804
rect 27620 10795 27672 10804
rect 27620 10761 27629 10795
rect 27629 10761 27663 10795
rect 27663 10761 27672 10795
rect 27620 10752 27672 10761
rect 27712 10795 27764 10804
rect 27712 10761 27721 10795
rect 27721 10761 27755 10795
rect 27755 10761 27764 10795
rect 27712 10752 27764 10761
rect 19248 10727 19300 10736
rect 19248 10693 19257 10727
rect 19257 10693 19291 10727
rect 19291 10693 19300 10727
rect 19248 10684 19300 10693
rect 9956 10548 10008 10600
rect 15752 10616 15804 10668
rect 16304 10659 16356 10668
rect 16304 10625 16313 10659
rect 16313 10625 16347 10659
rect 16347 10625 16356 10659
rect 16304 10616 16356 10625
rect 18144 10616 18196 10668
rect 16672 10548 16724 10600
rect 20076 10548 20128 10600
rect 12624 10480 12676 10532
rect 16948 10480 17000 10532
rect 21824 10616 21876 10668
rect 20996 10591 21048 10600
rect 20996 10557 21005 10591
rect 21005 10557 21039 10591
rect 21039 10557 21048 10591
rect 20996 10548 21048 10557
rect 20904 10480 20956 10532
rect 21456 10548 21508 10600
rect 24216 10548 24268 10600
rect 10140 10412 10192 10464
rect 15936 10455 15988 10464
rect 15936 10421 15945 10455
rect 15945 10421 15979 10455
rect 15979 10421 15988 10455
rect 15936 10412 15988 10421
rect 16764 10412 16816 10464
rect 20352 10412 20404 10464
rect 26700 10455 26752 10464
rect 26700 10421 26709 10455
rect 26709 10421 26743 10455
rect 26743 10421 26752 10455
rect 26700 10412 26752 10421
rect 3350 10310 3402 10362
rect 3414 10310 3466 10362
rect 3478 10310 3530 10362
rect 3542 10310 3594 10362
rect 3606 10310 3658 10362
rect 8150 10310 8202 10362
rect 8214 10310 8266 10362
rect 8278 10310 8330 10362
rect 8342 10310 8394 10362
rect 8406 10310 8458 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 17750 10310 17802 10362
rect 17814 10310 17866 10362
rect 17878 10310 17930 10362
rect 17942 10310 17994 10362
rect 18006 10310 18058 10362
rect 22550 10310 22602 10362
rect 22614 10310 22666 10362
rect 22678 10310 22730 10362
rect 22742 10310 22794 10362
rect 22806 10310 22858 10362
rect 27350 10310 27402 10362
rect 27414 10310 27466 10362
rect 27478 10310 27530 10362
rect 27542 10310 27594 10362
rect 27606 10310 27658 10362
rect 12716 10208 12768 10260
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 13728 10208 13780 10260
rect 13912 10208 13964 10260
rect 21824 10251 21876 10260
rect 21824 10217 21833 10251
rect 21833 10217 21867 10251
rect 21867 10217 21876 10251
rect 21824 10208 21876 10217
rect 4620 10183 4672 10192
rect 4620 10149 4629 10183
rect 4629 10149 4663 10183
rect 4663 10149 4672 10183
rect 4620 10140 4672 10149
rect 4988 10072 5040 10124
rect 6736 10140 6788 10192
rect 9772 10140 9824 10192
rect 10416 10140 10468 10192
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 5540 10004 5592 10056
rect 16120 10072 16172 10124
rect 17592 10072 17644 10124
rect 20352 10115 20404 10124
rect 20352 10081 20361 10115
rect 20361 10081 20395 10115
rect 20395 10081 20404 10115
rect 20352 10072 20404 10081
rect 4988 9936 5040 9988
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 6920 9936 6972 9988
rect 4528 9868 4580 9920
rect 9956 10004 10008 10056
rect 10324 10004 10376 10056
rect 12624 10004 12676 10056
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 13084 9936 13136 9988
rect 13728 10004 13780 10056
rect 18144 10004 18196 10056
rect 19432 10004 19484 10056
rect 20076 10047 20128 10056
rect 20076 10013 20085 10047
rect 20085 10013 20119 10047
rect 20119 10013 20128 10047
rect 20076 10004 20128 10013
rect 15936 9936 15988 9988
rect 8300 9868 8352 9920
rect 9680 9868 9732 9920
rect 10140 9911 10192 9920
rect 10140 9877 10149 9911
rect 10149 9877 10183 9911
rect 10183 9877 10192 9911
rect 10140 9868 10192 9877
rect 16764 9868 16816 9920
rect 23388 9936 23440 9988
rect 5750 9766 5802 9818
rect 5814 9766 5866 9818
rect 5878 9766 5930 9818
rect 5942 9766 5994 9818
rect 6006 9766 6058 9818
rect 10550 9766 10602 9818
rect 10614 9766 10666 9818
rect 10678 9766 10730 9818
rect 10742 9766 10794 9818
rect 10806 9766 10858 9818
rect 15350 9766 15402 9818
rect 15414 9766 15466 9818
rect 15478 9766 15530 9818
rect 15542 9766 15594 9818
rect 15606 9766 15658 9818
rect 20150 9766 20202 9818
rect 20214 9766 20266 9818
rect 20278 9766 20330 9818
rect 20342 9766 20394 9818
rect 20406 9766 20458 9818
rect 24950 9766 25002 9818
rect 25014 9766 25066 9818
rect 25078 9766 25130 9818
rect 25142 9766 25194 9818
rect 25206 9766 25258 9818
rect 4528 9664 4580 9716
rect 9680 9664 9732 9716
rect 10324 9664 10376 9716
rect 6920 9596 6972 9648
rect 11980 9639 12032 9648
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 8484 9571 8536 9580
rect 8484 9537 8493 9571
rect 8493 9537 8527 9571
rect 8527 9537 8536 9571
rect 8484 9528 8536 9537
rect 9588 9528 9640 9580
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 9956 9528 10008 9580
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 12716 9664 12768 9716
rect 11060 9528 11112 9580
rect 15936 9596 15988 9648
rect 16580 9528 16632 9580
rect 16948 9571 17000 9580
rect 16948 9537 16957 9571
rect 16957 9537 16991 9571
rect 16991 9537 17000 9571
rect 16948 9528 17000 9537
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 18512 9528 18564 9580
rect 24860 9528 24912 9580
rect 27160 9528 27212 9580
rect 28264 9528 28316 9580
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 4988 9460 5040 9512
rect 9496 9503 9548 9512
rect 8576 9392 8628 9444
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 9128 9435 9180 9444
rect 9128 9401 9137 9435
rect 9137 9401 9171 9435
rect 9171 9401 9180 9435
rect 9128 9392 9180 9401
rect 8760 9324 8812 9376
rect 12256 9460 12308 9512
rect 12716 9460 12768 9512
rect 13084 9460 13136 9512
rect 16764 9503 16816 9512
rect 16764 9469 16773 9503
rect 16773 9469 16807 9503
rect 16807 9469 16816 9503
rect 16764 9460 16816 9469
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 9680 9324 9732 9376
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 25964 9324 26016 9376
rect 26792 9324 26844 9376
rect 28356 9367 28408 9376
rect 28356 9333 28365 9367
rect 28365 9333 28399 9367
rect 28399 9333 28408 9367
rect 28356 9324 28408 9333
rect 3350 9222 3402 9274
rect 3414 9222 3466 9274
rect 3478 9222 3530 9274
rect 3542 9222 3594 9274
rect 3606 9222 3658 9274
rect 8150 9222 8202 9274
rect 8214 9222 8266 9274
rect 8278 9222 8330 9274
rect 8342 9222 8394 9274
rect 8406 9222 8458 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 17750 9222 17802 9274
rect 17814 9222 17866 9274
rect 17878 9222 17930 9274
rect 17942 9222 17994 9274
rect 18006 9222 18058 9274
rect 22550 9222 22602 9274
rect 22614 9222 22666 9274
rect 22678 9222 22730 9274
rect 22742 9222 22794 9274
rect 22806 9222 22858 9274
rect 27350 9222 27402 9274
rect 27414 9222 27466 9274
rect 27478 9222 27530 9274
rect 27542 9222 27594 9274
rect 27606 9222 27658 9274
rect 12256 9163 12308 9172
rect 12256 9129 12265 9163
rect 12265 9129 12299 9163
rect 12299 9129 12308 9163
rect 12256 9120 12308 9129
rect 12716 9163 12768 9172
rect 12716 9129 12725 9163
rect 12725 9129 12759 9163
rect 12759 9129 12768 9163
rect 12716 9120 12768 9129
rect 13084 9120 13136 9172
rect 4620 9095 4672 9104
rect 4620 9061 4629 9095
rect 4629 9061 4663 9095
rect 4663 9061 4672 9095
rect 4620 9052 4672 9061
rect 4252 9027 4304 9036
rect 4252 8993 4261 9027
rect 4261 8993 4295 9027
rect 4295 8993 4304 9027
rect 4252 8984 4304 8993
rect 9128 8984 9180 9036
rect 25964 9027 26016 9036
rect 25964 8993 25973 9027
rect 25973 8993 26007 9027
rect 26007 8993 26016 9027
rect 25964 8984 26016 8993
rect 26792 9027 26844 9036
rect 26792 8993 26801 9027
rect 26801 8993 26835 9027
rect 26835 8993 26844 9027
rect 26792 8984 26844 8993
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 8484 8916 8536 8968
rect 10876 8916 10928 8968
rect 8116 8891 8168 8900
rect 8116 8857 8125 8891
rect 8125 8857 8159 8891
rect 8159 8857 8168 8891
rect 8116 8848 8168 8857
rect 12716 8848 12768 8900
rect 19340 8916 19392 8968
rect 20076 8916 20128 8968
rect 23388 8916 23440 8968
rect 26516 8959 26568 8968
rect 26516 8925 26525 8959
rect 26525 8925 26559 8959
rect 26559 8925 26568 8959
rect 26516 8916 26568 8925
rect 21824 8891 21876 8900
rect 21824 8857 21833 8891
rect 21833 8857 21867 8891
rect 21867 8857 21876 8891
rect 21824 8848 21876 8857
rect 23940 8848 23992 8900
rect 27804 8848 27856 8900
rect 4528 8780 4580 8832
rect 5448 8780 5500 8832
rect 23296 8823 23348 8832
rect 23296 8789 23305 8823
rect 23305 8789 23339 8823
rect 23339 8789 23348 8823
rect 23296 8780 23348 8789
rect 24492 8823 24544 8832
rect 24492 8789 24501 8823
rect 24501 8789 24535 8823
rect 24535 8789 24544 8823
rect 24492 8780 24544 8789
rect 25964 8780 26016 8832
rect 27620 8780 27672 8832
rect 28264 8823 28316 8832
rect 28264 8789 28273 8823
rect 28273 8789 28307 8823
rect 28307 8789 28316 8823
rect 28264 8780 28316 8789
rect 5750 8678 5802 8730
rect 5814 8678 5866 8730
rect 5878 8678 5930 8730
rect 5942 8678 5994 8730
rect 6006 8678 6058 8730
rect 10550 8678 10602 8730
rect 10614 8678 10666 8730
rect 10678 8678 10730 8730
rect 10742 8678 10794 8730
rect 10806 8678 10858 8730
rect 15350 8678 15402 8730
rect 15414 8678 15466 8730
rect 15478 8678 15530 8730
rect 15542 8678 15594 8730
rect 15606 8678 15658 8730
rect 20150 8678 20202 8730
rect 20214 8678 20266 8730
rect 20278 8678 20330 8730
rect 20342 8678 20394 8730
rect 20406 8678 20458 8730
rect 24950 8678 25002 8730
rect 25014 8678 25066 8730
rect 25078 8678 25130 8730
rect 25142 8678 25194 8730
rect 25206 8678 25258 8730
rect 2964 8619 3016 8628
rect 2964 8585 2973 8619
rect 2973 8585 3007 8619
rect 3007 8585 3016 8619
rect 2964 8576 3016 8585
rect 8116 8576 8168 8628
rect 13084 8619 13136 8628
rect 13084 8585 13093 8619
rect 13093 8585 13127 8619
rect 13127 8585 13136 8619
rect 13084 8576 13136 8585
rect 16580 8576 16632 8628
rect 3240 8440 3292 8492
rect 7104 8440 7156 8492
rect 8576 8440 8628 8492
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 20444 8508 20496 8560
rect 21180 8551 21232 8560
rect 21180 8517 21189 8551
rect 21189 8517 21223 8551
rect 21223 8517 21232 8551
rect 21180 8508 21232 8517
rect 21824 8576 21876 8628
rect 24492 8576 24544 8628
rect 24860 8576 24912 8628
rect 27160 8576 27212 8628
rect 27620 8619 27672 8628
rect 27620 8585 27629 8619
rect 27629 8585 27663 8619
rect 27663 8585 27672 8619
rect 27620 8576 27672 8585
rect 28264 8576 28316 8628
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 13728 8440 13780 8492
rect 20904 8440 20956 8492
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 23296 8440 23348 8492
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 3884 8372 3936 8424
rect 7288 8372 7340 8424
rect 12624 8372 12676 8424
rect 13084 8415 13136 8424
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 24216 8415 24268 8424
rect 13084 8372 13136 8381
rect 24216 8381 24225 8415
rect 24225 8381 24259 8415
rect 24259 8381 24268 8415
rect 24676 8415 24728 8424
rect 24216 8372 24268 8381
rect 24676 8381 24685 8415
rect 24685 8381 24719 8415
rect 24719 8381 24728 8415
rect 24676 8372 24728 8381
rect 26700 8415 26752 8424
rect 26700 8381 26709 8415
rect 26709 8381 26743 8415
rect 26743 8381 26752 8415
rect 26700 8372 26752 8381
rect 27712 8372 27764 8424
rect 1952 8236 2004 8288
rect 7104 8279 7156 8288
rect 7104 8245 7113 8279
rect 7113 8245 7147 8279
rect 7147 8245 7156 8279
rect 7104 8236 7156 8245
rect 9036 8279 9088 8288
rect 9036 8245 9045 8279
rect 9045 8245 9079 8279
rect 9079 8245 9088 8279
rect 9036 8236 9088 8245
rect 19340 8236 19392 8288
rect 20996 8236 21048 8288
rect 3350 8134 3402 8186
rect 3414 8134 3466 8186
rect 3478 8134 3530 8186
rect 3542 8134 3594 8186
rect 3606 8134 3658 8186
rect 8150 8134 8202 8186
rect 8214 8134 8266 8186
rect 8278 8134 8330 8186
rect 8342 8134 8394 8186
rect 8406 8134 8458 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 17750 8134 17802 8186
rect 17814 8134 17866 8186
rect 17878 8134 17930 8186
rect 17942 8134 17994 8186
rect 18006 8134 18058 8186
rect 22550 8134 22602 8186
rect 22614 8134 22666 8186
rect 22678 8134 22730 8186
rect 22742 8134 22794 8186
rect 22806 8134 22858 8186
rect 27350 8134 27402 8186
rect 27414 8134 27466 8186
rect 27478 8134 27530 8186
rect 27542 8134 27594 8186
rect 27606 8134 27658 8186
rect 5540 8032 5592 8084
rect 8576 8075 8628 8084
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 20444 8075 20496 8084
rect 20444 8041 20453 8075
rect 20453 8041 20487 8075
rect 20487 8041 20496 8075
rect 20444 8032 20496 8041
rect 22100 8032 22152 8084
rect 14188 8007 14240 8016
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 1952 7939 2004 7948
rect 1952 7905 1961 7939
rect 1961 7905 1995 7939
rect 1995 7905 2004 7939
rect 1952 7896 2004 7905
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 14188 7973 14197 8007
rect 14197 7973 14231 8007
rect 14231 7973 14240 8007
rect 14188 7964 14240 7973
rect 13728 7939 13780 7948
rect 13728 7905 13737 7939
rect 13737 7905 13771 7939
rect 13771 7905 13780 7939
rect 13728 7896 13780 7905
rect 7104 7828 7156 7880
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 9036 7828 9088 7880
rect 20444 7828 20496 7880
rect 22100 7828 22152 7880
rect 23388 7828 23440 7880
rect 3700 7760 3752 7812
rect 9864 7803 9916 7812
rect 9864 7769 9873 7803
rect 9873 7769 9907 7803
rect 9907 7769 9916 7803
rect 9864 7760 9916 7769
rect 22008 7760 22060 7812
rect 23296 7760 23348 7812
rect 3424 7735 3476 7744
rect 3424 7701 3433 7735
rect 3433 7701 3467 7735
rect 3467 7701 3476 7735
rect 3424 7692 3476 7701
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 14188 7735 14240 7744
rect 14188 7701 14197 7735
rect 14197 7701 14231 7735
rect 14231 7701 14240 7735
rect 14188 7692 14240 7701
rect 22284 7735 22336 7744
rect 22284 7701 22293 7735
rect 22293 7701 22327 7735
rect 22327 7701 22336 7735
rect 22284 7692 22336 7701
rect 23020 7735 23072 7744
rect 23020 7701 23029 7735
rect 23029 7701 23063 7735
rect 23063 7701 23072 7735
rect 23020 7692 23072 7701
rect 5750 7590 5802 7642
rect 5814 7590 5866 7642
rect 5878 7590 5930 7642
rect 5942 7590 5994 7642
rect 6006 7590 6058 7642
rect 10550 7590 10602 7642
rect 10614 7590 10666 7642
rect 10678 7590 10730 7642
rect 10742 7590 10794 7642
rect 10806 7590 10858 7642
rect 15350 7590 15402 7642
rect 15414 7590 15466 7642
rect 15478 7590 15530 7642
rect 15542 7590 15594 7642
rect 15606 7590 15658 7642
rect 20150 7590 20202 7642
rect 20214 7590 20266 7642
rect 20278 7590 20330 7642
rect 20342 7590 20394 7642
rect 20406 7590 20458 7642
rect 24950 7590 25002 7642
rect 25014 7590 25066 7642
rect 25078 7590 25130 7642
rect 25142 7590 25194 7642
rect 25206 7590 25258 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 5540 7488 5592 7540
rect 9680 7488 9732 7540
rect 3424 7352 3476 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 14188 7488 14240 7540
rect 19432 7488 19484 7540
rect 21180 7488 21232 7540
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 23020 7352 23072 7404
rect 9864 7284 9916 7336
rect 19156 7327 19208 7336
rect 19156 7293 19165 7327
rect 19165 7293 19199 7327
rect 19199 7293 19208 7327
rect 19156 7284 19208 7293
rect 19340 7284 19392 7336
rect 22100 7327 22152 7336
rect 22100 7293 22109 7327
rect 22109 7293 22143 7327
rect 22143 7293 22152 7327
rect 22100 7284 22152 7293
rect 7656 7259 7708 7268
rect 7656 7225 7665 7259
rect 7665 7225 7699 7259
rect 7699 7225 7708 7259
rect 7656 7216 7708 7225
rect 22008 7216 22060 7268
rect 23296 7284 23348 7336
rect 18604 7148 18656 7200
rect 3350 7046 3402 7098
rect 3414 7046 3466 7098
rect 3478 7046 3530 7098
rect 3542 7046 3594 7098
rect 3606 7046 3658 7098
rect 8150 7046 8202 7098
rect 8214 7046 8266 7098
rect 8278 7046 8330 7098
rect 8342 7046 8394 7098
rect 8406 7046 8458 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 17750 7046 17802 7098
rect 17814 7046 17866 7098
rect 17878 7046 17930 7098
rect 17942 7046 17994 7098
rect 18006 7046 18058 7098
rect 22550 7046 22602 7098
rect 22614 7046 22666 7098
rect 22678 7046 22730 7098
rect 22742 7046 22794 7098
rect 22806 7046 22858 7098
rect 27350 7046 27402 7098
rect 27414 7046 27466 7098
rect 27478 7046 27530 7098
rect 27542 7046 27594 7098
rect 27606 7046 27658 7098
rect 5540 6944 5592 6996
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 10416 6987 10468 6996
rect 9680 6944 9732 6953
rect 10416 6953 10425 6987
rect 10425 6953 10459 6987
rect 10459 6953 10468 6987
rect 10416 6944 10468 6953
rect 7288 6851 7340 6860
rect 7288 6817 7297 6851
rect 7297 6817 7331 6851
rect 7331 6817 7340 6851
rect 7288 6808 7340 6817
rect 9864 6808 9916 6860
rect 19156 6944 19208 6996
rect 20996 6987 21048 6996
rect 20996 6953 21005 6987
rect 21005 6953 21039 6987
rect 21039 6953 21048 6987
rect 20996 6944 21048 6953
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 8208 6740 8260 6792
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 20996 6808 21048 6860
rect 10416 6740 10468 6749
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 22100 6808 22152 6860
rect 22284 6808 22336 6860
rect 22192 6740 22244 6792
rect 25688 6740 25740 6792
rect 27252 6783 27304 6792
rect 27252 6749 27261 6783
rect 27261 6749 27295 6783
rect 27295 6749 27304 6783
rect 27252 6740 27304 6749
rect 28264 6740 28316 6792
rect 18420 6672 18472 6724
rect 20812 6715 20864 6724
rect 20812 6681 20821 6715
rect 20821 6681 20855 6715
rect 20855 6681 20864 6715
rect 20812 6672 20864 6681
rect 21548 6672 21600 6724
rect 22008 6672 22060 6724
rect 22652 6715 22704 6724
rect 22652 6681 22661 6715
rect 22661 6681 22695 6715
rect 22695 6681 22704 6715
rect 22652 6672 22704 6681
rect 23940 6672 23992 6724
rect 24584 6672 24636 6724
rect 18880 6647 18932 6656
rect 18880 6613 18889 6647
rect 18889 6613 18923 6647
rect 18923 6613 18932 6647
rect 18880 6604 18932 6613
rect 21640 6604 21692 6656
rect 23388 6604 23440 6656
rect 24124 6647 24176 6656
rect 24124 6613 24133 6647
rect 24133 6613 24167 6647
rect 24167 6613 24176 6647
rect 24124 6604 24176 6613
rect 26240 6604 26292 6656
rect 26884 6604 26936 6656
rect 27804 6604 27856 6656
rect 28356 6647 28408 6656
rect 28356 6613 28365 6647
rect 28365 6613 28399 6647
rect 28399 6613 28408 6647
rect 28356 6604 28408 6613
rect 5750 6502 5802 6554
rect 5814 6502 5866 6554
rect 5878 6502 5930 6554
rect 5942 6502 5994 6554
rect 6006 6502 6058 6554
rect 10550 6502 10602 6554
rect 10614 6502 10666 6554
rect 10678 6502 10730 6554
rect 10742 6502 10794 6554
rect 10806 6502 10858 6554
rect 15350 6502 15402 6554
rect 15414 6502 15466 6554
rect 15478 6502 15530 6554
rect 15542 6502 15594 6554
rect 15606 6502 15658 6554
rect 20150 6502 20202 6554
rect 20214 6502 20266 6554
rect 20278 6502 20330 6554
rect 20342 6502 20394 6554
rect 20406 6502 20458 6554
rect 24950 6502 25002 6554
rect 25014 6502 25066 6554
rect 25078 6502 25130 6554
rect 25142 6502 25194 6554
rect 25206 6502 25258 6554
rect 5540 6400 5592 6452
rect 6644 6400 6696 6452
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7656 6264 7708 6316
rect 8208 6264 8260 6316
rect 20812 6400 20864 6452
rect 22192 6400 22244 6452
rect 22652 6400 22704 6452
rect 27252 6443 27304 6452
rect 27252 6409 27261 6443
rect 27261 6409 27295 6443
rect 27295 6409 27304 6443
rect 27252 6400 27304 6409
rect 7288 6128 7340 6180
rect 9864 6264 9916 6316
rect 18604 6264 18656 6316
rect 19248 6264 19300 6316
rect 22100 6332 22152 6384
rect 26240 6375 26292 6384
rect 26240 6341 26249 6375
rect 26249 6341 26283 6375
rect 26283 6341 26292 6375
rect 26240 6332 26292 6341
rect 20720 6264 20772 6316
rect 21548 6264 21600 6316
rect 21640 6264 21692 6316
rect 24584 6264 24636 6316
rect 12624 6103 12676 6112
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 20996 6196 21048 6248
rect 12624 6060 12676 6069
rect 19524 6060 19576 6112
rect 25228 6060 25280 6112
rect 26608 6196 26660 6248
rect 27804 6239 27856 6248
rect 27804 6205 27813 6239
rect 27813 6205 27847 6239
rect 27847 6205 27856 6239
rect 27804 6196 27856 6205
rect 28356 6128 28408 6180
rect 27896 6060 27948 6112
rect 3350 5958 3402 6010
rect 3414 5958 3466 6010
rect 3478 5958 3530 6010
rect 3542 5958 3594 6010
rect 3606 5958 3658 6010
rect 8150 5958 8202 6010
rect 8214 5958 8266 6010
rect 8278 5958 8330 6010
rect 8342 5958 8394 6010
rect 8406 5958 8458 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 17750 5958 17802 6010
rect 17814 5958 17866 6010
rect 17878 5958 17930 6010
rect 17942 5958 17994 6010
rect 18006 5958 18058 6010
rect 22550 5958 22602 6010
rect 22614 5958 22666 6010
rect 22678 5958 22730 6010
rect 22742 5958 22794 6010
rect 22806 5958 22858 6010
rect 27350 5958 27402 6010
rect 27414 5958 27466 6010
rect 27478 5958 27530 6010
rect 27542 5958 27594 6010
rect 27606 5958 27658 6010
rect 7288 5831 7340 5840
rect 7288 5797 7297 5831
rect 7297 5797 7331 5831
rect 7331 5797 7340 5831
rect 7288 5788 7340 5797
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 12624 5899 12676 5908
rect 11704 5831 11756 5840
rect 11704 5797 11713 5831
rect 11713 5797 11747 5831
rect 11747 5797 11756 5831
rect 12624 5865 12633 5899
rect 12633 5865 12667 5899
rect 12667 5865 12676 5899
rect 12624 5856 12676 5865
rect 24676 5899 24728 5908
rect 24676 5865 24685 5899
rect 24685 5865 24719 5899
rect 24719 5865 24728 5899
rect 24676 5856 24728 5865
rect 25688 5899 25740 5908
rect 25688 5865 25697 5899
rect 25697 5865 25731 5899
rect 25731 5865 25740 5899
rect 25688 5856 25740 5865
rect 28356 5899 28408 5908
rect 28356 5865 28365 5899
rect 28365 5865 28399 5899
rect 28399 5865 28408 5899
rect 28356 5856 28408 5865
rect 11704 5788 11756 5797
rect 9864 5720 9916 5772
rect 10968 5720 11020 5772
rect 19432 5788 19484 5840
rect 19248 5720 19300 5772
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 19524 5652 19576 5704
rect 25228 5763 25280 5772
rect 25228 5729 25237 5763
rect 25237 5729 25271 5763
rect 25271 5729 25280 5763
rect 25228 5720 25280 5729
rect 26884 5763 26936 5772
rect 26884 5729 26893 5763
rect 26893 5729 26927 5763
rect 26927 5729 26936 5763
rect 26884 5720 26936 5729
rect 24124 5652 24176 5704
rect 26608 5695 26660 5704
rect 26608 5661 26617 5695
rect 26617 5661 26651 5695
rect 26651 5661 26660 5695
rect 26608 5652 26660 5661
rect 27896 5584 27948 5636
rect 6644 5516 6696 5525
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 20720 5516 20772 5568
rect 5750 5414 5802 5466
rect 5814 5414 5866 5466
rect 5878 5414 5930 5466
rect 5942 5414 5994 5466
rect 6006 5414 6058 5466
rect 10550 5414 10602 5466
rect 10614 5414 10666 5466
rect 10678 5414 10730 5466
rect 10742 5414 10794 5466
rect 10806 5414 10858 5466
rect 15350 5414 15402 5466
rect 15414 5414 15466 5466
rect 15478 5414 15530 5466
rect 15542 5414 15594 5466
rect 15606 5414 15658 5466
rect 20150 5414 20202 5466
rect 20214 5414 20266 5466
rect 20278 5414 20330 5466
rect 20342 5414 20394 5466
rect 20406 5414 20458 5466
rect 24950 5414 25002 5466
rect 25014 5414 25066 5466
rect 25078 5414 25130 5466
rect 25142 5414 25194 5466
rect 25206 5414 25258 5466
rect 11704 5355 11756 5364
rect 10600 5176 10652 5228
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 20720 5312 20772 5364
rect 10968 5176 11020 5228
rect 19340 5244 19392 5296
rect 19616 5244 19668 5296
rect 19432 5108 19484 5160
rect 23572 4972 23624 5024
rect 3350 4870 3402 4922
rect 3414 4870 3466 4922
rect 3478 4870 3530 4922
rect 3542 4870 3594 4922
rect 3606 4870 3658 4922
rect 8150 4870 8202 4922
rect 8214 4870 8266 4922
rect 8278 4870 8330 4922
rect 8342 4870 8394 4922
rect 8406 4870 8458 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 17750 4870 17802 4922
rect 17814 4870 17866 4922
rect 17878 4870 17930 4922
rect 17942 4870 17994 4922
rect 18006 4870 18058 4922
rect 22550 4870 22602 4922
rect 22614 4870 22666 4922
rect 22678 4870 22730 4922
rect 22742 4870 22794 4922
rect 22806 4870 22858 4922
rect 27350 4870 27402 4922
rect 27414 4870 27466 4922
rect 27478 4870 27530 4922
rect 27542 4870 27594 4922
rect 27606 4870 27658 4922
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 23572 4632 23624 4684
rect 24676 4632 24728 4684
rect 20720 4564 20772 4616
rect 23020 4564 23072 4616
rect 26240 4564 26292 4616
rect 26608 4564 26660 4616
rect 26976 4539 27028 4548
rect 26976 4505 26985 4539
rect 26985 4505 27019 4539
rect 27019 4505 27028 4539
rect 26976 4496 27028 4505
rect 27988 4496 28040 4548
rect 3148 4428 3200 4480
rect 22100 4471 22152 4480
rect 22100 4437 22109 4471
rect 22109 4437 22143 4471
rect 22143 4437 22152 4471
rect 22100 4428 22152 4437
rect 23020 4428 23072 4480
rect 23204 4428 23256 4480
rect 23572 4471 23624 4480
rect 23572 4437 23581 4471
rect 23581 4437 23615 4471
rect 23615 4437 23624 4471
rect 28448 4471 28500 4480
rect 23572 4428 23624 4437
rect 28448 4437 28457 4471
rect 28457 4437 28491 4471
rect 28491 4437 28500 4471
rect 28448 4428 28500 4437
rect 5750 4326 5802 4378
rect 5814 4326 5866 4378
rect 5878 4326 5930 4378
rect 5942 4326 5994 4378
rect 6006 4326 6058 4378
rect 10550 4326 10602 4378
rect 10614 4326 10666 4378
rect 10678 4326 10730 4378
rect 10742 4326 10794 4378
rect 10806 4326 10858 4378
rect 15350 4326 15402 4378
rect 15414 4326 15466 4378
rect 15478 4326 15530 4378
rect 15542 4326 15594 4378
rect 15606 4326 15658 4378
rect 20150 4326 20202 4378
rect 20214 4326 20266 4378
rect 20278 4326 20330 4378
rect 20342 4326 20394 4378
rect 20406 4326 20458 4378
rect 24950 4326 25002 4378
rect 25014 4326 25066 4378
rect 25078 4326 25130 4378
rect 25142 4326 25194 4378
rect 25206 4326 25258 4378
rect 10232 4224 10284 4276
rect 28448 4224 28500 4276
rect 11612 4156 11664 4208
rect 19616 4156 19668 4208
rect 20076 4156 20128 4208
rect 21088 4088 21140 4140
rect 22100 4088 22152 4140
rect 23204 4131 23256 4140
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 25412 4131 25464 4140
rect 25412 4097 25421 4131
rect 25421 4097 25455 4131
rect 25455 4097 25464 4131
rect 25412 4088 25464 4097
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 3148 4063 3200 4072
rect 3148 4029 3157 4063
rect 3157 4029 3191 4063
rect 3191 4029 3200 4063
rect 3148 4020 3200 4029
rect 21640 3952 21692 4004
rect 27804 4063 27856 4072
rect 27804 4029 27813 4063
rect 27813 4029 27847 4063
rect 27847 4029 27856 4063
rect 27804 4020 27856 4029
rect 23388 3995 23440 4004
rect 23388 3961 23397 3995
rect 23397 3961 23431 3995
rect 23431 3961 23440 3995
rect 23388 3952 23440 3961
rect 25780 3952 25832 4004
rect 2504 3927 2556 3936
rect 2504 3893 2513 3927
rect 2513 3893 2547 3927
rect 2547 3893 2556 3927
rect 2504 3884 2556 3893
rect 3700 3884 3752 3936
rect 18788 3884 18840 3936
rect 23848 3884 23900 3936
rect 25136 3884 25188 3936
rect 27252 3927 27304 3936
rect 27252 3893 27261 3927
rect 27261 3893 27295 3927
rect 27295 3893 27304 3927
rect 27252 3884 27304 3893
rect 3350 3782 3402 3834
rect 3414 3782 3466 3834
rect 3478 3782 3530 3834
rect 3542 3782 3594 3834
rect 3606 3782 3658 3834
rect 8150 3782 8202 3834
rect 8214 3782 8266 3834
rect 8278 3782 8330 3834
rect 8342 3782 8394 3834
rect 8406 3782 8458 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 17750 3782 17802 3834
rect 17814 3782 17866 3834
rect 17878 3782 17930 3834
rect 17942 3782 17994 3834
rect 18006 3782 18058 3834
rect 22550 3782 22602 3834
rect 22614 3782 22666 3834
rect 22678 3782 22730 3834
rect 22742 3782 22794 3834
rect 22806 3782 22858 3834
rect 27350 3782 27402 3834
rect 27414 3782 27466 3834
rect 27478 3782 27530 3834
rect 27542 3782 27594 3834
rect 27606 3782 27658 3834
rect 2964 3680 3016 3732
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 23020 3680 23072 3732
rect 26976 3680 27028 3732
rect 28356 3723 28408 3732
rect 28356 3689 28365 3723
rect 28365 3689 28399 3723
rect 28399 3689 28408 3723
rect 28356 3680 28408 3689
rect 26240 3612 26292 3664
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 3792 3544 3844 3596
rect 13820 3544 13872 3596
rect 19340 3587 19392 3596
rect 3056 3476 3108 3528
rect 3884 3519 3936 3528
rect 3884 3485 3893 3519
rect 3893 3485 3927 3519
rect 3927 3485 3936 3519
rect 3884 3476 3936 3485
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 18788 3519 18840 3528
rect 18788 3485 18797 3519
rect 18797 3485 18831 3519
rect 18831 3485 18840 3519
rect 18788 3476 18840 3485
rect 18880 3519 18932 3528
rect 18880 3485 18894 3519
rect 18894 3485 18928 3519
rect 18928 3485 18932 3519
rect 18880 3476 18932 3485
rect 2228 3408 2280 3460
rect 18236 3451 18288 3460
rect 18236 3417 18245 3451
rect 18245 3417 18279 3451
rect 18279 3417 18288 3451
rect 18236 3408 18288 3417
rect 19340 3553 19349 3587
rect 19349 3553 19383 3587
rect 19383 3553 19392 3587
rect 19340 3544 19392 3553
rect 21640 3587 21692 3596
rect 21640 3553 21649 3587
rect 21649 3553 21683 3587
rect 21683 3553 21692 3587
rect 21640 3544 21692 3553
rect 22284 3544 22336 3596
rect 27252 3519 27304 3528
rect 27252 3485 27261 3519
rect 27261 3485 27295 3519
rect 27295 3485 27304 3519
rect 27252 3476 27304 3485
rect 28448 3476 28500 3528
rect 20076 3408 20128 3460
rect 23848 3408 23900 3460
rect 25136 3451 25188 3460
rect 25136 3417 25145 3451
rect 25145 3417 25179 3451
rect 25179 3417 25188 3451
rect 25136 3408 25188 3417
rect 26424 3408 26476 3460
rect 27896 3408 27948 3460
rect 1768 3340 1820 3392
rect 2964 3340 3016 3392
rect 21088 3340 21140 3392
rect 26148 3340 26200 3392
rect 26608 3383 26660 3392
rect 26608 3349 26617 3383
rect 26617 3349 26651 3383
rect 26651 3349 26660 3383
rect 26608 3340 26660 3349
rect 5750 3238 5802 3290
rect 5814 3238 5866 3290
rect 5878 3238 5930 3290
rect 5942 3238 5994 3290
rect 6006 3238 6058 3290
rect 10550 3238 10602 3290
rect 10614 3238 10666 3290
rect 10678 3238 10730 3290
rect 10742 3238 10794 3290
rect 10806 3238 10858 3290
rect 15350 3238 15402 3290
rect 15414 3238 15466 3290
rect 15478 3238 15530 3290
rect 15542 3238 15594 3290
rect 15606 3238 15658 3290
rect 20150 3238 20202 3290
rect 20214 3238 20266 3290
rect 20278 3238 20330 3290
rect 20342 3238 20394 3290
rect 20406 3238 20458 3290
rect 24950 3238 25002 3290
rect 25014 3238 25066 3290
rect 25078 3238 25130 3290
rect 25142 3238 25194 3290
rect 25206 3238 25258 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 3056 3136 3108 3188
rect 19708 3179 19760 3188
rect 19708 3145 19717 3179
rect 19717 3145 19751 3179
rect 19751 3145 19760 3179
rect 19708 3136 19760 3145
rect 20076 3111 20128 3120
rect 20076 3077 20085 3111
rect 20085 3077 20119 3111
rect 20119 3077 20128 3111
rect 20076 3068 20128 3077
rect 23388 3136 23440 3188
rect 23572 3136 23624 3188
rect 25412 3179 25464 3188
rect 25412 3145 25421 3179
rect 25421 3145 25455 3179
rect 25455 3145 25464 3179
rect 25412 3136 25464 3145
rect 25780 3179 25832 3188
rect 25780 3145 25789 3179
rect 25789 3145 25823 3179
rect 25823 3145 25832 3179
rect 25780 3136 25832 3145
rect 23848 3068 23900 3120
rect 26424 3068 26476 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 2504 3000 2556 3052
rect 3700 3000 3752 3052
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 26608 3000 26660 3052
rect 18880 2932 18932 2984
rect 19708 2864 19760 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 3350 2694 3402 2746
rect 3414 2694 3466 2746
rect 3478 2694 3530 2746
rect 3542 2694 3594 2746
rect 3606 2694 3658 2746
rect 8150 2694 8202 2746
rect 8214 2694 8266 2746
rect 8278 2694 8330 2746
rect 8342 2694 8394 2746
rect 8406 2694 8458 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 17750 2694 17802 2746
rect 17814 2694 17866 2746
rect 17878 2694 17930 2746
rect 17942 2694 17994 2746
rect 18006 2694 18058 2746
rect 22550 2694 22602 2746
rect 22614 2694 22666 2746
rect 22678 2694 22730 2746
rect 22742 2694 22794 2746
rect 22806 2694 22858 2746
rect 27350 2694 27402 2746
rect 27414 2694 27466 2746
rect 27478 2694 27530 2746
rect 27542 2694 27594 2746
rect 27606 2694 27658 2746
rect 11612 2635 11664 2644
rect 11612 2601 11621 2635
rect 11621 2601 11655 2635
rect 11655 2601 11664 2635
rect 11612 2592 11664 2601
rect 18512 2592 18564 2644
rect 11244 2388 11296 2440
rect 18696 2388 18748 2440
rect 26240 2431 26292 2440
rect 26240 2397 26249 2431
rect 26249 2397 26283 2431
rect 26283 2397 26292 2431
rect 26240 2388 26292 2397
rect 26608 2388 26660 2440
rect 26148 2252 26200 2304
rect 28356 2295 28408 2304
rect 28356 2261 28365 2295
rect 28365 2261 28399 2295
rect 28399 2261 28408 2295
rect 28356 2252 28408 2261
rect 5750 2150 5802 2202
rect 5814 2150 5866 2202
rect 5878 2150 5930 2202
rect 5942 2150 5994 2202
rect 6006 2150 6058 2202
rect 10550 2150 10602 2202
rect 10614 2150 10666 2202
rect 10678 2150 10730 2202
rect 10742 2150 10794 2202
rect 10806 2150 10858 2202
rect 15350 2150 15402 2202
rect 15414 2150 15466 2202
rect 15478 2150 15530 2202
rect 15542 2150 15594 2202
rect 15606 2150 15658 2202
rect 20150 2150 20202 2202
rect 20214 2150 20266 2202
rect 20278 2150 20330 2202
rect 20342 2150 20394 2202
rect 20406 2150 20458 2202
rect 24950 2150 25002 2202
rect 25014 2150 25066 2202
rect 25078 2150 25130 2202
rect 25142 2150 25194 2202
rect 25206 2150 25258 2202
<< metal2 >>
rect 28354 28384 28410 28393
rect 28354 28319 28410 28328
rect 3350 27772 3658 27781
rect 3350 27770 3356 27772
rect 3412 27770 3436 27772
rect 3492 27770 3516 27772
rect 3572 27770 3596 27772
rect 3652 27770 3658 27772
rect 3412 27718 3414 27770
rect 3594 27718 3596 27770
rect 3350 27716 3356 27718
rect 3412 27716 3436 27718
rect 3492 27716 3516 27718
rect 3572 27716 3596 27718
rect 3652 27716 3658 27718
rect 3350 27707 3658 27716
rect 8150 27772 8458 27781
rect 8150 27770 8156 27772
rect 8212 27770 8236 27772
rect 8292 27770 8316 27772
rect 8372 27770 8396 27772
rect 8452 27770 8458 27772
rect 8212 27718 8214 27770
rect 8394 27718 8396 27770
rect 8150 27716 8156 27718
rect 8212 27716 8236 27718
rect 8292 27716 8316 27718
rect 8372 27716 8396 27718
rect 8452 27716 8458 27718
rect 8150 27707 8458 27716
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 17750 27772 18058 27781
rect 17750 27770 17756 27772
rect 17812 27770 17836 27772
rect 17892 27770 17916 27772
rect 17972 27770 17996 27772
rect 18052 27770 18058 27772
rect 17812 27718 17814 27770
rect 17994 27718 17996 27770
rect 17750 27716 17756 27718
rect 17812 27716 17836 27718
rect 17892 27716 17916 27718
rect 17972 27716 17996 27718
rect 18052 27716 18058 27718
rect 17750 27707 18058 27716
rect 22550 27772 22858 27781
rect 22550 27770 22556 27772
rect 22612 27770 22636 27772
rect 22692 27770 22716 27772
rect 22772 27770 22796 27772
rect 22852 27770 22858 27772
rect 22612 27718 22614 27770
rect 22794 27718 22796 27770
rect 22550 27716 22556 27718
rect 22612 27716 22636 27718
rect 22692 27716 22716 27718
rect 22772 27716 22796 27718
rect 22852 27716 22858 27718
rect 22550 27707 22858 27716
rect 27350 27772 27658 27781
rect 27350 27770 27356 27772
rect 27412 27770 27436 27772
rect 27492 27770 27516 27772
rect 27572 27770 27596 27772
rect 27652 27770 27658 27772
rect 27412 27718 27414 27770
rect 27594 27718 27596 27770
rect 27350 27716 27356 27718
rect 27412 27716 27436 27718
rect 27492 27716 27516 27718
rect 27572 27716 27596 27718
rect 27652 27716 27658 27718
rect 27350 27707 27658 27716
rect 28368 27606 28396 28319
rect 28356 27600 28408 27606
rect 28356 27542 28408 27548
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 27804 27464 27856 27470
rect 27804 27406 27856 27412
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1596 27169 1624 27270
rect 1582 27160 1638 27169
rect 1582 27095 1638 27104
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22273 1624 22374
rect 1582 22264 1638 22273
rect 1582 22199 1638 22208
rect 3068 21690 3096 27406
rect 5750 27228 6058 27237
rect 5750 27226 5756 27228
rect 5812 27226 5836 27228
rect 5892 27226 5916 27228
rect 5972 27226 5996 27228
rect 6052 27226 6058 27228
rect 5812 27174 5814 27226
rect 5994 27174 5996 27226
rect 5750 27172 5756 27174
rect 5812 27172 5836 27174
rect 5892 27172 5916 27174
rect 5972 27172 5996 27174
rect 6052 27172 6058 27174
rect 5750 27163 6058 27172
rect 10550 27228 10858 27237
rect 10550 27226 10556 27228
rect 10612 27226 10636 27228
rect 10692 27226 10716 27228
rect 10772 27226 10796 27228
rect 10852 27226 10858 27228
rect 10612 27174 10614 27226
rect 10794 27174 10796 27226
rect 10550 27172 10556 27174
rect 10612 27172 10636 27174
rect 10692 27172 10716 27174
rect 10772 27172 10796 27174
rect 10852 27172 10858 27174
rect 10550 27163 10858 27172
rect 15350 27228 15658 27237
rect 15350 27226 15356 27228
rect 15412 27226 15436 27228
rect 15492 27226 15516 27228
rect 15572 27226 15596 27228
rect 15652 27226 15658 27228
rect 15412 27174 15414 27226
rect 15594 27174 15596 27226
rect 15350 27172 15356 27174
rect 15412 27172 15436 27174
rect 15492 27172 15516 27174
rect 15572 27172 15596 27174
rect 15652 27172 15658 27174
rect 15350 27163 15658 27172
rect 20150 27228 20458 27237
rect 20150 27226 20156 27228
rect 20212 27226 20236 27228
rect 20292 27226 20316 27228
rect 20372 27226 20396 27228
rect 20452 27226 20458 27228
rect 20212 27174 20214 27226
rect 20394 27174 20396 27226
rect 20150 27172 20156 27174
rect 20212 27172 20236 27174
rect 20292 27172 20316 27174
rect 20372 27172 20396 27174
rect 20452 27172 20458 27174
rect 20150 27163 20458 27172
rect 24950 27228 25258 27237
rect 24950 27226 24956 27228
rect 25012 27226 25036 27228
rect 25092 27226 25116 27228
rect 25172 27226 25196 27228
rect 25252 27226 25258 27228
rect 25012 27174 25014 27226
rect 25194 27174 25196 27226
rect 24950 27172 24956 27174
rect 25012 27172 25036 27174
rect 25092 27172 25116 27174
rect 25172 27172 25196 27174
rect 25252 27172 25258 27174
rect 24950 27163 25258 27172
rect 3350 26684 3658 26693
rect 3350 26682 3356 26684
rect 3412 26682 3436 26684
rect 3492 26682 3516 26684
rect 3572 26682 3596 26684
rect 3652 26682 3658 26684
rect 3412 26630 3414 26682
rect 3594 26630 3596 26682
rect 3350 26628 3356 26630
rect 3412 26628 3436 26630
rect 3492 26628 3516 26630
rect 3572 26628 3596 26630
rect 3652 26628 3658 26630
rect 3350 26619 3658 26628
rect 8150 26684 8458 26693
rect 8150 26682 8156 26684
rect 8212 26682 8236 26684
rect 8292 26682 8316 26684
rect 8372 26682 8396 26684
rect 8452 26682 8458 26684
rect 8212 26630 8214 26682
rect 8394 26630 8396 26682
rect 8150 26628 8156 26630
rect 8212 26628 8236 26630
rect 8292 26628 8316 26630
rect 8372 26628 8396 26630
rect 8452 26628 8458 26630
rect 8150 26619 8458 26628
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 17750 26684 18058 26693
rect 17750 26682 17756 26684
rect 17812 26682 17836 26684
rect 17892 26682 17916 26684
rect 17972 26682 17996 26684
rect 18052 26682 18058 26684
rect 17812 26630 17814 26682
rect 17994 26630 17996 26682
rect 17750 26628 17756 26630
rect 17812 26628 17836 26630
rect 17892 26628 17916 26630
rect 17972 26628 17996 26630
rect 18052 26628 18058 26630
rect 17750 26619 18058 26628
rect 22550 26684 22858 26693
rect 22550 26682 22556 26684
rect 22612 26682 22636 26684
rect 22692 26682 22716 26684
rect 22772 26682 22796 26684
rect 22852 26682 22858 26684
rect 22612 26630 22614 26682
rect 22794 26630 22796 26682
rect 22550 26628 22556 26630
rect 22612 26628 22636 26630
rect 22692 26628 22716 26630
rect 22772 26628 22796 26630
rect 22852 26628 22858 26630
rect 22550 26619 22858 26628
rect 27350 26684 27658 26693
rect 27350 26682 27356 26684
rect 27412 26682 27436 26684
rect 27492 26682 27516 26684
rect 27572 26682 27596 26684
rect 27652 26682 27658 26684
rect 27412 26630 27414 26682
rect 27594 26630 27596 26682
rect 27350 26628 27356 26630
rect 27412 26628 27436 26630
rect 27492 26628 27516 26630
rect 27572 26628 27596 26630
rect 27652 26628 27658 26630
rect 27350 26619 27658 26628
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 5750 26140 6058 26149
rect 5750 26138 5756 26140
rect 5812 26138 5836 26140
rect 5892 26138 5916 26140
rect 5972 26138 5996 26140
rect 6052 26138 6058 26140
rect 5812 26086 5814 26138
rect 5994 26086 5996 26138
rect 5750 26084 5756 26086
rect 5812 26084 5836 26086
rect 5892 26084 5916 26086
rect 5972 26084 5996 26086
rect 6052 26084 6058 26086
rect 5750 26075 6058 26084
rect 10550 26140 10858 26149
rect 10550 26138 10556 26140
rect 10612 26138 10636 26140
rect 10692 26138 10716 26140
rect 10772 26138 10796 26140
rect 10852 26138 10858 26140
rect 10612 26086 10614 26138
rect 10794 26086 10796 26138
rect 10550 26084 10556 26086
rect 10612 26084 10636 26086
rect 10692 26084 10716 26086
rect 10772 26084 10796 26086
rect 10852 26084 10858 26086
rect 10550 26075 10858 26084
rect 15350 26140 15658 26149
rect 15350 26138 15356 26140
rect 15412 26138 15436 26140
rect 15492 26138 15516 26140
rect 15572 26138 15596 26140
rect 15652 26138 15658 26140
rect 15412 26086 15414 26138
rect 15594 26086 15596 26138
rect 15350 26084 15356 26086
rect 15412 26084 15436 26086
rect 15492 26084 15516 26086
rect 15572 26084 15596 26086
rect 15652 26084 15658 26086
rect 15350 26075 15658 26084
rect 20150 26140 20458 26149
rect 20150 26138 20156 26140
rect 20212 26138 20236 26140
rect 20292 26138 20316 26140
rect 20372 26138 20396 26140
rect 20452 26138 20458 26140
rect 20212 26086 20214 26138
rect 20394 26086 20396 26138
rect 20150 26084 20156 26086
rect 20212 26084 20236 26086
rect 20292 26084 20316 26086
rect 20372 26084 20396 26086
rect 20452 26084 20458 26086
rect 20150 26075 20458 26084
rect 24950 26140 25258 26149
rect 24950 26138 24956 26140
rect 25012 26138 25036 26140
rect 25092 26138 25116 26140
rect 25172 26138 25196 26140
rect 25252 26138 25258 26140
rect 25012 26086 25014 26138
rect 25194 26086 25196 26138
rect 24950 26084 24956 26086
rect 25012 26084 25036 26086
rect 25092 26084 25116 26086
rect 25172 26084 25196 26086
rect 25252 26084 25258 26086
rect 24950 26075 25258 26084
rect 3350 25596 3658 25605
rect 3350 25594 3356 25596
rect 3412 25594 3436 25596
rect 3492 25594 3516 25596
rect 3572 25594 3596 25596
rect 3652 25594 3658 25596
rect 3412 25542 3414 25594
rect 3594 25542 3596 25594
rect 3350 25540 3356 25542
rect 3412 25540 3436 25542
rect 3492 25540 3516 25542
rect 3572 25540 3596 25542
rect 3652 25540 3658 25542
rect 3350 25531 3658 25540
rect 8150 25596 8458 25605
rect 8150 25594 8156 25596
rect 8212 25594 8236 25596
rect 8292 25594 8316 25596
rect 8372 25594 8396 25596
rect 8452 25594 8458 25596
rect 8212 25542 8214 25594
rect 8394 25542 8396 25594
rect 8150 25540 8156 25542
rect 8212 25540 8236 25542
rect 8292 25540 8316 25542
rect 8372 25540 8396 25542
rect 8452 25540 8458 25542
rect 8150 25531 8458 25540
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 17750 25596 18058 25605
rect 17750 25594 17756 25596
rect 17812 25594 17836 25596
rect 17892 25594 17916 25596
rect 17972 25594 17996 25596
rect 18052 25594 18058 25596
rect 17812 25542 17814 25594
rect 17994 25542 17996 25594
rect 17750 25540 17756 25542
rect 17812 25540 17836 25542
rect 17892 25540 17916 25542
rect 17972 25540 17996 25542
rect 18052 25540 18058 25542
rect 17750 25531 18058 25540
rect 22550 25596 22858 25605
rect 22550 25594 22556 25596
rect 22612 25594 22636 25596
rect 22692 25594 22716 25596
rect 22772 25594 22796 25596
rect 22852 25594 22858 25596
rect 22612 25542 22614 25594
rect 22794 25542 22796 25594
rect 22550 25540 22556 25542
rect 22612 25540 22636 25542
rect 22692 25540 22716 25542
rect 22772 25540 22796 25542
rect 22852 25540 22858 25542
rect 22550 25531 22858 25540
rect 27350 25596 27658 25605
rect 27350 25594 27356 25596
rect 27412 25594 27436 25596
rect 27492 25594 27516 25596
rect 27572 25594 27596 25596
rect 27652 25594 27658 25596
rect 27412 25542 27414 25594
rect 27594 25542 27596 25594
rect 27350 25540 27356 25542
rect 27412 25540 27436 25542
rect 27492 25540 27516 25542
rect 27572 25540 27596 25542
rect 27652 25540 27658 25542
rect 27350 25531 27658 25540
rect 5750 25052 6058 25061
rect 5750 25050 5756 25052
rect 5812 25050 5836 25052
rect 5892 25050 5916 25052
rect 5972 25050 5996 25052
rect 6052 25050 6058 25052
rect 5812 24998 5814 25050
rect 5994 24998 5996 25050
rect 5750 24996 5756 24998
rect 5812 24996 5836 24998
rect 5892 24996 5916 24998
rect 5972 24996 5996 24998
rect 6052 24996 6058 24998
rect 5750 24987 6058 24996
rect 10550 25052 10858 25061
rect 10550 25050 10556 25052
rect 10612 25050 10636 25052
rect 10692 25050 10716 25052
rect 10772 25050 10796 25052
rect 10852 25050 10858 25052
rect 10612 24998 10614 25050
rect 10794 24998 10796 25050
rect 10550 24996 10556 24998
rect 10612 24996 10636 24998
rect 10692 24996 10716 24998
rect 10772 24996 10796 24998
rect 10852 24996 10858 24998
rect 10550 24987 10858 24996
rect 15350 25052 15658 25061
rect 15350 25050 15356 25052
rect 15412 25050 15436 25052
rect 15492 25050 15516 25052
rect 15572 25050 15596 25052
rect 15652 25050 15658 25052
rect 15412 24998 15414 25050
rect 15594 24998 15596 25050
rect 15350 24996 15356 24998
rect 15412 24996 15436 24998
rect 15492 24996 15516 24998
rect 15572 24996 15596 24998
rect 15652 24996 15658 24998
rect 15350 24987 15658 24996
rect 20150 25052 20458 25061
rect 20150 25050 20156 25052
rect 20212 25050 20236 25052
rect 20292 25050 20316 25052
rect 20372 25050 20396 25052
rect 20452 25050 20458 25052
rect 20212 24998 20214 25050
rect 20394 24998 20396 25050
rect 20150 24996 20156 24998
rect 20212 24996 20236 24998
rect 20292 24996 20316 24998
rect 20372 24996 20396 24998
rect 20452 24996 20458 24998
rect 20150 24987 20458 24996
rect 24950 25052 25258 25061
rect 24950 25050 24956 25052
rect 25012 25050 25036 25052
rect 25092 25050 25116 25052
rect 25172 25050 25196 25052
rect 25252 25050 25258 25052
rect 25012 24998 25014 25050
rect 25194 24998 25196 25050
rect 24950 24996 24956 24998
rect 25012 24996 25036 24998
rect 25092 24996 25116 24998
rect 25172 24996 25196 24998
rect 25252 24996 25258 24998
rect 24950 24987 25258 24996
rect 3350 24508 3658 24517
rect 3350 24506 3356 24508
rect 3412 24506 3436 24508
rect 3492 24506 3516 24508
rect 3572 24506 3596 24508
rect 3652 24506 3658 24508
rect 3412 24454 3414 24506
rect 3594 24454 3596 24506
rect 3350 24452 3356 24454
rect 3412 24452 3436 24454
rect 3492 24452 3516 24454
rect 3572 24452 3596 24454
rect 3652 24452 3658 24454
rect 3350 24443 3658 24452
rect 8150 24508 8458 24517
rect 8150 24506 8156 24508
rect 8212 24506 8236 24508
rect 8292 24506 8316 24508
rect 8372 24506 8396 24508
rect 8452 24506 8458 24508
rect 8212 24454 8214 24506
rect 8394 24454 8396 24506
rect 8150 24452 8156 24454
rect 8212 24452 8236 24454
rect 8292 24452 8316 24454
rect 8372 24452 8396 24454
rect 8452 24452 8458 24454
rect 8150 24443 8458 24452
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 17750 24508 18058 24517
rect 17750 24506 17756 24508
rect 17812 24506 17836 24508
rect 17892 24506 17916 24508
rect 17972 24506 17996 24508
rect 18052 24506 18058 24508
rect 17812 24454 17814 24506
rect 17994 24454 17996 24506
rect 17750 24452 17756 24454
rect 17812 24452 17836 24454
rect 17892 24452 17916 24454
rect 17972 24452 17996 24454
rect 18052 24452 18058 24454
rect 17750 24443 18058 24452
rect 22550 24508 22858 24517
rect 22550 24506 22556 24508
rect 22612 24506 22636 24508
rect 22692 24506 22716 24508
rect 22772 24506 22796 24508
rect 22852 24506 22858 24508
rect 22612 24454 22614 24506
rect 22794 24454 22796 24506
rect 22550 24452 22556 24454
rect 22612 24452 22636 24454
rect 22692 24452 22716 24454
rect 22772 24452 22796 24454
rect 22852 24452 22858 24454
rect 22550 24443 22858 24452
rect 27350 24508 27658 24517
rect 27350 24506 27356 24508
rect 27412 24506 27436 24508
rect 27492 24506 27516 24508
rect 27572 24506 27596 24508
rect 27652 24506 27658 24508
rect 27412 24454 27414 24506
rect 27594 24454 27596 24506
rect 27350 24452 27356 24454
rect 27412 24452 27436 24454
rect 27492 24452 27516 24454
rect 27572 24452 27596 24454
rect 27652 24452 27658 24454
rect 27350 24443 27658 24452
rect 5750 23964 6058 23973
rect 5750 23962 5756 23964
rect 5812 23962 5836 23964
rect 5892 23962 5916 23964
rect 5972 23962 5996 23964
rect 6052 23962 6058 23964
rect 5812 23910 5814 23962
rect 5994 23910 5996 23962
rect 5750 23908 5756 23910
rect 5812 23908 5836 23910
rect 5892 23908 5916 23910
rect 5972 23908 5996 23910
rect 6052 23908 6058 23910
rect 5750 23899 6058 23908
rect 10550 23964 10858 23973
rect 10550 23962 10556 23964
rect 10612 23962 10636 23964
rect 10692 23962 10716 23964
rect 10772 23962 10796 23964
rect 10852 23962 10858 23964
rect 10612 23910 10614 23962
rect 10794 23910 10796 23962
rect 10550 23908 10556 23910
rect 10612 23908 10636 23910
rect 10692 23908 10716 23910
rect 10772 23908 10796 23910
rect 10852 23908 10858 23910
rect 10550 23899 10858 23908
rect 15350 23964 15658 23973
rect 15350 23962 15356 23964
rect 15412 23962 15436 23964
rect 15492 23962 15516 23964
rect 15572 23962 15596 23964
rect 15652 23962 15658 23964
rect 15412 23910 15414 23962
rect 15594 23910 15596 23962
rect 15350 23908 15356 23910
rect 15412 23908 15436 23910
rect 15492 23908 15516 23910
rect 15572 23908 15596 23910
rect 15652 23908 15658 23910
rect 15350 23899 15658 23908
rect 20150 23964 20458 23973
rect 20150 23962 20156 23964
rect 20212 23962 20236 23964
rect 20292 23962 20316 23964
rect 20372 23962 20396 23964
rect 20452 23962 20458 23964
rect 20212 23910 20214 23962
rect 20394 23910 20396 23962
rect 20150 23908 20156 23910
rect 20212 23908 20236 23910
rect 20292 23908 20316 23910
rect 20372 23908 20396 23910
rect 20452 23908 20458 23910
rect 20150 23899 20458 23908
rect 24950 23964 25258 23973
rect 24950 23962 24956 23964
rect 25012 23962 25036 23964
rect 25092 23962 25116 23964
rect 25172 23962 25196 23964
rect 25252 23962 25258 23964
rect 25012 23910 25014 23962
rect 25194 23910 25196 23962
rect 24950 23908 24956 23910
rect 25012 23908 25036 23910
rect 25092 23908 25116 23910
rect 25172 23908 25196 23910
rect 25252 23908 25258 23910
rect 24950 23899 25258 23908
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 3350 23420 3658 23429
rect 3350 23418 3356 23420
rect 3412 23418 3436 23420
rect 3492 23418 3516 23420
rect 3572 23418 3596 23420
rect 3652 23418 3658 23420
rect 3412 23366 3414 23418
rect 3594 23366 3596 23418
rect 3350 23364 3356 23366
rect 3412 23364 3436 23366
rect 3492 23364 3516 23366
rect 3572 23364 3596 23366
rect 3652 23364 3658 23366
rect 3350 23355 3658 23364
rect 8150 23420 8458 23429
rect 8150 23418 8156 23420
rect 8212 23418 8236 23420
rect 8292 23418 8316 23420
rect 8372 23418 8396 23420
rect 8452 23418 8458 23420
rect 8212 23366 8214 23418
rect 8394 23366 8396 23418
rect 8150 23364 8156 23366
rect 8212 23364 8236 23366
rect 8292 23364 8316 23366
rect 8372 23364 8396 23366
rect 8452 23364 8458 23366
rect 8150 23355 8458 23364
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 17750 23420 18058 23429
rect 17750 23418 17756 23420
rect 17812 23418 17836 23420
rect 17892 23418 17916 23420
rect 17972 23418 17996 23420
rect 18052 23418 18058 23420
rect 17812 23366 17814 23418
rect 17994 23366 17996 23418
rect 17750 23364 17756 23366
rect 17812 23364 17836 23366
rect 17892 23364 17916 23366
rect 17972 23364 17996 23366
rect 18052 23364 18058 23366
rect 17750 23355 18058 23364
rect 22550 23420 22858 23429
rect 22550 23418 22556 23420
rect 22612 23418 22636 23420
rect 22692 23418 22716 23420
rect 22772 23418 22796 23420
rect 22852 23418 22858 23420
rect 22612 23366 22614 23418
rect 22794 23366 22796 23418
rect 22550 23364 22556 23366
rect 22612 23364 22636 23366
rect 22692 23364 22716 23366
rect 22772 23364 22796 23366
rect 22852 23364 22858 23366
rect 22550 23355 22858 23364
rect 5750 22876 6058 22885
rect 5750 22874 5756 22876
rect 5812 22874 5836 22876
rect 5892 22874 5916 22876
rect 5972 22874 5996 22876
rect 6052 22874 6058 22876
rect 5812 22822 5814 22874
rect 5994 22822 5996 22874
rect 5750 22820 5756 22822
rect 5812 22820 5836 22822
rect 5892 22820 5916 22822
rect 5972 22820 5996 22822
rect 6052 22820 6058 22822
rect 5750 22811 6058 22820
rect 10550 22876 10858 22885
rect 10550 22874 10556 22876
rect 10612 22874 10636 22876
rect 10692 22874 10716 22876
rect 10772 22874 10796 22876
rect 10852 22874 10858 22876
rect 10612 22822 10614 22874
rect 10794 22822 10796 22874
rect 10550 22820 10556 22822
rect 10612 22820 10636 22822
rect 10692 22820 10716 22822
rect 10772 22820 10796 22822
rect 10852 22820 10858 22822
rect 10550 22811 10858 22820
rect 15350 22876 15658 22885
rect 15350 22874 15356 22876
rect 15412 22874 15436 22876
rect 15492 22874 15516 22876
rect 15572 22874 15596 22876
rect 15652 22874 15658 22876
rect 15412 22822 15414 22874
rect 15594 22822 15596 22874
rect 15350 22820 15356 22822
rect 15412 22820 15436 22822
rect 15492 22820 15516 22822
rect 15572 22820 15596 22822
rect 15652 22820 15658 22822
rect 15350 22811 15658 22820
rect 20150 22876 20458 22885
rect 20150 22874 20156 22876
rect 20212 22874 20236 22876
rect 20292 22874 20316 22876
rect 20372 22874 20396 22876
rect 20452 22874 20458 22876
rect 20212 22822 20214 22874
rect 20394 22822 20396 22874
rect 20150 22820 20156 22822
rect 20212 22820 20236 22822
rect 20292 22820 20316 22822
rect 20372 22820 20396 22822
rect 20452 22820 20458 22822
rect 20150 22811 20458 22820
rect 24228 22778 24256 23666
rect 27350 23420 27658 23429
rect 27350 23418 27356 23420
rect 27412 23418 27436 23420
rect 27492 23418 27516 23420
rect 27572 23418 27596 23420
rect 27652 23418 27658 23420
rect 27412 23366 27414 23418
rect 27594 23366 27596 23418
rect 27350 23364 27356 23366
rect 27412 23364 27436 23366
rect 27492 23364 27516 23366
rect 27572 23364 27596 23366
rect 27652 23364 27658 23366
rect 27350 23355 27658 23364
rect 24950 22876 25258 22885
rect 24950 22874 24956 22876
rect 25012 22874 25036 22876
rect 25092 22874 25116 22876
rect 25172 22874 25196 22876
rect 25252 22874 25258 22876
rect 25012 22822 25014 22874
rect 25194 22822 25196 22874
rect 24950 22820 24956 22822
rect 25012 22820 25036 22822
rect 25092 22820 25116 22822
rect 25172 22820 25196 22822
rect 25252 22820 25258 22822
rect 24950 22811 25258 22820
rect 24216 22772 24268 22778
rect 24216 22714 24268 22720
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 2780 21616 2832 21622
rect 2780 21558 2832 21564
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 1780 21010 1808 21422
rect 1768 21004 1820 21010
rect 1768 20946 1820 20952
rect 2044 20868 2096 20874
rect 2044 20810 2096 20816
rect 2056 20058 2084 20810
rect 2148 20602 2176 21422
rect 2792 20874 2820 21558
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 2792 18630 2820 20810
rect 3068 20602 3096 21626
rect 3160 21146 3188 22578
rect 3350 22332 3658 22341
rect 3350 22330 3356 22332
rect 3412 22330 3436 22332
rect 3492 22330 3516 22332
rect 3572 22330 3596 22332
rect 3652 22330 3658 22332
rect 3412 22278 3414 22330
rect 3594 22278 3596 22330
rect 3350 22276 3356 22278
rect 3412 22276 3436 22278
rect 3492 22276 3516 22278
rect 3572 22276 3596 22278
rect 3652 22276 3658 22278
rect 3350 22267 3658 22276
rect 8150 22332 8458 22341
rect 8150 22330 8156 22332
rect 8212 22330 8236 22332
rect 8292 22330 8316 22332
rect 8372 22330 8396 22332
rect 8452 22330 8458 22332
rect 8212 22278 8214 22330
rect 8394 22278 8396 22330
rect 8150 22276 8156 22278
rect 8212 22276 8236 22278
rect 8292 22276 8316 22278
rect 8372 22276 8396 22278
rect 8452 22276 8458 22278
rect 8150 22267 8458 22276
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 17750 22332 18058 22341
rect 17750 22330 17756 22332
rect 17812 22330 17836 22332
rect 17892 22330 17916 22332
rect 17972 22330 17996 22332
rect 18052 22330 18058 22332
rect 17812 22278 17814 22330
rect 17994 22278 17996 22330
rect 17750 22276 17756 22278
rect 17812 22276 17836 22278
rect 17892 22276 17916 22278
rect 17972 22276 17996 22278
rect 18052 22276 18058 22278
rect 17750 22267 18058 22276
rect 22550 22332 22858 22341
rect 22550 22330 22556 22332
rect 22612 22330 22636 22332
rect 22692 22330 22716 22332
rect 22772 22330 22796 22332
rect 22852 22330 22858 22332
rect 22612 22278 22614 22330
rect 22794 22278 22796 22330
rect 22550 22276 22556 22278
rect 22612 22276 22636 22278
rect 22692 22276 22716 22278
rect 22772 22276 22796 22278
rect 22852 22276 22858 22278
rect 22550 22267 22858 22276
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 5750 21788 6058 21797
rect 5750 21786 5756 21788
rect 5812 21786 5836 21788
rect 5892 21786 5916 21788
rect 5972 21786 5996 21788
rect 6052 21786 6058 21788
rect 5812 21734 5814 21786
rect 5994 21734 5996 21786
rect 5750 21732 5756 21734
rect 5812 21732 5836 21734
rect 5892 21732 5916 21734
rect 5972 21732 5996 21734
rect 6052 21732 6058 21734
rect 5750 21723 6058 21732
rect 10550 21788 10858 21797
rect 10550 21786 10556 21788
rect 10612 21786 10636 21788
rect 10692 21786 10716 21788
rect 10772 21786 10796 21788
rect 10852 21786 10858 21788
rect 10612 21734 10614 21786
rect 10794 21734 10796 21786
rect 10550 21732 10556 21734
rect 10612 21732 10636 21734
rect 10692 21732 10716 21734
rect 10772 21732 10796 21734
rect 10852 21732 10858 21734
rect 10550 21723 10858 21732
rect 15350 21788 15658 21797
rect 15350 21786 15356 21788
rect 15412 21786 15436 21788
rect 15492 21786 15516 21788
rect 15572 21786 15596 21788
rect 15652 21786 15658 21788
rect 15412 21734 15414 21786
rect 15594 21734 15596 21786
rect 15350 21732 15356 21734
rect 15412 21732 15436 21734
rect 15492 21732 15516 21734
rect 15572 21732 15596 21734
rect 15652 21732 15658 21734
rect 15350 21723 15658 21732
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 3350 21244 3658 21253
rect 3350 21242 3356 21244
rect 3412 21242 3436 21244
rect 3492 21242 3516 21244
rect 3572 21242 3596 21244
rect 3652 21242 3658 21244
rect 3412 21190 3414 21242
rect 3594 21190 3596 21242
rect 3350 21188 3356 21190
rect 3412 21188 3436 21190
rect 3492 21188 3516 21190
rect 3572 21188 3596 21190
rect 3652 21188 3658 21190
rect 3350 21179 3658 21188
rect 8150 21244 8458 21253
rect 8150 21242 8156 21244
rect 8212 21242 8236 21244
rect 8292 21242 8316 21244
rect 8372 21242 8396 21244
rect 8452 21242 8458 21244
rect 8212 21190 8214 21242
rect 8394 21190 8396 21242
rect 8150 21188 8156 21190
rect 8212 21188 8236 21190
rect 8292 21188 8316 21190
rect 8372 21188 8396 21190
rect 8452 21188 8458 21190
rect 8150 21179 8458 21188
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 17750 21244 18058 21253
rect 17750 21242 17756 21244
rect 17812 21242 17836 21244
rect 17892 21242 17916 21244
rect 17972 21242 17996 21244
rect 18052 21242 18058 21244
rect 17812 21190 17814 21242
rect 17994 21190 17996 21242
rect 17750 21188 17756 21190
rect 17812 21188 17836 21190
rect 17892 21188 17916 21190
rect 17972 21188 17996 21190
rect 18052 21188 18058 21190
rect 17750 21179 18058 21188
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3240 21004 3292 21010
rect 3240 20946 3292 20952
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2792 18358 2820 18566
rect 3160 18426 3188 20402
rect 3252 18766 3280 20946
rect 4908 20806 4936 20946
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 6736 20868 6788 20874
rect 6736 20810 6788 20816
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3350 20156 3658 20165
rect 3350 20154 3356 20156
rect 3412 20154 3436 20156
rect 3492 20154 3516 20156
rect 3572 20154 3596 20156
rect 3652 20154 3658 20156
rect 3412 20102 3414 20154
rect 3594 20102 3596 20154
rect 3350 20100 3356 20102
rect 3412 20100 3436 20102
rect 3492 20100 3516 20102
rect 3572 20100 3596 20102
rect 3652 20100 3658 20102
rect 3350 20091 3658 20100
rect 3350 19068 3658 19077
rect 3350 19066 3356 19068
rect 3412 19066 3436 19068
rect 3492 19066 3516 19068
rect 3572 19066 3596 19068
rect 3652 19066 3658 19068
rect 3412 19014 3414 19066
rect 3594 19014 3596 19066
rect 3350 19012 3356 19014
rect 3412 19012 3436 19014
rect 3492 19012 3516 19014
rect 3572 19012 3596 19014
rect 3652 19012 3658 19014
rect 3350 19003 3658 19012
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17202 1532 17478
rect 1582 17368 1638 17377
rect 2240 17338 2268 18226
rect 2792 17762 2820 18294
rect 3252 18086 3280 18702
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 2700 17734 2820 17762
rect 2884 17746 2912 18022
rect 3252 17746 3280 18022
rect 3350 17980 3658 17989
rect 3350 17978 3356 17980
rect 3412 17978 3436 17980
rect 3492 17978 3516 17980
rect 3572 17978 3596 17980
rect 3652 17978 3658 17980
rect 3412 17926 3414 17978
rect 3594 17926 3596 17978
rect 3350 17924 3356 17926
rect 3412 17924 3436 17926
rect 3492 17924 3516 17926
rect 3572 17924 3596 17926
rect 3652 17924 3658 17926
rect 3350 17915 3658 17924
rect 2872 17740 2924 17746
rect 2700 17610 2728 17734
rect 2872 17682 2924 17688
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 1582 17303 1584 17312
rect 1636 17303 1638 17312
rect 2228 17332 2280 17338
rect 1584 17274 1636 17280
rect 2228 17274 2280 17280
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2608 16114 2636 17138
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2608 15706 2636 16050
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2700 15434 2728 17546
rect 3252 15570 3280 17682
rect 3804 17134 3832 20198
rect 3896 19854 3924 20742
rect 4908 20398 4936 20742
rect 5750 20700 6058 20709
rect 5750 20698 5756 20700
rect 5812 20698 5836 20700
rect 5892 20698 5916 20700
rect 5972 20698 5996 20700
rect 6052 20698 6058 20700
rect 5812 20646 5814 20698
rect 5994 20646 5996 20698
rect 5750 20644 5756 20646
rect 5812 20644 5836 20646
rect 5892 20644 5916 20646
rect 5972 20644 5996 20646
rect 6052 20644 6058 20646
rect 5750 20635 6058 20644
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 5750 19612 6058 19621
rect 5750 19610 5756 19612
rect 5812 19610 5836 19612
rect 5892 19610 5916 19612
rect 5972 19610 5996 19612
rect 6052 19610 6058 19612
rect 5812 19558 5814 19610
rect 5994 19558 5996 19610
rect 5750 19556 5756 19558
rect 5812 19556 5836 19558
rect 5892 19556 5916 19558
rect 5972 19556 5996 19558
rect 6052 19556 6058 19558
rect 5750 19547 6058 19556
rect 6748 18970 6776 20810
rect 10550 20700 10858 20709
rect 10550 20698 10556 20700
rect 10612 20698 10636 20700
rect 10692 20698 10716 20700
rect 10772 20698 10796 20700
rect 10852 20698 10858 20700
rect 10612 20646 10614 20698
rect 10794 20646 10796 20698
rect 10550 20644 10556 20646
rect 10612 20644 10636 20646
rect 10692 20644 10716 20646
rect 10772 20644 10796 20646
rect 10852 20644 10858 20646
rect 10550 20635 10858 20644
rect 15350 20700 15658 20709
rect 15350 20698 15356 20700
rect 15412 20698 15436 20700
rect 15492 20698 15516 20700
rect 15572 20698 15596 20700
rect 15652 20698 15658 20700
rect 15412 20646 15414 20698
rect 15594 20646 15596 20698
rect 15350 20644 15356 20646
rect 15412 20644 15436 20646
rect 15492 20644 15516 20646
rect 15572 20644 15596 20646
rect 15652 20644 15658 20646
rect 15350 20635 15658 20644
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 8150 20156 8458 20165
rect 8150 20154 8156 20156
rect 8212 20154 8236 20156
rect 8292 20154 8316 20156
rect 8372 20154 8396 20156
rect 8452 20154 8458 20156
rect 8212 20102 8214 20154
rect 8394 20102 8396 20154
rect 8150 20100 8156 20102
rect 8212 20100 8236 20102
rect 8292 20100 8316 20102
rect 8372 20100 8396 20102
rect 8452 20100 8458 20102
rect 8150 20091 8458 20100
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 16776 19922 16804 20198
rect 16868 20058 16896 20878
rect 18248 20806 18276 21626
rect 19168 21554 19196 22034
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19444 21622 19472 21830
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19524 21616 19576 21622
rect 19524 21558 19576 21564
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18248 20534 18276 20742
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 19168 20466 19196 21490
rect 19536 21486 19564 21558
rect 19524 21480 19576 21486
rect 19352 21440 19524 21468
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 10550 19612 10858 19621
rect 10550 19610 10556 19612
rect 10612 19610 10636 19612
rect 10692 19610 10716 19612
rect 10772 19610 10796 19612
rect 10852 19610 10858 19612
rect 10612 19558 10614 19610
rect 10794 19558 10796 19610
rect 10550 19556 10556 19558
rect 10612 19556 10636 19558
rect 10692 19556 10716 19558
rect 10772 19556 10796 19558
rect 10852 19556 10858 19558
rect 10550 19547 10858 19556
rect 15350 19612 15658 19621
rect 15350 19610 15356 19612
rect 15412 19610 15436 19612
rect 15492 19610 15516 19612
rect 15572 19610 15596 19612
rect 15652 19610 15658 19612
rect 15412 19558 15414 19610
rect 15594 19558 15596 19610
rect 15350 19556 15356 19558
rect 15412 19556 15436 19558
rect 15492 19556 15516 19558
rect 15572 19556 15596 19558
rect 15652 19556 15658 19558
rect 15350 19547 15658 19556
rect 17144 19446 17172 20402
rect 17750 20156 18058 20165
rect 17750 20154 17756 20156
rect 17812 20154 17836 20156
rect 17892 20154 17916 20156
rect 17972 20154 17996 20156
rect 18052 20154 18058 20156
rect 17812 20102 17814 20154
rect 17994 20102 17996 20154
rect 17750 20100 17756 20102
rect 17812 20100 17836 20102
rect 17892 20100 17916 20102
rect 17972 20100 17996 20102
rect 18052 20100 18058 20102
rect 17750 20091 18058 20100
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 8150 19068 8458 19077
rect 8150 19066 8156 19068
rect 8212 19066 8236 19068
rect 8292 19066 8316 19068
rect 8372 19066 8396 19068
rect 8452 19066 8458 19068
rect 8212 19014 8214 19066
rect 8394 19014 8396 19066
rect 8150 19012 8156 19014
rect 8212 19012 8236 19014
rect 8292 19012 8316 19014
rect 8372 19012 8396 19014
rect 8452 19012 8458 19014
rect 8150 19003 8458 19012
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3350 16892 3658 16901
rect 3350 16890 3356 16892
rect 3412 16890 3436 16892
rect 3492 16890 3516 16892
rect 3572 16890 3596 16892
rect 3652 16890 3658 16892
rect 3412 16838 3414 16890
rect 3594 16838 3596 16890
rect 3350 16836 3356 16838
rect 3412 16836 3436 16838
rect 3492 16836 3516 16838
rect 3572 16836 3596 16838
rect 3652 16836 3658 16838
rect 3350 16827 3658 16836
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3350 15804 3658 15813
rect 3350 15802 3356 15804
rect 3412 15802 3436 15804
rect 3492 15802 3516 15804
rect 3572 15802 3596 15804
rect 3652 15802 3658 15804
rect 3412 15750 3414 15802
rect 3594 15750 3596 15802
rect 3350 15748 3356 15750
rect 3412 15748 3436 15750
rect 3492 15748 3516 15750
rect 3572 15748 3596 15750
rect 3652 15748 3658 15750
rect 3350 15739 3658 15748
rect 3712 15706 3740 15846
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 3148 15020 3200 15026
rect 3252 15008 3280 15506
rect 3988 15094 4016 18566
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4080 17678 4108 18362
rect 4436 18216 4488 18222
rect 4436 18158 4488 18164
rect 4448 17882 4476 18158
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 4344 17808 4396 17814
rect 4344 17750 4396 17756
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 4080 17270 4108 17614
rect 4356 17542 4384 17750
rect 5092 17678 5120 18022
rect 5276 17882 5304 18634
rect 5750 18524 6058 18533
rect 5750 18522 5756 18524
rect 5812 18522 5836 18524
rect 5892 18522 5916 18524
rect 5972 18522 5996 18524
rect 6052 18522 6058 18524
rect 5812 18470 5814 18522
rect 5994 18470 5996 18522
rect 5750 18468 5756 18470
rect 5812 18468 5836 18470
rect 5892 18468 5916 18470
rect 5972 18468 5996 18470
rect 6052 18468 6058 18470
rect 5750 18459 6058 18468
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 6748 17678 6776 18906
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18358 8340 18566
rect 10550 18524 10858 18533
rect 10550 18522 10556 18524
rect 10612 18522 10636 18524
rect 10692 18522 10716 18524
rect 10772 18522 10796 18524
rect 10852 18522 10858 18524
rect 10612 18470 10614 18522
rect 10794 18470 10796 18522
rect 10550 18468 10556 18470
rect 10612 18468 10636 18470
rect 10692 18468 10716 18470
rect 10772 18468 10796 18470
rect 10852 18468 10858 18470
rect 10550 18459 10858 18468
rect 15350 18524 15658 18533
rect 15350 18522 15356 18524
rect 15412 18522 15436 18524
rect 15492 18522 15516 18524
rect 15572 18522 15596 18524
rect 15652 18522 15658 18524
rect 15412 18470 15414 18522
rect 15594 18470 15596 18522
rect 15350 18468 15356 18470
rect 15412 18468 15436 18470
rect 15492 18468 15516 18470
rect 15572 18468 15596 18470
rect 15652 18468 15658 18470
rect 15350 18459 15658 18468
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5264 17672 5316 17678
rect 5724 17672 5776 17678
rect 5264 17614 5316 17620
rect 5552 17632 5724 17660
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 3200 14980 3280 15008
rect 3148 14962 3200 14968
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 12918 1808 13126
rect 1768 12912 1820 12918
rect 1768 12854 1820 12860
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1490 12472 1546 12481
rect 1490 12407 1492 12416
rect 1544 12407 1546 12416
rect 1492 12378 1544 12384
rect 1780 11694 1808 12718
rect 2424 12442 2452 13262
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2608 12170 2636 14758
rect 3350 14716 3658 14725
rect 3350 14714 3356 14716
rect 3412 14714 3436 14716
rect 3492 14714 3516 14716
rect 3572 14714 3596 14716
rect 3652 14714 3658 14716
rect 3412 14662 3414 14714
rect 3594 14662 3596 14714
rect 3350 14660 3356 14662
rect 3412 14660 3436 14662
rect 3492 14660 3516 14662
rect 3572 14660 3596 14662
rect 3652 14660 3658 14662
rect 3350 14651 3658 14660
rect 3896 14618 3924 14894
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 4080 14498 4108 17070
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4172 15706 4200 16050
rect 4356 15978 4384 17478
rect 4540 16998 4568 17614
rect 5276 17066 5304 17614
rect 5552 17066 5580 17632
rect 5724 17614 5776 17620
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 5750 17436 6058 17445
rect 5750 17434 5756 17436
rect 5812 17434 5836 17436
rect 5892 17434 5916 17436
rect 5972 17434 5996 17436
rect 6052 17434 6058 17436
rect 5812 17382 5814 17434
rect 5994 17382 5996 17434
rect 5750 17380 5756 17382
rect 5812 17380 5836 17382
rect 5892 17380 5916 17382
rect 5972 17380 5996 17382
rect 6052 17380 6058 17382
rect 5750 17371 6058 17380
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 3896 14470 4108 14498
rect 3350 13628 3658 13637
rect 3350 13626 3356 13628
rect 3412 13626 3436 13628
rect 3492 13626 3516 13628
rect 3572 13626 3596 13628
rect 3652 13626 3658 13628
rect 3412 13574 3414 13626
rect 3594 13574 3596 13626
rect 3350 13572 3356 13574
rect 3412 13572 3436 13574
rect 3492 13572 3516 13574
rect 3572 13572 3596 13574
rect 3652 13572 3658 13574
rect 3350 13563 3658 13572
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1676 7948 1728 7954
rect 1780 7936 1808 11630
rect 2976 11558 3004 13194
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 3160 12102 3188 12854
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3252 12238 3280 12582
rect 3350 12540 3658 12549
rect 3350 12538 3356 12540
rect 3412 12538 3436 12540
rect 3492 12538 3516 12540
rect 3572 12538 3596 12540
rect 3652 12538 3658 12540
rect 3412 12486 3414 12538
rect 3594 12486 3596 12538
rect 3350 12484 3356 12486
rect 3412 12484 3436 12486
rect 3492 12484 3516 12486
rect 3572 12484 3596 12486
rect 3652 12484 3658 12486
rect 3350 12475 3658 12484
rect 3896 12306 3924 14470
rect 4172 14414 4200 14758
rect 4356 14550 4384 15914
rect 5276 15910 5304 17002
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3988 12918 4016 13194
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 4356 12714 4384 14486
rect 5184 14414 5212 15846
rect 5276 15706 5304 15846
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5276 14346 5304 15642
rect 5644 15094 5672 16934
rect 5750 16348 6058 16357
rect 5750 16346 5756 16348
rect 5812 16346 5836 16348
rect 5892 16346 5916 16348
rect 5972 16346 5996 16348
rect 6052 16346 6058 16348
rect 5812 16294 5814 16346
rect 5994 16294 5996 16346
rect 5750 16292 5756 16294
rect 5812 16292 5836 16294
rect 5892 16292 5916 16294
rect 5972 16292 5996 16294
rect 6052 16292 6058 16294
rect 5750 16283 6058 16292
rect 5750 15260 6058 15269
rect 5750 15258 5756 15260
rect 5812 15258 5836 15260
rect 5892 15258 5916 15260
rect 5972 15258 5996 15260
rect 6052 15258 6058 15260
rect 5812 15206 5814 15258
rect 5994 15206 5996 15258
rect 5750 15204 5756 15206
rect 5812 15204 5836 15206
rect 5892 15204 5916 15206
rect 5972 15204 5996 15206
rect 6052 15204 6058 15206
rect 5750 15195 6058 15204
rect 5632 15088 5684 15094
rect 5632 15030 5684 15036
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5828 14346 5856 14962
rect 6288 14414 6316 17478
rect 7392 16454 7420 18294
rect 8312 18170 8340 18294
rect 8312 18142 8616 18170
rect 8150 17980 8458 17989
rect 8150 17978 8156 17980
rect 8212 17978 8236 17980
rect 8292 17978 8316 17980
rect 8372 17978 8396 17980
rect 8452 17978 8458 17980
rect 8212 17926 8214 17978
rect 8394 17926 8396 17978
rect 8150 17924 8156 17926
rect 8212 17924 8236 17926
rect 8292 17924 8316 17926
rect 8372 17924 8396 17926
rect 8452 17924 8458 17926
rect 8150 17915 8458 17924
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7484 17270 7512 17478
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7484 14958 7512 16050
rect 7576 15162 7604 17070
rect 7668 15978 7696 17614
rect 7748 17604 7800 17610
rect 7800 17564 7880 17592
rect 7748 17546 7800 17552
rect 7852 16454 7880 17564
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7944 16590 7972 17274
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 8036 16522 8064 17614
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8150 16892 8458 16901
rect 8150 16890 8156 16892
rect 8212 16890 8236 16892
rect 8292 16890 8316 16892
rect 8372 16890 8396 16892
rect 8452 16890 8458 16892
rect 8212 16838 8214 16890
rect 8394 16838 8396 16890
rect 8150 16836 8156 16838
rect 8212 16836 8236 16838
rect 8292 16836 8316 16838
rect 8372 16836 8396 16838
rect 8452 16836 8458 16838
rect 8150 16827 8458 16836
rect 8496 16658 8524 17546
rect 8588 17270 8616 18142
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9140 17610 9168 18022
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 10550 17436 10858 17445
rect 10550 17434 10556 17436
rect 10612 17434 10636 17436
rect 10692 17434 10716 17436
rect 10772 17434 10796 17436
rect 10852 17434 10858 17436
rect 10612 17382 10614 17434
rect 10794 17382 10796 17434
rect 10550 17380 10556 17382
rect 10612 17380 10636 17382
rect 10692 17380 10716 17382
rect 10772 17380 10796 17382
rect 10852 17380 10858 17382
rect 10550 17371 10858 17380
rect 15350 17436 15658 17445
rect 15350 17434 15356 17436
rect 15412 17434 15436 17436
rect 15492 17434 15516 17436
rect 15572 17434 15596 17436
rect 15652 17434 15658 17436
rect 15412 17382 15414 17434
rect 15594 17382 15596 17434
rect 15350 17380 15356 17382
rect 15412 17380 15436 17382
rect 15492 17380 15516 17382
rect 15572 17380 15596 17382
rect 15652 17380 15658 17382
rect 15350 17371 15658 17380
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 7840 16448 7892 16454
rect 7760 16408 7840 16436
rect 7760 16250 7788 16408
rect 7840 16390 7892 16396
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 8036 16182 8064 16458
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 8220 16046 8248 16526
rect 8496 16182 8524 16594
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7576 15026 7604 15098
rect 7852 15094 7880 15846
rect 8150 15804 8458 15813
rect 8150 15802 8156 15804
rect 8212 15802 8236 15804
rect 8292 15802 8316 15804
rect 8372 15802 8396 15804
rect 8452 15802 8458 15804
rect 8212 15750 8214 15802
rect 8394 15750 8396 15802
rect 8150 15748 8156 15750
rect 8212 15748 8236 15750
rect 8292 15748 8316 15750
rect 8372 15748 8396 15750
rect 8452 15748 8458 15750
rect 8150 15739 8458 15748
rect 8588 15706 8616 17206
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 9140 15910 9168 16458
rect 9324 16114 9352 16934
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16182 9720 16526
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8588 15094 8616 15642
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 9140 14958 9168 15846
rect 9784 15366 9812 16934
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9968 16046 9996 16458
rect 10060 16114 10088 17070
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 10428 15892 10456 16526
rect 10888 16522 10916 16934
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12072 16584 12124 16590
rect 11992 16532 12072 16538
rect 11992 16526 12124 16532
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 11992 16510 12112 16526
rect 10550 16348 10858 16357
rect 10550 16346 10556 16348
rect 10612 16346 10636 16348
rect 10692 16346 10716 16348
rect 10772 16346 10796 16348
rect 10852 16346 10858 16348
rect 10612 16294 10614 16346
rect 10794 16294 10796 16346
rect 10550 16292 10556 16294
rect 10612 16292 10636 16294
rect 10692 16292 10716 16294
rect 10772 16292 10796 16294
rect 10852 16292 10858 16294
rect 10550 16283 10858 16292
rect 11992 16182 12020 16510
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 10600 15904 10652 15910
rect 10428 15864 10600 15892
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 11072 15502 11100 15982
rect 11244 15972 11296 15978
rect 11244 15914 11296 15920
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 4816 12918 4844 14214
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4816 12646 4844 12854
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3896 12102 3924 12242
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3712 11830 3740 12038
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 8634 3004 11494
rect 3350 11452 3658 11461
rect 3350 11450 3356 11452
rect 3412 11450 3436 11452
rect 3492 11450 3516 11452
rect 3572 11450 3596 11452
rect 3652 11450 3658 11452
rect 3412 11398 3414 11450
rect 3594 11398 3596 11450
rect 3350 11396 3356 11398
rect 3412 11396 3436 11398
rect 3492 11396 3516 11398
rect 3572 11396 3596 11398
rect 3652 11396 3658 11398
rect 3350 11387 3658 11396
rect 3350 10364 3658 10373
rect 3350 10362 3356 10364
rect 3412 10362 3436 10364
rect 3492 10362 3516 10364
rect 3572 10362 3596 10364
rect 3652 10362 3658 10364
rect 3412 10310 3414 10362
rect 3594 10310 3596 10362
rect 3350 10308 3356 10310
rect 3412 10308 3436 10310
rect 3492 10308 3516 10310
rect 3572 10308 3596 10310
rect 3652 10308 3658 10310
rect 3350 10299 3658 10308
rect 3350 9276 3658 9285
rect 3350 9274 3356 9276
rect 3412 9274 3436 9276
rect 3492 9274 3516 9276
rect 3572 9274 3596 9276
rect 3652 9274 3658 9276
rect 3412 9222 3414 9274
rect 3594 9222 3596 9274
rect 3350 9220 3356 9222
rect 3412 9220 3436 9222
rect 3492 9220 3516 9222
rect 3572 9220 3596 9222
rect 3652 9220 3658 9222
rect 3350 9211 3658 9220
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 7954 1992 8230
rect 1728 7908 1808 7936
rect 1952 7948 2004 7954
rect 1676 7890 1728 7896
rect 1952 7890 2004 7896
rect 1582 7576 1638 7585
rect 1582 7511 1584 7520
rect 1636 7511 1638 7520
rect 1584 7482 1636 7488
rect 1688 3602 1716 7890
rect 3160 4486 3188 8366
rect 3252 8072 3280 8434
rect 3350 8188 3658 8197
rect 3350 8186 3356 8188
rect 3412 8186 3436 8188
rect 3492 8186 3516 8188
rect 3572 8186 3596 8188
rect 3652 8186 3658 8188
rect 3412 8134 3414 8186
rect 3594 8134 3596 8186
rect 3350 8132 3356 8134
rect 3412 8132 3436 8134
rect 3492 8132 3516 8134
rect 3572 8132 3596 8134
rect 3652 8132 3658 8134
rect 3350 8123 3658 8132
rect 3252 8044 3464 8072
rect 3436 7750 3464 8044
rect 3712 7818 3740 11766
rect 3896 8430 3924 12038
rect 3988 11830 4016 12582
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 4816 11694 4844 12582
rect 5000 11898 5028 13262
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5092 12850 5120 13126
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4264 10606 4292 11086
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4540 10810 4568 10950
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4264 10062 4292 10542
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4540 9926 4568 10746
rect 4632 10674 4660 11086
rect 5552 10674 5580 14214
rect 5750 14172 6058 14181
rect 5750 14170 5756 14172
rect 5812 14170 5836 14172
rect 5892 14170 5916 14172
rect 5972 14170 5996 14172
rect 6052 14170 6058 14172
rect 5812 14118 5814 14170
rect 5994 14118 5996 14170
rect 5750 14116 5756 14118
rect 5812 14116 5836 14118
rect 5892 14116 5916 14118
rect 5972 14116 5996 14118
rect 6052 14116 6058 14118
rect 5750 14107 6058 14116
rect 6564 14006 6592 14758
rect 8150 14716 8458 14725
rect 8150 14714 8156 14716
rect 8212 14714 8236 14716
rect 8292 14714 8316 14716
rect 8372 14714 8396 14716
rect 8452 14714 8458 14716
rect 8212 14662 8214 14714
rect 8394 14662 8396 14714
rect 8150 14660 8156 14662
rect 8212 14660 8236 14662
rect 8292 14660 8316 14662
rect 8372 14660 8396 14662
rect 8452 14660 8458 14662
rect 8150 14651 8458 14660
rect 8496 14482 8524 14758
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 5750 13084 6058 13093
rect 5750 13082 5756 13084
rect 5812 13082 5836 13084
rect 5892 13082 5916 13084
rect 5972 13082 5996 13084
rect 6052 13082 6058 13084
rect 5812 13030 5814 13082
rect 5994 13030 5996 13082
rect 5750 13028 5756 13030
rect 5812 13028 5836 13030
rect 5892 13028 5916 13030
rect 5972 13028 5996 13030
rect 6052 13028 6058 13030
rect 5750 13019 6058 13028
rect 6656 12918 6684 14282
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6748 12782 6776 13738
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12238 6408 12582
rect 6748 12374 6776 12718
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 5750 11996 6058 12005
rect 5750 11994 5756 11996
rect 5812 11994 5836 11996
rect 5892 11994 5916 11996
rect 5972 11994 5996 11996
rect 6052 11994 6058 11996
rect 5812 11942 5814 11994
rect 5994 11942 5996 11994
rect 5750 11940 5756 11942
rect 5812 11940 5836 11942
rect 5892 11940 5916 11942
rect 5972 11940 5996 11942
rect 6052 11940 6058 11942
rect 5750 11931 6058 11940
rect 6380 11762 6408 12174
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 5750 10908 6058 10917
rect 5750 10906 5756 10908
rect 5812 10906 5836 10908
rect 5892 10906 5916 10908
rect 5972 10906 5996 10908
rect 6052 10906 6058 10908
rect 5812 10854 5814 10906
rect 5994 10854 5996 10906
rect 5750 10852 5756 10854
rect 5812 10852 5836 10854
rect 5892 10852 5916 10854
rect 5972 10852 5996 10854
rect 6052 10852 6058 10854
rect 5750 10843 6058 10852
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 4632 10198 4660 10610
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 9722 4568 9862
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4264 9042 4292 9454
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4540 8838 4568 9658
rect 4632 9586 4660 10134
rect 5000 10130 5028 10542
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 5000 9994 5028 10066
rect 5552 10062 5580 10610
rect 6748 10198 6776 12310
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6840 10062 6868 12038
rect 7024 11150 7052 12038
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4632 9110 4660 9522
rect 5000 9518 5028 9930
rect 5750 9820 6058 9829
rect 5750 9818 5756 9820
rect 5812 9818 5836 9820
rect 5892 9818 5916 9820
rect 5972 9818 5996 9820
rect 6052 9818 6058 9820
rect 5812 9766 5814 9818
rect 5994 9766 5996 9818
rect 5750 9764 5756 9766
rect 5812 9764 5836 9766
rect 5892 9764 5916 9766
rect 5972 9764 5996 9766
rect 6052 9764 6058 9766
rect 5750 9755 6058 9764
rect 6932 9654 6960 9930
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 7116 8974 7144 14282
rect 8150 13628 8458 13637
rect 8150 13626 8156 13628
rect 8212 13626 8236 13628
rect 8292 13626 8316 13628
rect 8372 13626 8396 13628
rect 8452 13626 8458 13628
rect 8212 13574 8214 13626
rect 8394 13574 8396 13626
rect 8150 13572 8156 13574
rect 8212 13572 8236 13574
rect 8292 13572 8316 13574
rect 8372 13572 8396 13574
rect 8452 13572 8458 13574
rect 8150 13563 8458 13572
rect 8496 12986 8524 14418
rect 9784 13530 9812 15302
rect 10550 15260 10858 15269
rect 10550 15258 10556 15260
rect 10612 15258 10636 15260
rect 10692 15258 10716 15260
rect 10772 15258 10796 15260
rect 10852 15258 10858 15260
rect 10612 15206 10614 15258
rect 10794 15206 10796 15258
rect 10550 15204 10556 15206
rect 10612 15204 10636 15206
rect 10692 15204 10716 15206
rect 10772 15204 10796 15206
rect 10852 15204 10858 15206
rect 10550 15195 10858 15204
rect 11164 15094 11192 15642
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 10550 14172 10858 14181
rect 10550 14170 10556 14172
rect 10612 14170 10636 14172
rect 10692 14170 10716 14172
rect 10772 14170 10796 14172
rect 10852 14170 10858 14172
rect 10612 14118 10614 14170
rect 10794 14118 10796 14170
rect 10550 14116 10556 14118
rect 10612 14116 10636 14118
rect 10692 14116 10716 14118
rect 10772 14116 10796 14118
rect 10852 14116 10858 14118
rect 10550 14107 10858 14116
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8588 12850 8616 13330
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 7392 12306 7420 12582
rect 8150 12540 8458 12549
rect 8150 12538 8156 12540
rect 8212 12538 8236 12540
rect 8292 12538 8316 12540
rect 8372 12538 8396 12540
rect 8452 12538 8458 12540
rect 8212 12486 8214 12538
rect 8394 12486 8396 12538
rect 8150 12484 8156 12486
rect 8212 12484 8236 12486
rect 8292 12484 8316 12486
rect 8372 12484 8396 12486
rect 8452 12484 8458 12486
rect 8150 12475 8458 12484
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11218 7604 11494
rect 8150 11452 8458 11461
rect 8150 11450 8156 11452
rect 8212 11450 8236 11452
rect 8292 11450 8316 11452
rect 8372 11450 8396 11452
rect 8452 11450 8458 11452
rect 8212 11398 8214 11450
rect 8394 11398 8396 11450
rect 8150 11396 8156 11398
rect 8212 11396 8236 11398
rect 8292 11396 8316 11398
rect 8372 11396 8396 11398
rect 8452 11396 8458 11398
rect 8150 11387 8458 11396
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 8680 11150 8708 12582
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8150 10364 8458 10373
rect 8150 10362 8156 10364
rect 8212 10362 8236 10364
rect 8292 10362 8316 10364
rect 8372 10362 8396 10364
rect 8452 10362 8458 10364
rect 8212 10310 8214 10362
rect 8394 10310 8396 10362
rect 8150 10308 8156 10310
rect 8212 10308 8236 10310
rect 8292 10308 8316 10310
rect 8372 10308 8396 10310
rect 8452 10308 8458 10310
rect 8150 10299 8458 10308
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9586 8340 9862
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8150 9276 8458 9285
rect 8150 9274 8156 9276
rect 8212 9274 8236 9276
rect 8292 9274 8316 9276
rect 8372 9274 8396 9276
rect 8452 9274 8458 9276
rect 8212 9222 8214 9274
rect 8394 9222 8396 9274
rect 8150 9220 8156 9222
rect 8212 9220 8236 9222
rect 8292 9220 8316 9222
rect 8372 9220 8396 9222
rect 8452 9220 8458 9222
rect 8150 9211 8458 9220
rect 8496 8974 8524 9522
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 5460 8072 5488 8774
rect 5750 8732 6058 8741
rect 5750 8730 5756 8732
rect 5812 8730 5836 8732
rect 5892 8730 5916 8732
rect 5972 8730 5996 8732
rect 6052 8730 6058 8732
rect 5812 8678 5814 8730
rect 5994 8678 5996 8730
rect 5750 8676 5756 8678
rect 5812 8676 5836 8678
rect 5892 8676 5916 8678
rect 5972 8676 5996 8678
rect 6052 8676 6058 8678
rect 5750 8667 6058 8676
rect 7116 8498 7144 8910
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8128 8634 8156 8842
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8588 8498 8616 9386
rect 8772 9382 8800 11630
rect 9048 11626 9076 13262
rect 9784 13258 9812 13466
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9600 12986 9628 13194
rect 10550 13084 10858 13093
rect 10550 13082 10556 13084
rect 10612 13082 10636 13084
rect 10692 13082 10716 13084
rect 10772 13082 10796 13084
rect 10852 13082 10858 13084
rect 10612 13030 10614 13082
rect 10794 13030 10796 13082
rect 10550 13028 10556 13030
rect 10612 13028 10636 13030
rect 10692 13028 10716 13030
rect 10772 13028 10796 13030
rect 10852 13028 10858 13030
rect 10550 13019 10858 13028
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 10980 12850 11008 13466
rect 11164 13190 11192 15030
rect 11256 15026 11284 15914
rect 11624 15706 11652 15982
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11624 15162 11652 15642
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11256 13326 11284 14962
rect 11900 14890 11928 15982
rect 11992 15026 12020 16118
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 12084 15094 12112 15370
rect 12176 15162 12204 16390
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 12268 14482 12296 16594
rect 12360 16182 12388 16934
rect 12820 16658 12848 16934
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 14568 16794 14596 17070
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 15120 16658 15148 17206
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 12820 16250 12848 16594
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 14844 16114 14872 16526
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12360 14822 12388 15982
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15026 12480 15846
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 15120 15570 15148 16594
rect 15212 16522 15240 17002
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15350 16348 15658 16357
rect 15350 16346 15356 16348
rect 15412 16346 15436 16348
rect 15492 16346 15516 16348
rect 15572 16346 15596 16348
rect 15652 16346 15658 16348
rect 15412 16294 15414 16346
rect 15594 16294 15596 16346
rect 15350 16292 15356 16294
rect 15412 16292 15436 16294
rect 15492 16292 15516 16294
rect 15572 16292 15596 16294
rect 15652 16292 15658 16294
rect 15350 16283 15658 16292
rect 15764 16182 15792 17070
rect 15856 16658 15884 17478
rect 16500 16794 16528 17614
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 16592 16590 16620 19382
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17236 17270 17264 19314
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16960 16658 16988 17070
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11256 12986 11284 13262
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 9692 12646 9720 12786
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 9048 10810 9076 11562
rect 9600 11218 9628 12242
rect 9876 12170 9904 12718
rect 11348 12714 11376 12922
rect 12268 12850 12296 13126
rect 12452 12986 12480 13806
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13462 12572 13670
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13556 13530 13584 13874
rect 14108 13530 14136 13874
rect 15120 13802 15148 14282
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12544 12918 12572 13398
rect 14200 13326 14228 13738
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14844 13530 14872 13670
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 15212 13394 15240 16050
rect 15764 15434 15792 16118
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15350 15260 15658 15269
rect 15350 15258 15356 15260
rect 15412 15258 15436 15260
rect 15492 15258 15516 15260
rect 15572 15258 15596 15260
rect 15652 15258 15658 15260
rect 15412 15206 15414 15258
rect 15594 15206 15596 15258
rect 15350 15204 15356 15206
rect 15412 15204 15436 15206
rect 15492 15204 15516 15206
rect 15572 15204 15596 15206
rect 15652 15204 15658 15206
rect 15350 15195 15658 15204
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15350 14172 15658 14181
rect 15350 14170 15356 14172
rect 15412 14170 15436 14172
rect 15492 14170 15516 14172
rect 15572 14170 15596 14172
rect 15652 14170 15658 14172
rect 15412 14118 15414 14170
rect 15594 14118 15596 14170
rect 15350 14116 15356 14118
rect 15412 14116 15436 14118
rect 15492 14116 15516 14118
rect 15572 14116 15596 14118
rect 15652 14116 15658 14118
rect 15350 14107 15658 14116
rect 15764 14074 15792 14758
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15764 13954 15792 14010
rect 15384 13932 15436 13938
rect 15764 13926 15884 13954
rect 15384 13874 15436 13880
rect 15396 13530 15424 13874
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10428 12434 10456 12582
rect 10244 12406 10456 12434
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9508 9518 9536 10678
rect 9600 9586 9628 11154
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9722 9720 9862
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8772 8498 8800 9318
rect 9140 9042 9168 9386
rect 9692 9382 9720 9658
rect 9784 9586 9812 10134
rect 9968 10062 9996 10542
rect 10152 10470 10180 12038
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9968 9586 9996 9998
rect 10152 9926 10180 10406
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 5540 8084 5592 8090
rect 5460 8044 5540 8072
rect 5540 8026 5592 8032
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3436 7410 3464 7686
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3350 7100 3658 7109
rect 3350 7098 3356 7100
rect 3412 7098 3436 7100
rect 3492 7098 3516 7100
rect 3572 7098 3596 7100
rect 3652 7098 3658 7100
rect 3412 7046 3414 7098
rect 3594 7046 3596 7098
rect 3350 7044 3356 7046
rect 3412 7044 3436 7046
rect 3492 7044 3516 7046
rect 3572 7044 3596 7046
rect 3652 7044 3658 7046
rect 3350 7035 3658 7044
rect 3350 6012 3658 6021
rect 3350 6010 3356 6012
rect 3412 6010 3436 6012
rect 3492 6010 3516 6012
rect 3572 6010 3596 6012
rect 3652 6010 3658 6012
rect 3412 5958 3414 6010
rect 3594 5958 3596 6010
rect 3350 5956 3356 5958
rect 3412 5956 3436 5958
rect 3492 5956 3516 5958
rect 3572 5956 3596 5958
rect 3652 5956 3658 5958
rect 3350 5947 3658 5956
rect 3350 4924 3658 4933
rect 3350 4922 3356 4924
rect 3412 4922 3436 4924
rect 3492 4922 3516 4924
rect 3572 4922 3596 4924
rect 3652 4922 3658 4924
rect 3412 4870 3414 4922
rect 3594 4870 3596 4922
rect 3350 4868 3356 4870
rect 3412 4868 3436 4870
rect 3492 4868 3516 4870
rect 3572 4868 3596 4870
rect 3652 4868 3658 4870
rect 3350 4859 3658 4868
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 4078 3188 4422
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1780 3058 1808 3334
rect 2240 3194 2268 3402
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2516 3058 2544 3878
rect 2976 3738 3004 4014
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3350 3836 3658 3845
rect 3350 3834 3356 3836
rect 3412 3834 3436 3836
rect 3492 3834 3516 3836
rect 3572 3834 3596 3836
rect 3652 3834 3658 3836
rect 3412 3782 3414 3834
rect 3594 3782 3596 3834
rect 3350 3780 3356 3782
rect 3412 3780 3436 3782
rect 3492 3780 3516 3782
rect 3572 3780 3596 3782
rect 3652 3780 3658 3782
rect 3350 3771 3658 3780
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2976 3398 3004 3674
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 3068 3194 3096 3470
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3712 3058 3740 3878
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2689 1624 2790
rect 3350 2748 3658 2757
rect 3350 2746 3356 2748
rect 3412 2746 3436 2748
rect 3492 2746 3516 2748
rect 3572 2746 3596 2748
rect 3652 2746 3658 2748
rect 3412 2694 3414 2746
rect 3594 2694 3596 2746
rect 3350 2692 3356 2694
rect 3412 2692 3436 2694
rect 3492 2692 3516 2694
rect 3572 2692 3596 2694
rect 3652 2692 3658 2694
rect 1582 2680 1638 2689
rect 3350 2683 3658 2692
rect 1582 2615 1638 2624
rect 3804 800 3832 3538
rect 3896 3534 3924 7686
rect 5552 7546 5580 8026
rect 7116 7886 7144 8230
rect 7300 7954 7328 8366
rect 8150 8188 8458 8197
rect 8150 8186 8156 8188
rect 8212 8186 8236 8188
rect 8292 8186 8316 8188
rect 8372 8186 8396 8188
rect 8452 8186 8458 8188
rect 8212 8134 8214 8186
rect 8394 8134 8396 8186
rect 8150 8132 8156 8134
rect 8212 8132 8236 8134
rect 8292 8132 8316 8134
rect 8372 8132 8396 8134
rect 8452 8132 8458 8134
rect 8150 8123 8458 8132
rect 8588 8090 8616 8434
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 5750 7644 6058 7653
rect 5750 7642 5756 7644
rect 5812 7642 5836 7644
rect 5892 7642 5916 7644
rect 5972 7642 5996 7644
rect 6052 7642 6058 7644
rect 5812 7590 5814 7642
rect 5994 7590 5996 7642
rect 5750 7588 5756 7590
rect 5812 7588 5836 7590
rect 5892 7588 5916 7590
rect 5972 7588 5996 7590
rect 6052 7588 6058 7590
rect 5750 7579 6058 7588
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5552 7002 5580 7482
rect 7300 7410 7328 7890
rect 9048 7886 9076 8230
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5552 6458 5580 6938
rect 7300 6866 7328 7346
rect 7668 7274 7696 7822
rect 9692 7546 9720 9318
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 5750 6556 6058 6565
rect 5750 6554 5756 6556
rect 5812 6554 5836 6556
rect 5892 6554 5916 6556
rect 5972 6554 5996 6556
rect 6052 6554 6058 6556
rect 5812 6502 5814 6554
rect 5994 6502 5996 6554
rect 5750 6500 5756 6502
rect 5812 6500 5836 6502
rect 5892 6500 5916 6502
rect 5972 6500 5996 6502
rect 6052 6500 6058 6502
rect 5750 6491 6058 6500
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6656 5574 6684 6394
rect 7300 6322 7328 6802
rect 7668 6798 7696 7210
rect 8150 7100 8458 7109
rect 8150 7098 8156 7100
rect 8212 7098 8236 7100
rect 8292 7098 8316 7100
rect 8372 7098 8396 7100
rect 8452 7098 8458 7100
rect 8212 7046 8214 7098
rect 8394 7046 8396 7098
rect 8150 7044 8156 7046
rect 8212 7044 8236 7046
rect 8292 7044 8316 7046
rect 8372 7044 8396 7046
rect 8452 7044 8458 7046
rect 8150 7035 8458 7044
rect 9692 7002 9720 7482
rect 9876 7342 9904 7754
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9876 6866 9904 7278
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6322 8248 6734
rect 9876 6322 9904 6802
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7300 5846 7328 6122
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7668 5778 7696 6258
rect 8150 6012 8458 6021
rect 8150 6010 8156 6012
rect 8212 6010 8236 6012
rect 8292 6010 8316 6012
rect 8372 6010 8396 6012
rect 8452 6010 8458 6012
rect 8212 5958 8214 6010
rect 8394 5958 8396 6010
rect 8150 5956 8156 5958
rect 8212 5956 8236 5958
rect 8292 5956 8316 5958
rect 8372 5956 8396 5958
rect 8452 5956 8458 5958
rect 8150 5947 8458 5956
rect 9876 5778 9904 6258
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 5750 5468 6058 5477
rect 5750 5466 5756 5468
rect 5812 5466 5836 5468
rect 5892 5466 5916 5468
rect 5972 5466 5996 5468
rect 6052 5466 6058 5468
rect 5812 5414 5814 5466
rect 5994 5414 5996 5466
rect 5750 5412 5756 5414
rect 5812 5412 5836 5414
rect 5892 5412 5916 5414
rect 5972 5412 5996 5414
rect 6052 5412 6058 5414
rect 5750 5403 6058 5412
rect 8150 4924 8458 4933
rect 8150 4922 8156 4924
rect 8212 4922 8236 4924
rect 8292 4922 8316 4924
rect 8372 4922 8396 4924
rect 8452 4922 8458 4924
rect 8212 4870 8214 4922
rect 8394 4870 8396 4922
rect 8150 4868 8156 4870
rect 8212 4868 8236 4870
rect 8292 4868 8316 4870
rect 8372 4868 8396 4870
rect 8452 4868 8458 4870
rect 8150 4859 8458 4868
rect 5750 4380 6058 4389
rect 5750 4378 5756 4380
rect 5812 4378 5836 4380
rect 5892 4378 5916 4380
rect 5972 4378 5996 4380
rect 6052 4378 6058 4380
rect 5812 4326 5814 4378
rect 5994 4326 5996 4378
rect 5750 4324 5756 4326
rect 5812 4324 5836 4326
rect 5892 4324 5916 4326
rect 5972 4324 5996 4326
rect 6052 4324 6058 4326
rect 5750 4315 6058 4324
rect 10244 4282 10272 12406
rect 12268 12238 12296 12786
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12360 12374 12388 12582
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 10550 11996 10858 12005
rect 10550 11994 10556 11996
rect 10612 11994 10636 11996
rect 10692 11994 10716 11996
rect 10772 11994 10796 11996
rect 10852 11994 10858 11996
rect 10612 11942 10614 11994
rect 10794 11942 10796 11994
rect 10550 11940 10556 11942
rect 10612 11940 10636 11942
rect 10692 11940 10716 11942
rect 10772 11940 10796 11942
rect 10852 11940 10858 11942
rect 10550 11931 10858 11940
rect 10980 11354 11008 12106
rect 12820 12102 12848 13126
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12646 13860 12786
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11354 12848 12038
rect 12912 11762 12940 12174
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11830 13584 12038
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10428 10674 10456 10950
rect 10550 10908 10858 10917
rect 10550 10906 10556 10908
rect 10612 10906 10636 10908
rect 10692 10906 10716 10908
rect 10772 10906 10796 10908
rect 10852 10906 10858 10908
rect 10612 10854 10614 10906
rect 10794 10854 10796 10906
rect 10550 10852 10556 10854
rect 10612 10852 10636 10854
rect 10692 10852 10716 10854
rect 10772 10852 10796 10854
rect 10852 10852 10858 10854
rect 10550 10843 10858 10852
rect 10980 10742 11008 11290
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 11072 10674 11100 11154
rect 12820 10810 12848 11290
rect 13372 11218 13400 11494
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12820 10690 12848 10746
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12728 10662 12848 10690
rect 10336 10062 10364 10610
rect 10428 10198 10456 10610
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9722 10364 9998
rect 10550 9820 10858 9829
rect 10550 9818 10556 9820
rect 10612 9818 10636 9820
rect 10692 9818 10716 9820
rect 10772 9818 10796 9820
rect 10852 9818 10858 9820
rect 10612 9766 10614 9818
rect 10794 9766 10796 9818
rect 10550 9764 10556 9766
rect 10612 9764 10636 9766
rect 10692 9764 10716 9766
rect 10772 9764 10796 9766
rect 10852 9764 10858 9766
rect 10550 9755 10858 9764
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 11072 9586 11100 10610
rect 11992 9654 12020 10610
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 10062 12664 10474
rect 12728 10266 12756 10662
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12728 9722 12756 10202
rect 13188 10062 13216 10202
rect 13740 10062 13768 10202
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 12728 9518 12756 9658
rect 13096 9518 13124 9930
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 8974 10916 9318
rect 12268 9178 12296 9454
rect 12728 9178 12756 9454
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 10550 8732 10858 8741
rect 10550 8730 10556 8732
rect 10612 8730 10636 8732
rect 10692 8730 10716 8732
rect 10772 8730 10796 8732
rect 10852 8730 10858 8732
rect 10612 8678 10614 8730
rect 10794 8678 10796 8730
rect 10550 8676 10556 8678
rect 10612 8676 10636 8678
rect 10692 8676 10716 8678
rect 10772 8676 10796 8678
rect 10852 8676 10858 8678
rect 10550 8667 10858 8676
rect 12728 8498 12756 8842
rect 13096 8634 13124 9114
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 13096 8430 13124 8570
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12636 8090 12664 8366
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 13740 7954 13768 8434
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 10550 7644 10858 7653
rect 10550 7642 10556 7644
rect 10612 7642 10636 7644
rect 10692 7642 10716 7644
rect 10772 7642 10796 7644
rect 10852 7642 10858 7644
rect 10612 7590 10614 7642
rect 10794 7590 10796 7642
rect 10550 7588 10556 7590
rect 10612 7588 10636 7590
rect 10692 7588 10716 7590
rect 10772 7588 10796 7590
rect 10852 7588 10858 7590
rect 10550 7579 10858 7588
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10428 6798 10456 6938
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10550 6556 10858 6565
rect 10550 6554 10556 6556
rect 10612 6554 10636 6556
rect 10692 6554 10716 6556
rect 10772 6554 10796 6556
rect 10852 6554 10858 6556
rect 10612 6502 10614 6554
rect 10794 6502 10796 6554
rect 10550 6500 10556 6502
rect 10612 6500 10636 6502
rect 10692 6500 10716 6502
rect 10772 6500 10796 6502
rect 10852 6500 10858 6502
rect 10550 6491 10858 6500
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12636 5914 12664 6054
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10550 5468 10858 5477
rect 10550 5466 10556 5468
rect 10612 5466 10636 5468
rect 10692 5466 10716 5468
rect 10772 5466 10796 5468
rect 10852 5466 10858 5468
rect 10612 5414 10614 5466
rect 10794 5414 10796 5466
rect 10550 5412 10556 5414
rect 10612 5412 10636 5414
rect 10692 5412 10716 5414
rect 10772 5412 10796 5414
rect 10852 5412 10858 5414
rect 10550 5403 10858 5412
rect 10980 5234 11008 5714
rect 11716 5574 11744 5782
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11716 5370 11744 5510
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10612 4826 10640 5170
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10550 4380 10858 4389
rect 10550 4378 10556 4380
rect 10612 4378 10636 4380
rect 10692 4378 10716 4380
rect 10772 4378 10796 4380
rect 10852 4378 10858 4380
rect 10612 4326 10614 4378
rect 10794 4326 10796 4378
rect 10550 4324 10556 4326
rect 10612 4324 10636 4326
rect 10692 4324 10716 4326
rect 10772 4324 10796 4326
rect 10852 4324 10858 4326
rect 10550 4315 10858 4324
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 8150 3836 8458 3845
rect 8150 3834 8156 3836
rect 8212 3834 8236 3836
rect 8292 3834 8316 3836
rect 8372 3834 8396 3836
rect 8452 3834 8458 3836
rect 8212 3782 8214 3834
rect 8394 3782 8396 3834
rect 8150 3780 8156 3782
rect 8212 3780 8236 3782
rect 8292 3780 8316 3782
rect 8372 3780 8396 3782
rect 8452 3780 8458 3782
rect 8150 3771 8458 3780
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 5750 3292 6058 3301
rect 5750 3290 5756 3292
rect 5812 3290 5836 3292
rect 5892 3290 5916 3292
rect 5972 3290 5996 3292
rect 6052 3290 6058 3292
rect 5812 3238 5814 3290
rect 5994 3238 5996 3290
rect 5750 3236 5756 3238
rect 5812 3236 5836 3238
rect 5892 3236 5916 3238
rect 5972 3236 5996 3238
rect 6052 3236 6058 3238
rect 5750 3227 6058 3236
rect 10550 3292 10858 3301
rect 10550 3290 10556 3292
rect 10612 3290 10636 3292
rect 10692 3290 10716 3292
rect 10772 3290 10796 3292
rect 10852 3290 10858 3292
rect 10612 3238 10614 3290
rect 10794 3238 10796 3290
rect 10550 3236 10556 3238
rect 10612 3236 10636 3238
rect 10692 3236 10716 3238
rect 10772 3236 10796 3238
rect 10852 3236 10858 3238
rect 10550 3227 10858 3236
rect 8150 2748 8458 2757
rect 8150 2746 8156 2748
rect 8212 2746 8236 2748
rect 8292 2746 8316 2748
rect 8372 2746 8396 2748
rect 8452 2746 8458 2748
rect 8212 2694 8214 2746
rect 8394 2694 8396 2746
rect 8150 2692 8156 2694
rect 8212 2692 8236 2694
rect 8292 2692 8316 2694
rect 8372 2692 8396 2694
rect 8452 2692 8458 2694
rect 8150 2683 8458 2692
rect 11624 2650 11652 4150
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13832 3602 13860 12582
rect 15212 12442 15240 13126
rect 15350 13084 15658 13093
rect 15350 13082 15356 13084
rect 15412 13082 15436 13084
rect 15492 13082 15516 13084
rect 15572 13082 15596 13084
rect 15652 13082 15658 13084
rect 15412 13030 15414 13082
rect 15594 13030 15596 13082
rect 15350 13028 15356 13030
rect 15412 13028 15436 13030
rect 15492 13028 15516 13030
rect 15572 13028 15596 13030
rect 15652 13028 15658 13030
rect 15350 13019 15658 13028
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15350 11996 15658 12005
rect 15350 11994 15356 11996
rect 15412 11994 15436 11996
rect 15492 11994 15516 11996
rect 15572 11994 15596 11996
rect 15652 11994 15658 11996
rect 15412 11942 15414 11994
rect 15594 11942 15596 11994
rect 15350 11940 15356 11942
rect 15412 11940 15436 11942
rect 15492 11940 15516 11942
rect 15572 11940 15596 11942
rect 15652 11940 15658 11942
rect 15350 11931 15658 11940
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13924 10266 13952 11494
rect 15764 11014 15792 13806
rect 15856 13258 15884 13926
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15948 12782 15976 15302
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16224 13870 16252 14418
rect 16592 14346 16620 16526
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 14414 17264 14826
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 14006 16712 14214
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15350 10908 15658 10917
rect 15350 10906 15356 10908
rect 15412 10906 15436 10908
rect 15492 10906 15516 10908
rect 15572 10906 15596 10908
rect 15652 10906 15658 10908
rect 15412 10854 15414 10906
rect 15594 10854 15596 10906
rect 15350 10852 15356 10854
rect 15412 10852 15436 10854
rect 15492 10852 15516 10854
rect 15572 10852 15596 10854
rect 15652 10852 15658 10854
rect 15350 10843 15658 10852
rect 15764 10674 15792 10950
rect 16224 10810 16252 13806
rect 16684 13326 16712 13942
rect 16960 13394 16988 14282
rect 17420 14074 17448 19858
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17512 17678 17540 19654
rect 19352 19514 19380 21440
rect 19524 21422 19576 21428
rect 19536 21357 19564 21422
rect 19996 21146 20024 21966
rect 20150 21788 20458 21797
rect 20150 21786 20156 21788
rect 20212 21786 20236 21788
rect 20292 21786 20316 21788
rect 20372 21786 20396 21788
rect 20452 21786 20458 21788
rect 20212 21734 20214 21786
rect 20394 21734 20396 21786
rect 20150 21732 20156 21734
rect 20212 21732 20236 21734
rect 20292 21732 20316 21734
rect 20372 21732 20396 21734
rect 20452 21732 20458 21734
rect 20150 21723 20458 21732
rect 23492 21622 23520 22646
rect 24124 22432 24176 22438
rect 24124 22374 24176 22380
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 23664 22092 23716 22098
rect 23664 22034 23716 22040
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20456 21010 20484 21286
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19536 19514 19564 20742
rect 20150 20700 20458 20709
rect 20150 20698 20156 20700
rect 20212 20698 20236 20700
rect 20292 20698 20316 20700
rect 20372 20698 20396 20700
rect 20452 20698 20458 20700
rect 20212 20646 20214 20698
rect 20394 20646 20396 20698
rect 20150 20644 20156 20646
rect 20212 20644 20236 20646
rect 20292 20644 20316 20646
rect 20372 20644 20396 20646
rect 20452 20644 20458 20646
rect 20150 20635 20458 20644
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 17750 19068 18058 19077
rect 17750 19066 17756 19068
rect 17812 19066 17836 19068
rect 17892 19066 17916 19068
rect 17972 19066 17996 19068
rect 18052 19066 18058 19068
rect 17812 19014 17814 19066
rect 17994 19014 17996 19066
rect 17750 19012 17756 19014
rect 17812 19012 17836 19014
rect 17892 19012 17916 19014
rect 17972 19012 17996 19014
rect 18052 19012 18058 19014
rect 17750 19003 18058 19012
rect 18156 18970 18184 19246
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 17750 17980 18058 17989
rect 17750 17978 17756 17980
rect 17812 17978 17836 17980
rect 17892 17978 17916 17980
rect 17972 17978 17996 17980
rect 18052 17978 18058 17980
rect 17812 17926 17814 17978
rect 17994 17926 17996 17978
rect 17750 17924 17756 17926
rect 17812 17924 17836 17926
rect 17892 17924 17916 17926
rect 17972 17924 17996 17926
rect 18052 17924 18058 17926
rect 17750 17915 18058 17924
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17512 17270 17540 17614
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 17512 16658 17540 17206
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17604 16538 17632 16934
rect 17750 16892 18058 16901
rect 17750 16890 17756 16892
rect 17812 16890 17836 16892
rect 17892 16890 17916 16892
rect 17972 16890 17996 16892
rect 18052 16890 18058 16892
rect 17812 16838 17814 16890
rect 17994 16838 17996 16890
rect 17750 16836 17756 16838
rect 17812 16836 17836 16838
rect 17892 16836 17916 16838
rect 17972 16836 17996 16838
rect 18052 16836 18058 16838
rect 17750 16827 18058 16836
rect 17604 16522 17724 16538
rect 18156 16522 18184 17750
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18248 17202 18276 17614
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18800 16998 18828 18702
rect 19352 18358 19380 19450
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19536 17814 19564 19450
rect 19812 18290 19840 20402
rect 20732 19922 20760 20946
rect 22008 20936 22060 20942
rect 22008 20878 22060 20884
rect 22020 20602 22048 20878
rect 22388 20602 22416 21286
rect 22550 21244 22858 21253
rect 22550 21242 22556 21244
rect 22612 21242 22636 21244
rect 22692 21242 22716 21244
rect 22772 21242 22796 21244
rect 22852 21242 22858 21244
rect 22612 21190 22614 21242
rect 22794 21190 22796 21242
rect 22550 21188 22556 21190
rect 22612 21188 22636 21190
rect 22692 21188 22716 21190
rect 22772 21188 22796 21190
rect 22852 21188 22858 21190
rect 22550 21179 22858 21188
rect 23492 21146 23520 21558
rect 23676 21486 23704 22034
rect 23952 21690 23980 22170
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 24136 21554 24164 22374
rect 24228 22234 24256 22714
rect 25872 22636 25924 22642
rect 25872 22578 25924 22584
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25700 22234 25728 22374
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 25688 22228 25740 22234
rect 25688 22170 25740 22176
rect 25320 22024 25372 22030
rect 25320 21966 25372 21972
rect 24950 21788 25258 21797
rect 24950 21786 24956 21788
rect 25012 21786 25036 21788
rect 25092 21786 25116 21788
rect 25172 21786 25196 21788
rect 25252 21786 25258 21788
rect 25012 21734 25014 21786
rect 25194 21734 25196 21786
rect 24950 21732 24956 21734
rect 25012 21732 25036 21734
rect 25092 21732 25116 21734
rect 25172 21732 25196 21734
rect 25252 21732 25258 21734
rect 24950 21723 25258 21732
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 24950 20700 25258 20709
rect 24950 20698 24956 20700
rect 25012 20698 25036 20700
rect 25092 20698 25116 20700
rect 25172 20698 25196 20700
rect 25252 20698 25258 20700
rect 25012 20646 25014 20698
rect 25194 20646 25196 20698
rect 24950 20644 24956 20646
rect 25012 20644 25036 20646
rect 25092 20644 25116 20646
rect 25172 20644 25196 20646
rect 25252 20644 25258 20646
rect 24950 20635 25258 20644
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20150 19612 20458 19621
rect 20150 19610 20156 19612
rect 20212 19610 20236 19612
rect 20292 19610 20316 19612
rect 20372 19610 20396 19612
rect 20452 19610 20458 19612
rect 20212 19558 20214 19610
rect 20394 19558 20396 19610
rect 20150 19556 20156 19558
rect 20212 19556 20236 19558
rect 20292 19556 20316 19558
rect 20372 19556 20396 19558
rect 20452 19556 20458 19558
rect 20150 19547 20458 19556
rect 21284 18834 21312 20402
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 24308 20392 24360 20398
rect 24308 20334 24360 20340
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 22480 20058 22508 20334
rect 22550 20156 22858 20165
rect 22550 20154 22556 20156
rect 22612 20154 22636 20156
rect 22692 20154 22716 20156
rect 22772 20154 22796 20156
rect 22852 20154 22858 20156
rect 22612 20102 22614 20154
rect 22794 20102 22796 20154
rect 22550 20100 22556 20102
rect 22612 20100 22636 20102
rect 22692 20100 22716 20102
rect 22772 20100 22796 20102
rect 22852 20100 22858 20102
rect 22550 20091 22858 20100
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23308 19378 23336 19858
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 22550 19068 22858 19077
rect 22550 19066 22556 19068
rect 22612 19066 22636 19068
rect 22692 19066 22716 19068
rect 22772 19066 22796 19068
rect 22852 19066 22858 19068
rect 22612 19014 22614 19066
rect 22794 19014 22796 19066
rect 22550 19012 22556 19014
rect 22612 19012 22636 19014
rect 22692 19012 22716 19014
rect 22772 19012 22796 19014
rect 22852 19012 22858 19014
rect 22550 19003 22858 19012
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20150 18524 20458 18533
rect 20150 18522 20156 18524
rect 20212 18522 20236 18524
rect 20292 18522 20316 18524
rect 20372 18522 20396 18524
rect 20452 18522 20458 18524
rect 20212 18470 20214 18522
rect 20394 18470 20396 18522
rect 20150 18468 20156 18470
rect 20212 18468 20236 18470
rect 20292 18468 20316 18470
rect 20372 18468 20396 18470
rect 20452 18468 20458 18470
rect 20150 18459 20458 18468
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 20548 18086 20576 18294
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19812 17202 19840 17478
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19168 16658 19196 16730
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 17604 16516 17736 16522
rect 17604 16510 17684 16516
rect 17684 16458 17736 16464
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18236 16448 18288 16454
rect 18156 16396 18236 16402
rect 18156 16390 18288 16396
rect 18156 16374 18276 16390
rect 18156 15910 18184 16374
rect 18708 16182 18736 16458
rect 19168 16250 19196 16594
rect 19352 16574 19380 17002
rect 19432 16584 19484 16590
rect 19352 16546 19432 16574
rect 19432 16526 19484 16532
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 17750 15804 18058 15813
rect 17750 15802 17756 15804
rect 17812 15802 17836 15804
rect 17892 15802 17916 15804
rect 17972 15802 17996 15804
rect 18052 15802 18058 15804
rect 17812 15750 17814 15802
rect 17994 15750 17996 15802
rect 17750 15748 17756 15750
rect 17812 15748 17836 15750
rect 17892 15748 17916 15750
rect 17972 15748 17996 15750
rect 18052 15748 18058 15750
rect 17750 15739 18058 15748
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17512 13938 17540 14350
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16500 12322 16528 12718
rect 16592 12434 16620 13126
rect 16776 12986 16804 13194
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16960 12646 16988 13126
rect 17052 12850 17080 13194
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16592 12406 16712 12434
rect 16500 12294 16620 12322
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 15948 9994 15976 10406
rect 16224 10146 16252 10746
rect 16316 10674 16344 11154
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16132 10130 16252 10146
rect 16120 10124 16252 10130
rect 16172 10118 16252 10124
rect 16120 10066 16172 10072
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15350 9820 15658 9829
rect 15350 9818 15356 9820
rect 15412 9818 15436 9820
rect 15492 9818 15516 9820
rect 15572 9818 15596 9820
rect 15652 9818 15658 9820
rect 15412 9766 15414 9818
rect 15594 9766 15596 9818
rect 15350 9764 15356 9766
rect 15412 9764 15436 9766
rect 15492 9764 15516 9766
rect 15572 9764 15596 9766
rect 15652 9764 15658 9766
rect 15350 9755 15658 9764
rect 15948 9654 15976 9930
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 16592 9586 16620 12294
rect 16684 11898 16712 12406
rect 16960 12306 16988 12582
rect 17052 12374 17080 12786
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16776 11778 16804 12174
rect 16684 11750 16804 11778
rect 16684 11014 16712 11750
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16776 11014 16804 11086
rect 16960 11014 16988 12242
rect 17052 12238 17080 12310
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16684 10606 16712 10950
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16776 10470 16804 10950
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 15350 8732 15658 8741
rect 15350 8730 15356 8732
rect 15412 8730 15436 8732
rect 15492 8730 15516 8732
rect 15572 8730 15596 8732
rect 15652 8730 15658 8732
rect 15412 8678 15414 8730
rect 15594 8678 15596 8730
rect 15350 8676 15356 8678
rect 15412 8676 15436 8678
rect 15492 8676 15516 8678
rect 15572 8676 15596 8678
rect 15652 8676 15658 8678
rect 15350 8667 15658 8676
rect 16592 8634 16620 9522
rect 16776 9518 16804 9862
rect 16960 9586 16988 10474
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17144 9518 17172 11834
rect 17236 9586 17264 13262
rect 17328 12850 17356 13330
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17328 12238 17356 12786
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17328 11150 17356 12174
rect 17512 12102 17540 13874
rect 17604 13462 17632 15098
rect 17750 14716 18058 14725
rect 17750 14714 17756 14716
rect 17812 14714 17836 14716
rect 17892 14714 17916 14716
rect 17972 14714 17996 14716
rect 18052 14714 18058 14716
rect 17812 14662 17814 14714
rect 17994 14662 17996 14714
rect 17750 14660 17756 14662
rect 17812 14660 17836 14662
rect 17892 14660 17916 14662
rect 17972 14660 17996 14662
rect 18052 14660 18058 14662
rect 17750 14651 18058 14660
rect 17750 13628 18058 13637
rect 17750 13626 17756 13628
rect 17812 13626 17836 13628
rect 17892 13626 17916 13628
rect 17972 13626 17996 13628
rect 18052 13626 18058 13628
rect 17812 13574 17814 13626
rect 17994 13574 17996 13626
rect 17750 13572 17756 13574
rect 17812 13572 17836 13574
rect 17892 13572 17916 13574
rect 17972 13572 17996 13574
rect 18052 13572 18058 13574
rect 17750 13563 18058 13572
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17750 12540 18058 12549
rect 17750 12538 17756 12540
rect 17812 12538 17836 12540
rect 17892 12538 17916 12540
rect 17972 12538 17996 12540
rect 18052 12538 18058 12540
rect 17812 12486 17814 12538
rect 17994 12486 17996 12538
rect 17750 12484 17756 12486
rect 17812 12484 17836 12486
rect 17892 12484 17916 12486
rect 17972 12484 17996 12486
rect 18052 12484 18058 12486
rect 17750 12475 18058 12484
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17788 11762 17816 12038
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 18156 11558 18184 15846
rect 19168 14958 19196 16186
rect 19444 15706 19472 16526
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19352 15026 19380 15574
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18432 14006 18460 14758
rect 19444 14618 19472 15642
rect 19812 15570 19840 17138
rect 19996 16998 20024 17750
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20150 17436 20458 17445
rect 20150 17434 20156 17436
rect 20212 17434 20236 17436
rect 20292 17434 20316 17436
rect 20372 17434 20396 17436
rect 20452 17434 20458 17436
rect 20212 17382 20214 17434
rect 20394 17382 20396 17434
rect 20150 17380 20156 17382
rect 20212 17380 20236 17382
rect 20292 17380 20316 17382
rect 20372 17380 20396 17382
rect 20452 17380 20458 17382
rect 20150 17371 20458 17380
rect 20548 17338 20576 17478
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 20088 15638 20116 17206
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20180 16998 20208 17138
rect 20640 17066 20668 18158
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17202 20760 17614
rect 20824 17202 20852 17750
rect 20916 17678 20944 18566
rect 21284 18442 21312 18770
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21284 18426 21404 18442
rect 21284 18420 21416 18426
rect 21284 18414 21364 18420
rect 21364 18362 21416 18368
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20150 16348 20458 16357
rect 20150 16346 20156 16348
rect 20212 16346 20236 16348
rect 20292 16346 20316 16348
rect 20372 16346 20396 16348
rect 20452 16346 20458 16348
rect 20212 16294 20214 16346
rect 20394 16294 20396 16346
rect 20150 16292 20156 16294
rect 20212 16292 20236 16294
rect 20292 16292 20316 16294
rect 20372 16292 20396 16294
rect 20452 16292 20458 16294
rect 20150 16283 20458 16292
rect 21008 16250 21036 17138
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 15706 20576 16050
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20076 15632 20128 15638
rect 20076 15574 20128 15580
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20150 15260 20458 15269
rect 20150 15258 20156 15260
rect 20212 15258 20236 15260
rect 20292 15258 20316 15260
rect 20372 15258 20396 15260
rect 20452 15258 20458 15260
rect 20212 15206 20214 15258
rect 20394 15206 20396 15258
rect 20150 15204 20156 15206
rect 20212 15204 20236 15206
rect 20292 15204 20316 15206
rect 20372 15204 20396 15206
rect 20452 15204 20458 15206
rect 20150 15195 20458 15204
rect 20824 15162 20852 15370
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 17750 11452 18058 11461
rect 17750 11450 17756 11452
rect 17812 11450 17836 11452
rect 17892 11450 17916 11452
rect 17972 11450 17996 11452
rect 18052 11450 18058 11452
rect 17812 11398 17814 11450
rect 17994 11398 17996 11450
rect 17750 11396 17756 11398
rect 17812 11396 17836 11398
rect 17892 11396 17916 11398
rect 17972 11396 17996 11398
rect 18052 11396 18058 11398
rect 17750 11387 18058 11396
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17604 11014 17632 11086
rect 18248 11082 18276 11766
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10130 17632 10950
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 17750 10364 18058 10373
rect 17750 10362 17756 10364
rect 17812 10362 17836 10364
rect 17892 10362 17916 10364
rect 17972 10362 17996 10364
rect 18052 10362 18058 10364
rect 17812 10310 17814 10362
rect 17994 10310 17996 10362
rect 17750 10308 17756 10310
rect 17812 10308 17836 10310
rect 17892 10308 17916 10310
rect 17972 10308 17996 10310
rect 18052 10308 18058 10310
rect 17750 10299 18058 10308
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 18156 10062 18184 10610
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17750 9276 18058 9285
rect 17750 9274 17756 9276
rect 17812 9274 17836 9276
rect 17892 9274 17916 9276
rect 17972 9274 17996 9276
rect 18052 9274 18058 9276
rect 17812 9222 17814 9274
rect 17994 9222 17996 9274
rect 17750 9220 17756 9222
rect 17812 9220 17836 9222
rect 17892 9220 17916 9222
rect 17972 9220 17996 9222
rect 18052 9220 18058 9222
rect 17750 9211 18058 9220
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 17750 8188 18058 8197
rect 17750 8186 17756 8188
rect 17812 8186 17836 8188
rect 17892 8186 17916 8188
rect 17972 8186 17996 8188
rect 18052 8186 18058 8188
rect 17812 8134 17814 8186
rect 17994 8134 17996 8186
rect 17750 8132 17756 8134
rect 17812 8132 17836 8134
rect 17892 8132 17916 8134
rect 17972 8132 17996 8134
rect 18052 8132 18058 8134
rect 17750 8123 18058 8132
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14200 7750 14228 7958
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14200 7546 14228 7686
rect 15350 7644 15658 7653
rect 15350 7642 15356 7644
rect 15412 7642 15436 7644
rect 15492 7642 15516 7644
rect 15572 7642 15596 7644
rect 15652 7642 15658 7644
rect 15412 7590 15414 7642
rect 15594 7590 15596 7642
rect 15350 7588 15356 7590
rect 15412 7588 15436 7590
rect 15492 7588 15516 7590
rect 15572 7588 15596 7590
rect 15652 7588 15658 7590
rect 15350 7579 15658 7588
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 17750 7100 18058 7109
rect 17750 7098 17756 7100
rect 17812 7098 17836 7100
rect 17892 7098 17916 7100
rect 17972 7098 17996 7100
rect 18052 7098 18058 7100
rect 17812 7046 17814 7098
rect 17994 7046 17996 7098
rect 17750 7044 17756 7046
rect 17812 7044 17836 7046
rect 17892 7044 17916 7046
rect 17972 7044 17996 7046
rect 18052 7044 18058 7046
rect 17750 7035 18058 7044
rect 15350 6556 15658 6565
rect 15350 6554 15356 6556
rect 15412 6554 15436 6556
rect 15492 6554 15516 6556
rect 15572 6554 15596 6556
rect 15652 6554 15658 6556
rect 15412 6502 15414 6554
rect 15594 6502 15596 6554
rect 15350 6500 15356 6502
rect 15412 6500 15436 6502
rect 15492 6500 15516 6502
rect 15572 6500 15596 6502
rect 15652 6500 15658 6502
rect 15350 6491 15658 6500
rect 17750 6012 18058 6021
rect 17750 6010 17756 6012
rect 17812 6010 17836 6012
rect 17892 6010 17916 6012
rect 17972 6010 17996 6012
rect 18052 6010 18058 6012
rect 17812 5958 17814 6010
rect 17994 5958 17996 6010
rect 17750 5956 17756 5958
rect 17812 5956 17836 5958
rect 17892 5956 17916 5958
rect 17972 5956 17996 5958
rect 18052 5956 18058 5958
rect 17750 5947 18058 5956
rect 15350 5468 15658 5477
rect 15350 5466 15356 5468
rect 15412 5466 15436 5468
rect 15492 5466 15516 5468
rect 15572 5466 15596 5468
rect 15652 5466 15658 5468
rect 15412 5414 15414 5466
rect 15594 5414 15596 5466
rect 15350 5412 15356 5414
rect 15412 5412 15436 5414
rect 15492 5412 15516 5414
rect 15572 5412 15596 5414
rect 15652 5412 15658 5414
rect 15350 5403 15658 5412
rect 17750 4924 18058 4933
rect 17750 4922 17756 4924
rect 17812 4922 17836 4924
rect 17892 4922 17916 4924
rect 17972 4922 17996 4924
rect 18052 4922 18058 4924
rect 17812 4870 17814 4922
rect 17994 4870 17996 4922
rect 17750 4868 17756 4870
rect 17812 4868 17836 4870
rect 17892 4868 17916 4870
rect 17972 4868 17996 4870
rect 18052 4868 18058 4870
rect 17750 4859 18058 4868
rect 15350 4380 15658 4389
rect 15350 4378 15356 4380
rect 15412 4378 15436 4380
rect 15492 4378 15516 4380
rect 15572 4378 15596 4380
rect 15652 4378 15658 4380
rect 15412 4326 15414 4378
rect 15594 4326 15596 4378
rect 15350 4324 15356 4326
rect 15412 4324 15436 4326
rect 15492 4324 15516 4326
rect 15572 4324 15596 4326
rect 15652 4324 15658 4326
rect 15350 4315 15658 4324
rect 17750 3836 18058 3845
rect 17750 3834 17756 3836
rect 17812 3834 17836 3836
rect 17892 3834 17916 3836
rect 17972 3834 17996 3836
rect 18052 3834 18058 3836
rect 17812 3782 17814 3834
rect 17994 3782 17996 3834
rect 17750 3780 17756 3782
rect 17812 3780 17836 3782
rect 17892 3780 17916 3782
rect 17972 3780 17996 3782
rect 18052 3780 18058 3782
rect 17750 3771 18058 3780
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 18248 3466 18276 11018
rect 18432 6730 18460 11494
rect 19260 10742 19288 11562
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 18524 3534 18552 9522
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19352 8294 19380 8910
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 7342 19380 8230
rect 19444 7546 19472 9998
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18616 6798 18644 7142
rect 19168 7002 19196 7278
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 6322 18644 6734
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18800 3534 18828 3878
rect 18892 3534 18920 6598
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19260 5778 19288 6258
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19352 5302 19380 7278
rect 19444 7018 19472 7482
rect 19444 6990 19656 7018
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19432 5840 19484 5846
rect 19432 5782 19484 5788
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19352 3602 19380 5238
rect 19444 5166 19472 5782
rect 19536 5710 19564 6054
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19628 5302 19656 6990
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19628 4214 19656 5238
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 15350 3292 15658 3301
rect 15350 3290 15356 3292
rect 15412 3290 15436 3292
rect 15492 3290 15516 3292
rect 15572 3290 15596 3292
rect 15652 3290 15658 3292
rect 15412 3238 15414 3290
rect 15594 3238 15596 3290
rect 15350 3236 15356 3238
rect 15412 3236 15436 3238
rect 15492 3236 15516 3238
rect 15572 3236 15596 3238
rect 15652 3236 15658 3238
rect 15350 3227 15658 3236
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 17750 2748 18058 2757
rect 17750 2746 17756 2748
rect 17812 2746 17836 2748
rect 17892 2746 17916 2748
rect 17972 2746 17996 2748
rect 18052 2746 18058 2748
rect 17812 2694 17814 2746
rect 17994 2694 17996 2746
rect 17750 2692 17756 2694
rect 17812 2692 17836 2694
rect 17892 2692 17916 2694
rect 17972 2692 17996 2694
rect 18052 2692 18058 2694
rect 17750 2683 18058 2692
rect 18524 2650 18552 3470
rect 18892 2990 18920 3470
rect 19720 3194 19748 14826
rect 20150 14172 20458 14181
rect 20150 14170 20156 14172
rect 20212 14170 20236 14172
rect 20292 14170 20316 14172
rect 20372 14170 20396 14172
rect 20452 14170 20458 14172
rect 20212 14118 20214 14170
rect 20394 14118 20396 14170
rect 20150 14116 20156 14118
rect 20212 14116 20236 14118
rect 20292 14116 20316 14118
rect 20372 14116 20396 14118
rect 20452 14116 20458 14118
rect 20150 14107 20458 14116
rect 20732 13938 20760 14962
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20824 13530 20852 15098
rect 21008 13870 21036 16186
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20150 13084 20458 13093
rect 20150 13082 20156 13084
rect 20212 13082 20236 13084
rect 20292 13082 20316 13084
rect 20372 13082 20396 13084
rect 20452 13082 20458 13084
rect 20212 13030 20214 13082
rect 20394 13030 20396 13082
rect 20150 13028 20156 13030
rect 20212 13028 20236 13030
rect 20292 13028 20316 13030
rect 20372 13028 20396 13030
rect 20452 13028 20458 13030
rect 20150 13019 20458 13028
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19996 10810 20024 12242
rect 20150 11996 20458 12005
rect 20150 11994 20156 11996
rect 20212 11994 20236 11996
rect 20292 11994 20316 11996
rect 20372 11994 20396 11996
rect 20452 11994 20458 11996
rect 20212 11942 20214 11994
rect 20394 11942 20396 11994
rect 20150 11940 20156 11942
rect 20212 11940 20236 11942
rect 20292 11940 20316 11942
rect 20372 11940 20396 11942
rect 20452 11940 20458 11942
rect 20150 11931 20458 11940
rect 20150 10908 20458 10917
rect 20150 10906 20156 10908
rect 20212 10906 20236 10908
rect 20292 10906 20316 10908
rect 20372 10906 20396 10908
rect 20452 10906 20458 10908
rect 20212 10854 20214 10906
rect 20394 10854 20396 10906
rect 20150 10852 20156 10854
rect 20212 10852 20236 10854
rect 20292 10852 20316 10854
rect 20372 10852 20396 10854
rect 20452 10852 20458 10854
rect 20150 10843 20458 10852
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 20088 10062 20116 10542
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10130 20392 10406
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20088 8974 20116 9998
rect 20150 9820 20458 9829
rect 20150 9818 20156 9820
rect 20212 9818 20236 9820
rect 20292 9818 20316 9820
rect 20372 9818 20396 9820
rect 20452 9818 20458 9820
rect 20212 9766 20214 9818
rect 20394 9766 20396 9818
rect 20150 9764 20156 9766
rect 20212 9764 20236 9766
rect 20292 9764 20316 9766
rect 20372 9764 20396 9766
rect 20452 9764 20458 9766
rect 20150 9755 20458 9764
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20150 8732 20458 8741
rect 20150 8730 20156 8732
rect 20212 8730 20236 8732
rect 20292 8730 20316 8732
rect 20372 8730 20396 8732
rect 20452 8730 20458 8732
rect 20212 8678 20214 8730
rect 20394 8678 20396 8730
rect 20150 8676 20156 8678
rect 20212 8676 20236 8678
rect 20292 8676 20316 8678
rect 20372 8676 20396 8678
rect 20452 8676 20458 8678
rect 20150 8667 20458 8676
rect 20444 8560 20496 8566
rect 20548 8514 20576 13466
rect 20824 13326 20852 13466
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 21008 12918 21036 13806
rect 21192 13734 21220 18022
rect 21376 17746 21404 18362
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21560 17678 21588 18634
rect 22550 17980 22858 17989
rect 22550 17978 22556 17980
rect 22612 17978 22636 17980
rect 22692 17978 22716 17980
rect 22772 17978 22796 17980
rect 22852 17978 22858 17980
rect 22612 17926 22614 17978
rect 22794 17926 22796 17978
rect 22550 17924 22556 17926
rect 22612 17924 22636 17926
rect 22692 17924 22716 17926
rect 22772 17924 22796 17926
rect 22852 17924 22858 17926
rect 22550 17915 22858 17924
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21284 15026 21312 17614
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21468 15502 21496 17546
rect 23308 17202 23336 19314
rect 24320 18630 24348 20334
rect 24872 19310 24900 20334
rect 25332 19922 25360 21966
rect 25884 21690 25912 22578
rect 26608 22500 26660 22506
rect 26608 22442 26660 22448
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 26068 21842 26096 21898
rect 26332 21888 26384 21894
rect 26068 21814 26280 21842
rect 26332 21830 26384 21836
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 26056 20868 26108 20874
rect 26056 20810 26108 20816
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 24950 19612 25258 19621
rect 24950 19610 24956 19612
rect 25012 19610 25036 19612
rect 25092 19610 25116 19612
rect 25172 19610 25196 19612
rect 25252 19610 25258 19612
rect 25012 19558 25014 19610
rect 25194 19558 25196 19610
rect 24950 19556 24956 19558
rect 25012 19556 25036 19558
rect 25092 19556 25116 19558
rect 25172 19556 25196 19558
rect 25252 19556 25258 19558
rect 24950 19547 25258 19556
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24872 18970 24900 19246
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24964 18834 24992 19110
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24320 18426 24348 18566
rect 24950 18524 25258 18533
rect 24950 18522 24956 18524
rect 25012 18522 25036 18524
rect 25092 18522 25116 18524
rect 25172 18522 25196 18524
rect 25252 18522 25258 18524
rect 25012 18470 25014 18522
rect 25194 18470 25196 18522
rect 24950 18468 24956 18470
rect 25012 18468 25036 18470
rect 25092 18468 25116 18470
rect 25172 18468 25196 18470
rect 25252 18468 25258 18470
rect 24950 18459 25258 18468
rect 24308 18420 24360 18426
rect 24308 18362 24360 18368
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 22550 16892 22858 16901
rect 22550 16890 22556 16892
rect 22612 16890 22636 16892
rect 22692 16890 22716 16892
rect 22772 16890 22796 16892
rect 22852 16890 22858 16892
rect 22612 16838 22614 16890
rect 22794 16838 22796 16890
rect 22550 16836 22556 16838
rect 22612 16836 22636 16838
rect 22692 16836 22716 16838
rect 22772 16836 22796 16838
rect 22852 16836 22858 16838
rect 22550 16827 22858 16836
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 21284 13938 21312 14486
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11898 20668 12038
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20824 11762 20852 12582
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 21008 10606 21036 12854
rect 21468 12850 21496 15438
rect 21560 14618 21588 15506
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 15162 21956 15302
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21928 14550 21956 14894
rect 21916 14544 21968 14550
rect 21916 14486 21968 14492
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21836 12918 21864 14214
rect 21928 13734 21956 14486
rect 22020 13870 22048 16594
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 22112 16250 22140 16458
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22204 15026 22232 16390
rect 22550 15804 22858 15813
rect 22550 15802 22556 15804
rect 22612 15802 22636 15804
rect 22692 15802 22716 15804
rect 22772 15802 22796 15804
rect 22852 15802 22858 15804
rect 22612 15750 22614 15802
rect 22794 15750 22796 15802
rect 22550 15748 22556 15750
rect 22612 15748 22636 15750
rect 22692 15748 22716 15750
rect 22772 15748 22796 15750
rect 22852 15748 22858 15750
rect 22550 15739 22858 15748
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22204 14414 22232 14962
rect 22296 14482 22324 15030
rect 23124 14890 23152 17070
rect 23308 16658 23336 17138
rect 24320 16794 24348 18362
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24872 17882 24900 18158
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24492 17672 24544 17678
rect 24492 17614 24544 17620
rect 24504 16794 24532 17614
rect 24872 17354 24900 17818
rect 24950 17436 25258 17445
rect 24950 17434 24956 17436
rect 25012 17434 25036 17436
rect 25092 17434 25116 17436
rect 25172 17434 25196 17436
rect 25252 17434 25258 17436
rect 25012 17382 25014 17434
rect 25194 17382 25196 17434
rect 24950 17380 24956 17382
rect 25012 17380 25036 17382
rect 25092 17380 25116 17382
rect 25172 17380 25196 17382
rect 25252 17380 25258 17382
rect 24950 17371 25258 17380
rect 24780 17338 24900 17354
rect 24768 17332 24900 17338
rect 24820 17326 24900 17332
rect 24768 17274 24820 17280
rect 26068 17270 26096 20810
rect 26252 19718 26280 21814
rect 26344 21690 26372 21830
rect 26332 21684 26384 21690
rect 26332 21626 26384 21632
rect 26620 21486 26648 22442
rect 27350 22332 27658 22341
rect 27350 22330 27356 22332
rect 27412 22330 27436 22332
rect 27492 22330 27516 22332
rect 27572 22330 27596 22332
rect 27652 22330 27658 22332
rect 27412 22278 27414 22330
rect 27594 22278 27596 22330
rect 27350 22276 27356 22278
rect 27412 22276 27436 22278
rect 27492 22276 27516 22278
rect 27572 22276 27596 22278
rect 27652 22276 27658 22278
rect 27350 22267 27658 22276
rect 27724 22114 27752 26318
rect 27632 22098 27752 22114
rect 27816 22098 27844 27406
rect 28356 26512 28408 26518
rect 28356 26454 28408 26460
rect 28368 25945 28396 26454
rect 28354 25936 28410 25945
rect 28354 25871 28410 25880
rect 28356 23520 28408 23526
rect 28354 23488 28356 23497
rect 28408 23488 28410 23497
rect 28354 23423 28410 23432
rect 27620 22092 27752 22098
rect 27672 22086 27752 22092
rect 27804 22092 27856 22098
rect 27620 22034 27672 22040
rect 27804 22034 27856 22040
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27252 21888 27304 21894
rect 27252 21830 27304 21836
rect 27264 21554 27292 21830
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 26608 21480 26660 21486
rect 27356 21434 27384 21966
rect 27632 21690 27660 22034
rect 27712 21888 27764 21894
rect 27712 21830 27764 21836
rect 27620 21684 27672 21690
rect 27620 21626 27672 21632
rect 27724 21622 27752 21830
rect 27712 21616 27764 21622
rect 27712 21558 27764 21564
rect 26608 21422 26660 21428
rect 27264 21418 27384 21434
rect 26332 21412 26384 21418
rect 26332 21354 26384 21360
rect 27252 21412 27384 21418
rect 27304 21406 27384 21412
rect 27252 21354 27304 21360
rect 26344 20942 26372 21354
rect 26608 21344 26660 21350
rect 26608 21286 26660 21292
rect 26620 21010 26648 21286
rect 26608 21004 26660 21010
rect 26608 20946 26660 20952
rect 26332 20936 26384 20942
rect 26332 20878 26384 20884
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26344 17678 26372 20878
rect 27264 20330 27292 21354
rect 27350 21244 27658 21253
rect 27350 21242 27356 21244
rect 27412 21242 27436 21244
rect 27492 21242 27516 21244
rect 27572 21242 27596 21244
rect 27652 21242 27658 21244
rect 27412 21190 27414 21242
rect 27594 21190 27596 21242
rect 27350 21188 27356 21190
rect 27412 21188 27436 21190
rect 27492 21188 27516 21190
rect 27572 21188 27596 21190
rect 27652 21188 27658 21190
rect 27350 21179 27658 21188
rect 27816 21146 27844 22034
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 28184 20602 28212 21490
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28368 21049 28396 21286
rect 28354 21040 28410 21049
rect 28354 20975 28410 20984
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 26424 20256 26476 20262
rect 26424 20198 26476 20204
rect 26436 19922 26464 20198
rect 26424 19916 26476 19922
rect 26424 19858 26476 19864
rect 27264 18154 27292 20266
rect 27350 20156 27658 20165
rect 27350 20154 27356 20156
rect 27412 20154 27436 20156
rect 27492 20154 27516 20156
rect 27572 20154 27596 20156
rect 27652 20154 27658 20156
rect 27412 20102 27414 20154
rect 27594 20102 27596 20154
rect 27350 20100 27356 20102
rect 27412 20100 27436 20102
rect 27492 20100 27516 20102
rect 27572 20100 27596 20102
rect 27652 20100 27658 20102
rect 27350 20091 27658 20100
rect 28184 20058 28212 20538
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27350 19068 27658 19077
rect 27350 19066 27356 19068
rect 27412 19066 27436 19068
rect 27492 19066 27516 19068
rect 27572 19066 27596 19068
rect 27652 19066 27658 19068
rect 27412 19014 27414 19066
rect 27594 19014 27596 19066
rect 27350 19012 27356 19014
rect 27412 19012 27436 19014
rect 27492 19012 27516 19014
rect 27572 19012 27596 19014
rect 27652 19012 27658 19014
rect 27350 19003 27658 19012
rect 27252 18148 27304 18154
rect 27252 18090 27304 18096
rect 26608 18080 26660 18086
rect 26608 18022 26660 18028
rect 26620 17746 26648 18022
rect 26608 17740 26660 17746
rect 26608 17682 26660 17688
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26056 17264 26108 17270
rect 26056 17206 26108 17212
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24308 16788 24360 16794
rect 24492 16788 24544 16794
rect 24360 16748 24440 16776
rect 24308 16730 24360 16736
rect 23296 16652 23348 16658
rect 23296 16594 23348 16600
rect 24136 14958 24164 16730
rect 24412 16674 24440 16748
rect 24492 16730 24544 16736
rect 24584 16720 24636 16726
rect 24412 16668 24584 16674
rect 24412 16662 24636 16668
rect 24412 16646 24624 16662
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24872 15722 24900 16526
rect 24964 16522 24992 16934
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24950 16348 25258 16357
rect 24950 16346 24956 16348
rect 25012 16346 25036 16348
rect 25092 16346 25116 16348
rect 25172 16346 25196 16348
rect 25252 16346 25258 16348
rect 25012 16294 25014 16346
rect 25194 16294 25196 16346
rect 24950 16292 24956 16294
rect 25012 16292 25036 16294
rect 25092 16292 25116 16294
rect 25172 16292 25196 16294
rect 25252 16292 25258 16294
rect 24950 16283 25258 16292
rect 25964 16244 26016 16250
rect 25964 16186 26016 16192
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 24872 15694 24992 15722
rect 24860 15632 24912 15638
rect 24860 15574 24912 15580
rect 24872 15162 24900 15574
rect 24964 15502 24992 15694
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 24950 15260 25258 15269
rect 24950 15258 24956 15260
rect 25012 15258 25036 15260
rect 25092 15258 25116 15260
rect 25172 15258 25196 15260
rect 25252 15258 25258 15260
rect 25012 15206 25014 15258
rect 25194 15206 25196 15258
rect 24950 15204 24956 15206
rect 25012 15204 25036 15206
rect 25092 15204 25116 15206
rect 25172 15204 25196 15206
rect 25252 15204 25258 15206
rect 24950 15195 25258 15204
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 23112 14884 23164 14890
rect 23112 14826 23164 14832
rect 22550 14716 22858 14725
rect 22550 14714 22556 14716
rect 22612 14714 22636 14716
rect 22692 14714 22716 14716
rect 22772 14714 22796 14716
rect 22852 14714 22858 14716
rect 22612 14662 22614 14714
rect 22794 14662 22796 14714
rect 22550 14660 22556 14662
rect 22612 14660 22636 14662
rect 22692 14660 22716 14662
rect 22772 14660 22796 14662
rect 22852 14660 22858 14662
rect 22550 14651 22858 14660
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 21916 13728 21968 13734
rect 21916 13670 21968 13676
rect 21928 13326 21956 13670
rect 22020 13530 22048 13806
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21824 12912 21876 12918
rect 21824 12854 21876 12860
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21468 10606 21496 12786
rect 21836 12646 21864 12854
rect 21928 12714 21956 13262
rect 22112 12782 22140 14282
rect 22296 13938 22324 14418
rect 24228 14074 24256 14962
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22550 13628 22858 13637
rect 22550 13626 22556 13628
rect 22612 13626 22636 13628
rect 22692 13626 22716 13628
rect 22772 13626 22796 13628
rect 22852 13626 22858 13628
rect 22612 13574 22614 13626
rect 22794 13574 22796 13626
rect 22550 13572 22556 13574
rect 22612 13572 22636 13574
rect 22692 13572 22716 13574
rect 22772 13572 22796 13574
rect 22852 13572 22858 13574
rect 22550 13563 22858 13572
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 23032 12986 23060 13126
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22296 12782 22324 12854
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 21916 12708 21968 12714
rect 21916 12650 21968 12656
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21836 10674 21864 12582
rect 22296 12238 22324 12718
rect 22550 12540 22858 12549
rect 22550 12538 22556 12540
rect 22612 12538 22636 12540
rect 22692 12538 22716 12540
rect 22772 12538 22796 12540
rect 22852 12538 22858 12540
rect 22612 12486 22614 12538
rect 22794 12486 22796 12538
rect 22550 12484 22556 12486
rect 22612 12484 22636 12486
rect 22692 12484 22716 12486
rect 22772 12484 22796 12486
rect 22852 12484 22858 12486
rect 22550 12475 22858 12484
rect 24412 12306 24440 14758
rect 24950 14172 25258 14181
rect 24950 14170 24956 14172
rect 25012 14170 25036 14172
rect 25092 14170 25116 14172
rect 25172 14170 25196 14172
rect 25252 14170 25258 14172
rect 25012 14118 25014 14170
rect 25194 14118 25196 14170
rect 24950 14116 24956 14118
rect 25012 14116 25036 14118
rect 25092 14116 25116 14118
rect 25172 14116 25196 14118
rect 25252 14116 25258 14118
rect 24950 14107 25258 14116
rect 25332 14006 25360 15302
rect 25516 15162 25544 16050
rect 25976 15434 26004 16186
rect 26344 15570 26372 17614
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26620 15502 26648 16526
rect 27264 16182 27292 18090
rect 27350 17980 27658 17989
rect 27350 17978 27356 17980
rect 27412 17978 27436 17980
rect 27492 17978 27516 17980
rect 27572 17978 27596 17980
rect 27652 17978 27658 17980
rect 27412 17926 27414 17978
rect 27594 17926 27596 17978
rect 27350 17924 27356 17926
rect 27412 17924 27436 17926
rect 27492 17924 27516 17926
rect 27572 17924 27596 17926
rect 27652 17924 27658 17926
rect 27350 17915 27658 17924
rect 27724 17678 27752 19654
rect 28172 18760 28224 18766
rect 28172 18702 28224 18708
rect 28184 18290 28212 18702
rect 28356 18624 28408 18630
rect 28354 18592 28356 18601
rect 28408 18592 28410 18601
rect 28354 18527 28410 18536
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28184 17882 28212 18226
rect 28172 17876 28224 17882
rect 28172 17818 28224 17824
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27350 16892 27658 16901
rect 27350 16890 27356 16892
rect 27412 16890 27436 16892
rect 27492 16890 27516 16892
rect 27572 16890 27596 16892
rect 27652 16890 27658 16892
rect 27412 16838 27414 16890
rect 27594 16838 27596 16890
rect 27350 16836 27356 16838
rect 27412 16836 27436 16838
rect 27492 16836 27516 16838
rect 27572 16836 27596 16838
rect 27652 16836 27658 16838
rect 27350 16827 27658 16836
rect 27724 16574 27752 17614
rect 28172 16584 28224 16590
rect 27724 16546 27936 16574
rect 27252 16176 27304 16182
rect 27252 16118 27304 16124
rect 27264 16046 27292 16118
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 26884 15904 26936 15910
rect 26884 15846 26936 15852
rect 26896 15570 26924 15846
rect 27350 15804 27658 15813
rect 27350 15802 27356 15804
rect 27412 15802 27436 15804
rect 27492 15802 27516 15804
rect 27572 15802 27596 15804
rect 27652 15802 27658 15804
rect 27412 15750 27414 15802
rect 27594 15750 27596 15802
rect 27350 15748 27356 15750
rect 27412 15748 27436 15750
rect 27492 15748 27516 15750
rect 27572 15748 27596 15750
rect 27652 15748 27658 15750
rect 27350 15739 27658 15748
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 27908 15502 27936 16546
rect 28172 16526 28224 16532
rect 28184 16114 28212 16526
rect 28356 16448 28408 16454
rect 28356 16390 28408 16396
rect 28368 16153 28396 16390
rect 28354 16144 28410 16153
rect 28172 16108 28224 16114
rect 28354 16079 28410 16088
rect 28172 16050 28224 16056
rect 28184 15706 28212 16050
rect 28172 15700 28224 15706
rect 28172 15642 28224 15648
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 27896 15496 27948 15502
rect 27896 15438 27948 15444
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 25332 13258 25360 13942
rect 26620 13326 26648 15438
rect 27350 14716 27658 14725
rect 27350 14714 27356 14716
rect 27412 14714 27436 14716
rect 27492 14714 27516 14716
rect 27572 14714 27596 14716
rect 27652 14714 27658 14716
rect 27412 14662 27414 14714
rect 27594 14662 27596 14714
rect 27350 14660 27356 14662
rect 27412 14660 27436 14662
rect 27492 14660 27516 14662
rect 27572 14660 27596 14662
rect 27652 14660 27658 14662
rect 27350 14651 27658 14660
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 28172 13932 28224 13938
rect 28172 13874 28224 13880
rect 26884 13728 26936 13734
rect 26884 13670 26936 13676
rect 26896 13394 26924 13670
rect 26884 13388 26936 13394
rect 26884 13330 26936 13336
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 25320 13252 25372 13258
rect 25320 13194 25372 13200
rect 24950 13084 25258 13093
rect 24950 13082 24956 13084
rect 25012 13082 25036 13084
rect 25092 13082 25116 13084
rect 25172 13082 25196 13084
rect 25252 13082 25258 13084
rect 25012 13030 25014 13082
rect 25194 13030 25196 13082
rect 24950 13028 24956 13030
rect 25012 13028 25036 13030
rect 25092 13028 25116 13030
rect 25172 13028 25196 13030
rect 25252 13028 25258 13030
rect 24950 13019 25258 13028
rect 25332 12918 25360 13194
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24872 12306 24900 12582
rect 25424 12442 25452 13262
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25884 12918 25912 13126
rect 25872 12912 25924 12918
rect 25872 12854 25924 12860
rect 26620 12850 26648 13262
rect 27264 12986 27292 13874
rect 27350 13628 27658 13637
rect 27350 13626 27356 13628
rect 27412 13626 27436 13628
rect 27492 13626 27516 13628
rect 27572 13626 27596 13628
rect 27652 13626 27658 13628
rect 27412 13574 27414 13626
rect 27594 13574 27596 13626
rect 27350 13572 27356 13574
rect 27412 13572 27436 13574
rect 27492 13572 27516 13574
rect 27572 13572 27596 13574
rect 27652 13572 27658 13574
rect 27350 13563 27658 13572
rect 28184 13190 28212 13874
rect 28356 13728 28408 13734
rect 28354 13696 28356 13705
rect 28408 13696 28410 13705
rect 28354 13631 28410 13640
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 28172 13184 28224 13190
rect 28172 13126 28224 13132
rect 27724 12986 27752 13126
rect 27252 12980 27304 12986
rect 27252 12922 27304 12928
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 23388 12164 23440 12170
rect 23388 12106 23440 12112
rect 22550 11452 22858 11461
rect 22550 11450 22556 11452
rect 22612 11450 22636 11452
rect 22692 11450 22716 11452
rect 22772 11450 22796 11452
rect 22852 11450 22858 11452
rect 22612 11398 22614 11450
rect 22794 11398 22796 11450
rect 22550 11396 22556 11398
rect 22612 11396 22636 11398
rect 22692 11396 22716 11398
rect 22772 11396 22796 11398
rect 22852 11396 22858 11398
rect 22550 11387 22858 11396
rect 23400 11082 23428 12106
rect 24228 12102 24256 12242
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20496 8508 20576 8514
rect 20444 8502 20576 8508
rect 20456 8486 20576 8502
rect 20916 8498 20944 10474
rect 20904 8492 20956 8498
rect 20456 8090 20484 8486
rect 20904 8434 20956 8440
rect 21008 8294 21036 10542
rect 21836 10266 21864 10610
rect 22550 10364 22858 10373
rect 22550 10362 22556 10364
rect 22612 10362 22636 10364
rect 22692 10362 22716 10364
rect 22772 10362 22796 10364
rect 22852 10362 22858 10364
rect 22612 10310 22614 10362
rect 22794 10310 22796 10362
rect 22550 10308 22556 10310
rect 22612 10308 22636 10310
rect 22692 10308 22716 10310
rect 22772 10308 22796 10310
rect 22852 10308 22858 10310
rect 22550 10299 22858 10308
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 23400 9994 23428 11018
rect 23492 10810 23520 11154
rect 23860 11082 23888 11494
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23952 10810 23980 11698
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 24228 10606 24256 12038
rect 24950 11996 25258 12005
rect 24950 11994 24956 11996
rect 25012 11994 25036 11996
rect 25092 11994 25116 11996
rect 25172 11994 25196 11996
rect 25252 11994 25258 11996
rect 25012 11942 25014 11994
rect 25194 11942 25196 11994
rect 24950 11940 24956 11942
rect 25012 11940 25036 11942
rect 25092 11940 25116 11942
rect 25172 11940 25196 11942
rect 25252 11940 25258 11942
rect 24950 11931 25258 11940
rect 26712 11694 26740 12582
rect 27350 12540 27658 12549
rect 27350 12538 27356 12540
rect 27412 12538 27436 12540
rect 27492 12538 27516 12540
rect 27572 12538 27596 12540
rect 27652 12538 27658 12540
rect 27412 12486 27414 12538
rect 27594 12486 27596 12538
rect 27350 12484 27356 12486
rect 27412 12484 27436 12486
rect 27492 12484 27516 12486
rect 27572 12484 27596 12486
rect 27652 12484 27658 12486
rect 27350 12475 27658 12484
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 28172 11756 28224 11762
rect 28172 11698 28224 11704
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 24950 10908 25258 10917
rect 24950 10906 24956 10908
rect 25012 10906 25036 10908
rect 25092 10906 25116 10908
rect 25172 10906 25196 10908
rect 25252 10906 25258 10908
rect 25012 10854 25014 10906
rect 25194 10854 25196 10906
rect 24950 10852 24956 10854
rect 25012 10852 25036 10854
rect 25092 10852 25116 10854
rect 25172 10852 25196 10854
rect 25252 10852 25258 10854
rect 24950 10843 25258 10852
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 22550 9276 22858 9285
rect 22550 9274 22556 9276
rect 22612 9274 22636 9276
rect 22692 9274 22716 9276
rect 22772 9274 22796 9276
rect 22852 9274 22858 9276
rect 22612 9222 22614 9274
rect 22794 9222 22796 9274
rect 22550 9220 22556 9222
rect 22612 9220 22636 9222
rect 22692 9220 22716 9222
rect 22772 9220 22796 9222
rect 22852 9220 22858 9222
rect 22550 9211 22858 9220
rect 23400 8974 23428 9930
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 21836 8634 21864 8842
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21180 8560 21232 8566
rect 21180 8502 21232 8508
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20456 7886 20484 8026
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20150 7644 20458 7653
rect 20150 7642 20156 7644
rect 20212 7642 20236 7644
rect 20292 7642 20316 7644
rect 20372 7642 20396 7644
rect 20452 7642 20458 7644
rect 20212 7590 20214 7642
rect 20394 7590 20396 7642
rect 20150 7588 20156 7590
rect 20212 7588 20236 7590
rect 20292 7588 20316 7590
rect 20372 7588 20396 7590
rect 20452 7588 20458 7590
rect 20150 7579 20458 7588
rect 21008 7002 21036 8230
rect 21192 7546 21220 8502
rect 23308 8498 23336 8774
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 22112 8090 22140 8434
rect 22550 8188 22858 8197
rect 22550 8186 22556 8188
rect 22612 8186 22636 8188
rect 22692 8186 22716 8188
rect 22772 8186 22796 8188
rect 22852 8186 22858 8188
rect 22612 8134 22614 8186
rect 22794 8134 22796 8186
rect 22550 8132 22556 8134
rect 22612 8132 22636 8134
rect 22692 8132 22716 8134
rect 22772 8132 22796 8134
rect 22852 8132 22858 8134
rect 22550 8123 22858 8132
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 22020 7274 22048 7754
rect 22112 7342 22140 7822
rect 23308 7818 23336 8434
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23296 7812 23348 7818
rect 23296 7754 23348 7760
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 21008 6866 21036 6938
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20150 6556 20458 6565
rect 20150 6554 20156 6556
rect 20212 6554 20236 6556
rect 20292 6554 20316 6556
rect 20372 6554 20396 6556
rect 20452 6554 20458 6556
rect 20212 6502 20214 6554
rect 20394 6502 20396 6554
rect 20150 6500 20156 6502
rect 20212 6500 20236 6502
rect 20292 6500 20316 6502
rect 20372 6500 20396 6502
rect 20452 6500 20458 6502
rect 20150 6491 20458 6500
rect 20824 6458 20852 6666
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20732 5574 20760 6258
rect 21008 6254 21036 6802
rect 22020 6730 22048 7210
rect 22112 6866 22140 7278
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 21560 6322 21588 6666
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21652 6322 21680 6598
rect 22112 6390 22140 6802
rect 22204 6798 22232 7346
rect 22296 6866 22324 7686
rect 23032 7410 23060 7686
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 22550 7100 22858 7109
rect 22550 7098 22556 7100
rect 22612 7098 22636 7100
rect 22692 7098 22716 7100
rect 22772 7098 22796 7100
rect 22852 7098 22858 7100
rect 22612 7046 22614 7098
rect 22794 7046 22796 7098
rect 22550 7044 22556 7046
rect 22612 7044 22636 7046
rect 22692 7044 22716 7046
rect 22772 7044 22796 7046
rect 22852 7044 22858 7046
rect 22550 7035 22858 7044
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22204 6458 22232 6734
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 20996 6248 21048 6254
rect 20996 6190 21048 6196
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20150 5468 20458 5477
rect 20150 5466 20156 5468
rect 20212 5466 20236 5468
rect 20292 5466 20316 5468
rect 20372 5466 20396 5468
rect 20452 5466 20458 5468
rect 20212 5414 20214 5466
rect 20394 5414 20396 5466
rect 20150 5412 20156 5414
rect 20212 5412 20236 5414
rect 20292 5412 20316 5414
rect 20372 5412 20396 5414
rect 20452 5412 20458 5414
rect 20150 5403 20458 5412
rect 20732 5370 20760 5510
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20732 4622 20760 5306
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 20150 4380 20458 4389
rect 20150 4378 20156 4380
rect 20212 4378 20236 4380
rect 20292 4378 20316 4380
rect 20372 4378 20396 4380
rect 20452 4378 20458 4380
rect 20212 4326 20214 4378
rect 20394 4326 20396 4378
rect 20150 4324 20156 4326
rect 20212 4324 20236 4326
rect 20292 4324 20316 4326
rect 20372 4324 20396 4326
rect 20452 4324 20458 4326
rect 20150 4315 20458 4324
rect 20076 4208 20128 4214
rect 20076 4150 20128 4156
rect 20088 3466 20116 4150
rect 22112 4146 22140 4422
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 21100 3738 21128 4082
rect 21640 4004 21692 4010
rect 21640 3946 21692 3952
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 19720 2922 19748 3130
rect 20088 3126 20116 3402
rect 21100 3398 21128 3674
rect 21652 3602 21680 3946
rect 22296 3602 22324 6802
rect 22652 6724 22704 6730
rect 22652 6666 22704 6672
rect 22664 6458 22692 6666
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22550 6012 22858 6021
rect 22550 6010 22556 6012
rect 22612 6010 22636 6012
rect 22692 6010 22716 6012
rect 22772 6010 22796 6012
rect 22852 6010 22858 6012
rect 22612 5958 22614 6010
rect 22794 5958 22796 6010
rect 22550 5956 22556 5958
rect 22612 5956 22636 5958
rect 22692 5956 22716 5958
rect 22772 5956 22796 5958
rect 22852 5956 22858 5958
rect 22550 5947 22858 5956
rect 22550 4924 22858 4933
rect 22550 4922 22556 4924
rect 22612 4922 22636 4924
rect 22692 4922 22716 4924
rect 22772 4922 22796 4924
rect 22852 4922 22858 4924
rect 22612 4870 22614 4922
rect 22794 4870 22796 4922
rect 22550 4868 22556 4870
rect 22612 4868 22636 4870
rect 22692 4868 22716 4870
rect 22772 4868 22796 4870
rect 22852 4868 22858 4870
rect 22550 4859 22858 4868
rect 23032 4622 23060 7346
rect 23308 7342 23336 7754
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 23400 6662 23428 7822
rect 23952 6730 23980 8842
rect 24228 8430 24256 10542
rect 24950 9820 25258 9829
rect 24950 9818 24956 9820
rect 25012 9818 25036 9820
rect 25092 9818 25116 9820
rect 25172 9818 25196 9820
rect 25252 9818 25258 9820
rect 25012 9766 25014 9818
rect 25194 9766 25196 9818
rect 24950 9764 24956 9766
rect 25012 9764 25036 9766
rect 25092 9764 25116 9766
rect 25172 9764 25196 9766
rect 25252 9764 25258 9766
rect 24950 9755 25258 9764
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24504 8634 24532 8774
rect 24872 8634 24900 9522
rect 25964 9376 26016 9382
rect 25964 9318 26016 9324
rect 25976 9042 26004 9318
rect 25964 9036 26016 9042
rect 25964 8978 26016 8984
rect 25976 8838 26004 8978
rect 26528 8974 26556 11086
rect 26712 10470 26740 11630
rect 26792 11552 26844 11558
rect 26792 11494 26844 11500
rect 26804 11218 26832 11494
rect 26792 11212 26844 11218
rect 26792 11154 26844 11160
rect 27172 10810 27200 11698
rect 27350 11452 27658 11461
rect 27350 11450 27356 11452
rect 27412 11450 27436 11452
rect 27492 11450 27516 11452
rect 27572 11450 27596 11452
rect 27652 11450 27658 11452
rect 27412 11398 27414 11450
rect 27594 11398 27596 11450
rect 27350 11396 27356 11398
rect 27412 11396 27436 11398
rect 27492 11396 27516 11398
rect 27572 11396 27596 11398
rect 27652 11396 27658 11398
rect 27350 11387 27658 11396
rect 27804 11076 27856 11082
rect 27804 11018 27856 11024
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27632 10810 27660 10950
rect 27724 10810 27752 10950
rect 27160 10804 27212 10810
rect 27160 10746 27212 10752
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 24950 8732 25258 8741
rect 24950 8730 24956 8732
rect 25012 8730 25036 8732
rect 25092 8730 25116 8732
rect 25172 8730 25196 8732
rect 25252 8730 25258 8732
rect 25012 8678 25014 8730
rect 25194 8678 25196 8730
rect 24950 8676 24956 8678
rect 25012 8676 25036 8678
rect 25092 8676 25116 8678
rect 25172 8676 25196 8678
rect 25252 8676 25258 8678
rect 24950 8667 25258 8676
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 23940 6724 23992 6730
rect 23940 6666 23992 6672
rect 24584 6724 24636 6730
rect 24584 6666 24636 6672
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 24136 5710 24164 6598
rect 24596 6322 24624 6666
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24688 5914 24716 8366
rect 24950 7644 25258 7653
rect 24950 7642 24956 7644
rect 25012 7642 25036 7644
rect 25092 7642 25116 7644
rect 25172 7642 25196 7644
rect 25252 7642 25258 7644
rect 25012 7590 25014 7642
rect 25194 7590 25196 7642
rect 24950 7588 24956 7590
rect 25012 7588 25036 7590
rect 25092 7588 25116 7590
rect 25172 7588 25196 7590
rect 25252 7588 25258 7590
rect 24950 7579 25258 7588
rect 26528 6914 26556 8910
rect 26712 8430 26740 10406
rect 27350 10364 27658 10373
rect 27350 10362 27356 10364
rect 27412 10362 27436 10364
rect 27492 10362 27516 10364
rect 27572 10362 27596 10364
rect 27652 10362 27658 10364
rect 27412 10310 27414 10362
rect 27594 10310 27596 10362
rect 27350 10308 27356 10310
rect 27412 10308 27436 10310
rect 27492 10308 27516 10310
rect 27572 10308 27596 10310
rect 27652 10308 27658 10310
rect 27350 10299 27658 10308
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26804 9042 26832 9318
rect 26792 9036 26844 9042
rect 26792 8978 26844 8984
rect 27172 8634 27200 9522
rect 27350 9276 27658 9285
rect 27350 9274 27356 9276
rect 27412 9274 27436 9276
rect 27492 9274 27516 9276
rect 27572 9274 27596 9276
rect 27652 9274 27658 9276
rect 27412 9222 27414 9274
rect 27594 9222 27596 9274
rect 27350 9220 27356 9222
rect 27412 9220 27436 9222
rect 27492 9220 27516 9222
rect 27572 9220 27596 9222
rect 27652 9220 27658 9222
rect 27350 9211 27658 9220
rect 27816 8906 27844 11018
rect 28184 11014 28212 11698
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 28368 11257 28396 11494
rect 28354 11248 28410 11257
rect 28354 11183 28410 11192
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 28264 9580 28316 9586
rect 28264 9522 28316 9528
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27632 8634 27660 8774
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27350 8188 27658 8197
rect 27350 8186 27356 8188
rect 27412 8186 27436 8188
rect 27492 8186 27516 8188
rect 27572 8186 27596 8188
rect 27652 8186 27658 8188
rect 27412 8134 27414 8186
rect 27594 8134 27596 8186
rect 27350 8132 27356 8134
rect 27412 8132 27436 8134
rect 27492 8132 27516 8134
rect 27572 8132 27596 8134
rect 27652 8132 27658 8134
rect 27350 8123 27658 8132
rect 27350 7100 27658 7109
rect 27350 7098 27356 7100
rect 27412 7098 27436 7100
rect 27492 7098 27516 7100
rect 27572 7098 27596 7100
rect 27652 7098 27658 7100
rect 27412 7046 27414 7098
rect 27594 7046 27596 7098
rect 27350 7044 27356 7046
rect 27412 7044 27436 7046
rect 27492 7044 27516 7046
rect 27572 7044 27596 7046
rect 27652 7044 27658 7046
rect 27350 7035 27658 7044
rect 26528 6886 26648 6914
rect 25688 6792 25740 6798
rect 25688 6734 25740 6740
rect 24950 6556 25258 6565
rect 24950 6554 24956 6556
rect 25012 6554 25036 6556
rect 25092 6554 25116 6556
rect 25172 6554 25196 6556
rect 25252 6554 25258 6556
rect 25012 6502 25014 6554
rect 25194 6502 25196 6554
rect 24950 6500 24956 6502
rect 25012 6500 25036 6502
rect 25092 6500 25116 6502
rect 25172 6500 25196 6502
rect 25252 6500 25258 6502
rect 24950 6491 25258 6500
rect 25228 6112 25280 6118
rect 25228 6054 25280 6060
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4690 23612 4966
rect 24688 4690 24716 5850
rect 25240 5778 25268 6054
rect 25700 5914 25728 6734
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26252 6390 26280 6598
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 26620 6254 26648 6886
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27724 6746 27752 8366
rect 27816 6914 27844 8842
rect 28276 8838 28304 9522
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 28264 8832 28316 8838
rect 28368 8809 28396 9318
rect 28264 8774 28316 8780
rect 28354 8800 28410 8809
rect 28276 8634 28304 8774
rect 28354 8735 28410 8744
rect 28264 8628 28316 8634
rect 28264 8570 28316 8576
rect 27816 6886 27936 6914
rect 26884 6656 26936 6662
rect 26884 6598 26936 6604
rect 26608 6248 26660 6254
rect 26608 6190 26660 6196
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 26620 5710 26648 6190
rect 26896 5778 26924 6598
rect 27264 6458 27292 6734
rect 27724 6718 27844 6746
rect 27816 6662 27844 6718
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 27816 6254 27844 6598
rect 27804 6248 27856 6254
rect 27804 6190 27856 6196
rect 27350 6012 27658 6021
rect 27350 6010 27356 6012
rect 27412 6010 27436 6012
rect 27492 6010 27516 6012
rect 27572 6010 27596 6012
rect 27652 6010 27658 6012
rect 27412 5958 27414 6010
rect 27594 5958 27596 6010
rect 27350 5956 27356 5958
rect 27412 5956 27436 5958
rect 27492 5956 27516 5958
rect 27572 5956 27596 5958
rect 27652 5956 27658 5958
rect 27350 5947 27658 5956
rect 26884 5772 26936 5778
rect 26884 5714 26936 5720
rect 26608 5704 26660 5710
rect 26608 5646 26660 5652
rect 24950 5468 25258 5477
rect 24950 5466 24956 5468
rect 25012 5466 25036 5468
rect 25092 5466 25116 5468
rect 25172 5466 25196 5468
rect 25252 5466 25258 5468
rect 25012 5414 25014 5466
rect 25194 5414 25196 5466
rect 24950 5412 24956 5414
rect 25012 5412 25036 5414
rect 25092 5412 25116 5414
rect 25172 5412 25196 5414
rect 25252 5412 25258 5414
rect 24950 5403 25258 5412
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 26620 4622 26648 5646
rect 27350 4924 27658 4933
rect 27350 4922 27356 4924
rect 27412 4922 27436 4924
rect 27492 4922 27516 4924
rect 27572 4922 27596 4924
rect 27652 4922 27658 4924
rect 27412 4870 27414 4922
rect 27594 4870 27596 4922
rect 27350 4868 27356 4870
rect 27412 4868 27436 4870
rect 27492 4868 27516 4870
rect 27572 4868 27596 4870
rect 27652 4868 27658 4870
rect 27350 4859 27658 4868
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 22550 3836 22858 3845
rect 22550 3834 22556 3836
rect 22612 3834 22636 3836
rect 22692 3834 22716 3836
rect 22772 3834 22796 3836
rect 22852 3834 22858 3836
rect 22612 3782 22614 3834
rect 22794 3782 22796 3834
rect 22550 3780 22556 3782
rect 22612 3780 22636 3782
rect 22692 3780 22716 3782
rect 22772 3780 22796 3782
rect 22852 3780 22858 3782
rect 22550 3771 22858 3780
rect 23032 3738 23060 4422
rect 23216 4146 23244 4422
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23388 4004 23440 4010
rect 23388 3946 23440 3952
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 21640 3596 21692 3602
rect 21640 3538 21692 3544
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 20150 3292 20458 3301
rect 20150 3290 20156 3292
rect 20212 3290 20236 3292
rect 20292 3290 20316 3292
rect 20372 3290 20396 3292
rect 20452 3290 20458 3292
rect 20212 3238 20214 3290
rect 20394 3238 20396 3290
rect 20150 3236 20156 3238
rect 20212 3236 20236 3238
rect 20292 3236 20316 3238
rect 20372 3236 20396 3238
rect 20452 3236 20458 3238
rect 20150 3227 20458 3236
rect 20076 3120 20128 3126
rect 20076 3062 20128 3068
rect 22296 3058 22324 3538
rect 23400 3194 23428 3946
rect 23584 3194 23612 4422
rect 24950 4380 25258 4389
rect 24950 4378 24956 4380
rect 25012 4378 25036 4380
rect 25092 4378 25116 4380
rect 25172 4378 25196 4380
rect 25252 4378 25258 4380
rect 25012 4326 25014 4378
rect 25194 4326 25196 4378
rect 24950 4324 24956 4326
rect 25012 4324 25036 4326
rect 25092 4324 25116 4326
rect 25172 4324 25196 4326
rect 25252 4324 25258 4326
rect 24950 4315 25258 4324
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 23848 3936 23900 3942
rect 23848 3878 23900 3884
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 23860 3466 23888 3878
rect 25148 3466 25176 3878
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 25136 3460 25188 3466
rect 25136 3402 25188 3408
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23860 3126 23888 3402
rect 24950 3292 25258 3301
rect 24950 3290 24956 3292
rect 25012 3290 25036 3292
rect 25092 3290 25116 3292
rect 25172 3290 25196 3292
rect 25252 3290 25258 3292
rect 25012 3238 25014 3290
rect 25194 3238 25196 3290
rect 24950 3236 24956 3238
rect 25012 3236 25036 3238
rect 25092 3236 25116 3238
rect 25172 3236 25196 3238
rect 25252 3236 25258 3238
rect 24950 3227 25258 3236
rect 25424 3194 25452 4082
rect 25780 4004 25832 4010
rect 25780 3946 25832 3952
rect 25792 3194 25820 3946
rect 26252 3670 26280 4558
rect 26976 4548 27028 4554
rect 26976 4490 27028 4496
rect 26988 3738 27016 4490
rect 27816 4078 27844 6190
rect 27908 6118 27936 6886
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28276 6202 28304 6734
rect 28356 6656 28408 6662
rect 28356 6598 28408 6604
rect 28368 6361 28396 6598
rect 28354 6352 28410 6361
rect 28354 6287 28410 6296
rect 28276 6186 28396 6202
rect 28276 6180 28408 6186
rect 28276 6174 28356 6180
rect 28356 6122 28408 6128
rect 27896 6112 27948 6118
rect 27896 6054 27948 6060
rect 27908 5642 27936 6054
rect 28368 5914 28396 6122
rect 28356 5908 28408 5914
rect 28356 5850 28408 5856
rect 27896 5636 27948 5642
rect 27896 5578 27948 5584
rect 27908 4570 27936 5578
rect 27908 4554 28028 4570
rect 27908 4548 28040 4554
rect 27908 4542 27988 4548
rect 27804 4072 27856 4078
rect 27804 4014 27856 4020
rect 27252 3936 27304 3942
rect 27252 3878 27304 3884
rect 26976 3732 27028 3738
rect 26976 3674 27028 3680
rect 26240 3664 26292 3670
rect 26240 3606 26292 3612
rect 27264 3534 27292 3878
rect 27350 3836 27658 3845
rect 27350 3834 27356 3836
rect 27412 3834 27436 3836
rect 27492 3834 27516 3836
rect 27572 3834 27596 3836
rect 27652 3834 27658 3836
rect 27412 3782 27414 3834
rect 27594 3782 27596 3834
rect 27350 3780 27356 3782
rect 27412 3780 27436 3782
rect 27492 3780 27516 3782
rect 27572 3780 27596 3782
rect 27652 3780 27658 3782
rect 27350 3771 27658 3780
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 27908 3466 27936 4542
rect 27988 4490 28040 4496
rect 28448 4480 28500 4486
rect 28448 4422 28500 4428
rect 28460 4282 28488 4422
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 28354 3904 28410 3913
rect 28354 3839 28410 3848
rect 28368 3738 28396 3839
rect 28356 3732 28408 3738
rect 28356 3674 28408 3680
rect 28460 3534 28488 4218
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 26424 3460 26476 3466
rect 26424 3402 26476 3408
rect 27896 3460 27948 3466
rect 27896 3402 27948 3408
rect 26148 3392 26200 3398
rect 26200 3340 26280 3346
rect 26148 3334 26280 3340
rect 26160 3318 26280 3334
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 22550 2748 22858 2757
rect 22550 2746 22556 2748
rect 22612 2746 22636 2748
rect 22692 2746 22716 2748
rect 22772 2746 22796 2748
rect 22852 2746 22858 2748
rect 22612 2694 22614 2746
rect 22794 2694 22796 2746
rect 22550 2692 22556 2694
rect 22612 2692 22636 2694
rect 22692 2692 22716 2694
rect 22772 2692 22796 2694
rect 22852 2692 22858 2694
rect 22550 2683 22858 2692
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 26252 2446 26280 3318
rect 26436 3126 26464 3402
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 26424 3120 26476 3126
rect 26424 3062 26476 3068
rect 26620 3058 26648 3334
rect 26608 3052 26660 3058
rect 26608 2994 26660 3000
rect 26620 2446 26648 2994
rect 27350 2748 27658 2757
rect 27350 2746 27356 2748
rect 27412 2746 27436 2748
rect 27492 2746 27516 2748
rect 27572 2746 27596 2748
rect 27652 2746 27658 2748
rect 27412 2694 27414 2746
rect 27594 2694 27596 2746
rect 27350 2692 27356 2694
rect 27412 2692 27436 2694
rect 27492 2692 27516 2694
rect 27572 2692 27596 2694
rect 27652 2692 27658 2694
rect 27350 2683 27658 2692
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 5750 2204 6058 2213
rect 5750 2202 5756 2204
rect 5812 2202 5836 2204
rect 5892 2202 5916 2204
rect 5972 2202 5996 2204
rect 6052 2202 6058 2204
rect 5812 2150 5814 2202
rect 5994 2150 5996 2202
rect 5750 2148 5756 2150
rect 5812 2148 5836 2150
rect 5892 2148 5916 2150
rect 5972 2148 5996 2150
rect 6052 2148 6058 2150
rect 5750 2139 6058 2148
rect 10550 2204 10858 2213
rect 10550 2202 10556 2204
rect 10612 2202 10636 2204
rect 10692 2202 10716 2204
rect 10772 2202 10796 2204
rect 10852 2202 10858 2204
rect 10612 2150 10614 2202
rect 10794 2150 10796 2202
rect 10550 2148 10556 2150
rect 10612 2148 10636 2150
rect 10692 2148 10716 2150
rect 10772 2148 10796 2150
rect 10852 2148 10858 2150
rect 10550 2139 10858 2148
rect 11256 800 11284 2382
rect 15350 2204 15658 2213
rect 15350 2202 15356 2204
rect 15412 2202 15436 2204
rect 15492 2202 15516 2204
rect 15572 2202 15596 2204
rect 15652 2202 15658 2204
rect 15412 2150 15414 2202
rect 15594 2150 15596 2202
rect 15350 2148 15356 2150
rect 15412 2148 15436 2150
rect 15492 2148 15516 2150
rect 15572 2148 15596 2150
rect 15652 2148 15658 2150
rect 15350 2139 15658 2148
rect 18708 800 18736 2382
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 20150 2204 20458 2213
rect 20150 2202 20156 2204
rect 20212 2202 20236 2204
rect 20292 2202 20316 2204
rect 20372 2202 20396 2204
rect 20452 2202 20458 2204
rect 20212 2150 20214 2202
rect 20394 2150 20396 2202
rect 20150 2148 20156 2150
rect 20212 2148 20236 2150
rect 20292 2148 20316 2150
rect 20372 2148 20396 2150
rect 20452 2148 20458 2150
rect 20150 2139 20458 2148
rect 24950 2204 25258 2213
rect 24950 2202 24956 2204
rect 25012 2202 25036 2204
rect 25092 2202 25116 2204
rect 25172 2202 25196 2204
rect 25252 2202 25258 2204
rect 25012 2150 25014 2202
rect 25194 2150 25196 2202
rect 24950 2148 24956 2150
rect 25012 2148 25036 2150
rect 25092 2148 25116 2150
rect 25172 2148 25196 2150
rect 25252 2148 25258 2150
rect 24950 2139 25258 2148
rect 26160 800 26188 2246
rect 28368 1465 28396 2246
rect 28354 1456 28410 1465
rect 28354 1391 28410 1400
rect 3790 0 3846 800
rect 11242 0 11298 800
rect 18694 0 18750 800
rect 26146 0 26202 800
<< via2 >>
rect 28354 28328 28410 28384
rect 3356 27770 3412 27772
rect 3436 27770 3492 27772
rect 3516 27770 3572 27772
rect 3596 27770 3652 27772
rect 3356 27718 3402 27770
rect 3402 27718 3412 27770
rect 3436 27718 3466 27770
rect 3466 27718 3478 27770
rect 3478 27718 3492 27770
rect 3516 27718 3530 27770
rect 3530 27718 3542 27770
rect 3542 27718 3572 27770
rect 3596 27718 3606 27770
rect 3606 27718 3652 27770
rect 3356 27716 3412 27718
rect 3436 27716 3492 27718
rect 3516 27716 3572 27718
rect 3596 27716 3652 27718
rect 8156 27770 8212 27772
rect 8236 27770 8292 27772
rect 8316 27770 8372 27772
rect 8396 27770 8452 27772
rect 8156 27718 8202 27770
rect 8202 27718 8212 27770
rect 8236 27718 8266 27770
rect 8266 27718 8278 27770
rect 8278 27718 8292 27770
rect 8316 27718 8330 27770
rect 8330 27718 8342 27770
rect 8342 27718 8372 27770
rect 8396 27718 8406 27770
rect 8406 27718 8452 27770
rect 8156 27716 8212 27718
rect 8236 27716 8292 27718
rect 8316 27716 8372 27718
rect 8396 27716 8452 27718
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 17756 27770 17812 27772
rect 17836 27770 17892 27772
rect 17916 27770 17972 27772
rect 17996 27770 18052 27772
rect 17756 27718 17802 27770
rect 17802 27718 17812 27770
rect 17836 27718 17866 27770
rect 17866 27718 17878 27770
rect 17878 27718 17892 27770
rect 17916 27718 17930 27770
rect 17930 27718 17942 27770
rect 17942 27718 17972 27770
rect 17996 27718 18006 27770
rect 18006 27718 18052 27770
rect 17756 27716 17812 27718
rect 17836 27716 17892 27718
rect 17916 27716 17972 27718
rect 17996 27716 18052 27718
rect 22556 27770 22612 27772
rect 22636 27770 22692 27772
rect 22716 27770 22772 27772
rect 22796 27770 22852 27772
rect 22556 27718 22602 27770
rect 22602 27718 22612 27770
rect 22636 27718 22666 27770
rect 22666 27718 22678 27770
rect 22678 27718 22692 27770
rect 22716 27718 22730 27770
rect 22730 27718 22742 27770
rect 22742 27718 22772 27770
rect 22796 27718 22806 27770
rect 22806 27718 22852 27770
rect 22556 27716 22612 27718
rect 22636 27716 22692 27718
rect 22716 27716 22772 27718
rect 22796 27716 22852 27718
rect 27356 27770 27412 27772
rect 27436 27770 27492 27772
rect 27516 27770 27572 27772
rect 27596 27770 27652 27772
rect 27356 27718 27402 27770
rect 27402 27718 27412 27770
rect 27436 27718 27466 27770
rect 27466 27718 27478 27770
rect 27478 27718 27492 27770
rect 27516 27718 27530 27770
rect 27530 27718 27542 27770
rect 27542 27718 27572 27770
rect 27596 27718 27606 27770
rect 27606 27718 27652 27770
rect 27356 27716 27412 27718
rect 27436 27716 27492 27718
rect 27516 27716 27572 27718
rect 27596 27716 27652 27718
rect 1582 27104 1638 27160
rect 1582 22208 1638 22264
rect 5756 27226 5812 27228
rect 5836 27226 5892 27228
rect 5916 27226 5972 27228
rect 5996 27226 6052 27228
rect 5756 27174 5802 27226
rect 5802 27174 5812 27226
rect 5836 27174 5866 27226
rect 5866 27174 5878 27226
rect 5878 27174 5892 27226
rect 5916 27174 5930 27226
rect 5930 27174 5942 27226
rect 5942 27174 5972 27226
rect 5996 27174 6006 27226
rect 6006 27174 6052 27226
rect 5756 27172 5812 27174
rect 5836 27172 5892 27174
rect 5916 27172 5972 27174
rect 5996 27172 6052 27174
rect 10556 27226 10612 27228
rect 10636 27226 10692 27228
rect 10716 27226 10772 27228
rect 10796 27226 10852 27228
rect 10556 27174 10602 27226
rect 10602 27174 10612 27226
rect 10636 27174 10666 27226
rect 10666 27174 10678 27226
rect 10678 27174 10692 27226
rect 10716 27174 10730 27226
rect 10730 27174 10742 27226
rect 10742 27174 10772 27226
rect 10796 27174 10806 27226
rect 10806 27174 10852 27226
rect 10556 27172 10612 27174
rect 10636 27172 10692 27174
rect 10716 27172 10772 27174
rect 10796 27172 10852 27174
rect 15356 27226 15412 27228
rect 15436 27226 15492 27228
rect 15516 27226 15572 27228
rect 15596 27226 15652 27228
rect 15356 27174 15402 27226
rect 15402 27174 15412 27226
rect 15436 27174 15466 27226
rect 15466 27174 15478 27226
rect 15478 27174 15492 27226
rect 15516 27174 15530 27226
rect 15530 27174 15542 27226
rect 15542 27174 15572 27226
rect 15596 27174 15606 27226
rect 15606 27174 15652 27226
rect 15356 27172 15412 27174
rect 15436 27172 15492 27174
rect 15516 27172 15572 27174
rect 15596 27172 15652 27174
rect 20156 27226 20212 27228
rect 20236 27226 20292 27228
rect 20316 27226 20372 27228
rect 20396 27226 20452 27228
rect 20156 27174 20202 27226
rect 20202 27174 20212 27226
rect 20236 27174 20266 27226
rect 20266 27174 20278 27226
rect 20278 27174 20292 27226
rect 20316 27174 20330 27226
rect 20330 27174 20342 27226
rect 20342 27174 20372 27226
rect 20396 27174 20406 27226
rect 20406 27174 20452 27226
rect 20156 27172 20212 27174
rect 20236 27172 20292 27174
rect 20316 27172 20372 27174
rect 20396 27172 20452 27174
rect 24956 27226 25012 27228
rect 25036 27226 25092 27228
rect 25116 27226 25172 27228
rect 25196 27226 25252 27228
rect 24956 27174 25002 27226
rect 25002 27174 25012 27226
rect 25036 27174 25066 27226
rect 25066 27174 25078 27226
rect 25078 27174 25092 27226
rect 25116 27174 25130 27226
rect 25130 27174 25142 27226
rect 25142 27174 25172 27226
rect 25196 27174 25206 27226
rect 25206 27174 25252 27226
rect 24956 27172 25012 27174
rect 25036 27172 25092 27174
rect 25116 27172 25172 27174
rect 25196 27172 25252 27174
rect 3356 26682 3412 26684
rect 3436 26682 3492 26684
rect 3516 26682 3572 26684
rect 3596 26682 3652 26684
rect 3356 26630 3402 26682
rect 3402 26630 3412 26682
rect 3436 26630 3466 26682
rect 3466 26630 3478 26682
rect 3478 26630 3492 26682
rect 3516 26630 3530 26682
rect 3530 26630 3542 26682
rect 3542 26630 3572 26682
rect 3596 26630 3606 26682
rect 3606 26630 3652 26682
rect 3356 26628 3412 26630
rect 3436 26628 3492 26630
rect 3516 26628 3572 26630
rect 3596 26628 3652 26630
rect 8156 26682 8212 26684
rect 8236 26682 8292 26684
rect 8316 26682 8372 26684
rect 8396 26682 8452 26684
rect 8156 26630 8202 26682
rect 8202 26630 8212 26682
rect 8236 26630 8266 26682
rect 8266 26630 8278 26682
rect 8278 26630 8292 26682
rect 8316 26630 8330 26682
rect 8330 26630 8342 26682
rect 8342 26630 8372 26682
rect 8396 26630 8406 26682
rect 8406 26630 8452 26682
rect 8156 26628 8212 26630
rect 8236 26628 8292 26630
rect 8316 26628 8372 26630
rect 8396 26628 8452 26630
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 17756 26682 17812 26684
rect 17836 26682 17892 26684
rect 17916 26682 17972 26684
rect 17996 26682 18052 26684
rect 17756 26630 17802 26682
rect 17802 26630 17812 26682
rect 17836 26630 17866 26682
rect 17866 26630 17878 26682
rect 17878 26630 17892 26682
rect 17916 26630 17930 26682
rect 17930 26630 17942 26682
rect 17942 26630 17972 26682
rect 17996 26630 18006 26682
rect 18006 26630 18052 26682
rect 17756 26628 17812 26630
rect 17836 26628 17892 26630
rect 17916 26628 17972 26630
rect 17996 26628 18052 26630
rect 22556 26682 22612 26684
rect 22636 26682 22692 26684
rect 22716 26682 22772 26684
rect 22796 26682 22852 26684
rect 22556 26630 22602 26682
rect 22602 26630 22612 26682
rect 22636 26630 22666 26682
rect 22666 26630 22678 26682
rect 22678 26630 22692 26682
rect 22716 26630 22730 26682
rect 22730 26630 22742 26682
rect 22742 26630 22772 26682
rect 22796 26630 22806 26682
rect 22806 26630 22852 26682
rect 22556 26628 22612 26630
rect 22636 26628 22692 26630
rect 22716 26628 22772 26630
rect 22796 26628 22852 26630
rect 27356 26682 27412 26684
rect 27436 26682 27492 26684
rect 27516 26682 27572 26684
rect 27596 26682 27652 26684
rect 27356 26630 27402 26682
rect 27402 26630 27412 26682
rect 27436 26630 27466 26682
rect 27466 26630 27478 26682
rect 27478 26630 27492 26682
rect 27516 26630 27530 26682
rect 27530 26630 27542 26682
rect 27542 26630 27572 26682
rect 27596 26630 27606 26682
rect 27606 26630 27652 26682
rect 27356 26628 27412 26630
rect 27436 26628 27492 26630
rect 27516 26628 27572 26630
rect 27596 26628 27652 26630
rect 5756 26138 5812 26140
rect 5836 26138 5892 26140
rect 5916 26138 5972 26140
rect 5996 26138 6052 26140
rect 5756 26086 5802 26138
rect 5802 26086 5812 26138
rect 5836 26086 5866 26138
rect 5866 26086 5878 26138
rect 5878 26086 5892 26138
rect 5916 26086 5930 26138
rect 5930 26086 5942 26138
rect 5942 26086 5972 26138
rect 5996 26086 6006 26138
rect 6006 26086 6052 26138
rect 5756 26084 5812 26086
rect 5836 26084 5892 26086
rect 5916 26084 5972 26086
rect 5996 26084 6052 26086
rect 10556 26138 10612 26140
rect 10636 26138 10692 26140
rect 10716 26138 10772 26140
rect 10796 26138 10852 26140
rect 10556 26086 10602 26138
rect 10602 26086 10612 26138
rect 10636 26086 10666 26138
rect 10666 26086 10678 26138
rect 10678 26086 10692 26138
rect 10716 26086 10730 26138
rect 10730 26086 10742 26138
rect 10742 26086 10772 26138
rect 10796 26086 10806 26138
rect 10806 26086 10852 26138
rect 10556 26084 10612 26086
rect 10636 26084 10692 26086
rect 10716 26084 10772 26086
rect 10796 26084 10852 26086
rect 15356 26138 15412 26140
rect 15436 26138 15492 26140
rect 15516 26138 15572 26140
rect 15596 26138 15652 26140
rect 15356 26086 15402 26138
rect 15402 26086 15412 26138
rect 15436 26086 15466 26138
rect 15466 26086 15478 26138
rect 15478 26086 15492 26138
rect 15516 26086 15530 26138
rect 15530 26086 15542 26138
rect 15542 26086 15572 26138
rect 15596 26086 15606 26138
rect 15606 26086 15652 26138
rect 15356 26084 15412 26086
rect 15436 26084 15492 26086
rect 15516 26084 15572 26086
rect 15596 26084 15652 26086
rect 20156 26138 20212 26140
rect 20236 26138 20292 26140
rect 20316 26138 20372 26140
rect 20396 26138 20452 26140
rect 20156 26086 20202 26138
rect 20202 26086 20212 26138
rect 20236 26086 20266 26138
rect 20266 26086 20278 26138
rect 20278 26086 20292 26138
rect 20316 26086 20330 26138
rect 20330 26086 20342 26138
rect 20342 26086 20372 26138
rect 20396 26086 20406 26138
rect 20406 26086 20452 26138
rect 20156 26084 20212 26086
rect 20236 26084 20292 26086
rect 20316 26084 20372 26086
rect 20396 26084 20452 26086
rect 24956 26138 25012 26140
rect 25036 26138 25092 26140
rect 25116 26138 25172 26140
rect 25196 26138 25252 26140
rect 24956 26086 25002 26138
rect 25002 26086 25012 26138
rect 25036 26086 25066 26138
rect 25066 26086 25078 26138
rect 25078 26086 25092 26138
rect 25116 26086 25130 26138
rect 25130 26086 25142 26138
rect 25142 26086 25172 26138
rect 25196 26086 25206 26138
rect 25206 26086 25252 26138
rect 24956 26084 25012 26086
rect 25036 26084 25092 26086
rect 25116 26084 25172 26086
rect 25196 26084 25252 26086
rect 3356 25594 3412 25596
rect 3436 25594 3492 25596
rect 3516 25594 3572 25596
rect 3596 25594 3652 25596
rect 3356 25542 3402 25594
rect 3402 25542 3412 25594
rect 3436 25542 3466 25594
rect 3466 25542 3478 25594
rect 3478 25542 3492 25594
rect 3516 25542 3530 25594
rect 3530 25542 3542 25594
rect 3542 25542 3572 25594
rect 3596 25542 3606 25594
rect 3606 25542 3652 25594
rect 3356 25540 3412 25542
rect 3436 25540 3492 25542
rect 3516 25540 3572 25542
rect 3596 25540 3652 25542
rect 8156 25594 8212 25596
rect 8236 25594 8292 25596
rect 8316 25594 8372 25596
rect 8396 25594 8452 25596
rect 8156 25542 8202 25594
rect 8202 25542 8212 25594
rect 8236 25542 8266 25594
rect 8266 25542 8278 25594
rect 8278 25542 8292 25594
rect 8316 25542 8330 25594
rect 8330 25542 8342 25594
rect 8342 25542 8372 25594
rect 8396 25542 8406 25594
rect 8406 25542 8452 25594
rect 8156 25540 8212 25542
rect 8236 25540 8292 25542
rect 8316 25540 8372 25542
rect 8396 25540 8452 25542
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 17756 25594 17812 25596
rect 17836 25594 17892 25596
rect 17916 25594 17972 25596
rect 17996 25594 18052 25596
rect 17756 25542 17802 25594
rect 17802 25542 17812 25594
rect 17836 25542 17866 25594
rect 17866 25542 17878 25594
rect 17878 25542 17892 25594
rect 17916 25542 17930 25594
rect 17930 25542 17942 25594
rect 17942 25542 17972 25594
rect 17996 25542 18006 25594
rect 18006 25542 18052 25594
rect 17756 25540 17812 25542
rect 17836 25540 17892 25542
rect 17916 25540 17972 25542
rect 17996 25540 18052 25542
rect 22556 25594 22612 25596
rect 22636 25594 22692 25596
rect 22716 25594 22772 25596
rect 22796 25594 22852 25596
rect 22556 25542 22602 25594
rect 22602 25542 22612 25594
rect 22636 25542 22666 25594
rect 22666 25542 22678 25594
rect 22678 25542 22692 25594
rect 22716 25542 22730 25594
rect 22730 25542 22742 25594
rect 22742 25542 22772 25594
rect 22796 25542 22806 25594
rect 22806 25542 22852 25594
rect 22556 25540 22612 25542
rect 22636 25540 22692 25542
rect 22716 25540 22772 25542
rect 22796 25540 22852 25542
rect 27356 25594 27412 25596
rect 27436 25594 27492 25596
rect 27516 25594 27572 25596
rect 27596 25594 27652 25596
rect 27356 25542 27402 25594
rect 27402 25542 27412 25594
rect 27436 25542 27466 25594
rect 27466 25542 27478 25594
rect 27478 25542 27492 25594
rect 27516 25542 27530 25594
rect 27530 25542 27542 25594
rect 27542 25542 27572 25594
rect 27596 25542 27606 25594
rect 27606 25542 27652 25594
rect 27356 25540 27412 25542
rect 27436 25540 27492 25542
rect 27516 25540 27572 25542
rect 27596 25540 27652 25542
rect 5756 25050 5812 25052
rect 5836 25050 5892 25052
rect 5916 25050 5972 25052
rect 5996 25050 6052 25052
rect 5756 24998 5802 25050
rect 5802 24998 5812 25050
rect 5836 24998 5866 25050
rect 5866 24998 5878 25050
rect 5878 24998 5892 25050
rect 5916 24998 5930 25050
rect 5930 24998 5942 25050
rect 5942 24998 5972 25050
rect 5996 24998 6006 25050
rect 6006 24998 6052 25050
rect 5756 24996 5812 24998
rect 5836 24996 5892 24998
rect 5916 24996 5972 24998
rect 5996 24996 6052 24998
rect 10556 25050 10612 25052
rect 10636 25050 10692 25052
rect 10716 25050 10772 25052
rect 10796 25050 10852 25052
rect 10556 24998 10602 25050
rect 10602 24998 10612 25050
rect 10636 24998 10666 25050
rect 10666 24998 10678 25050
rect 10678 24998 10692 25050
rect 10716 24998 10730 25050
rect 10730 24998 10742 25050
rect 10742 24998 10772 25050
rect 10796 24998 10806 25050
rect 10806 24998 10852 25050
rect 10556 24996 10612 24998
rect 10636 24996 10692 24998
rect 10716 24996 10772 24998
rect 10796 24996 10852 24998
rect 15356 25050 15412 25052
rect 15436 25050 15492 25052
rect 15516 25050 15572 25052
rect 15596 25050 15652 25052
rect 15356 24998 15402 25050
rect 15402 24998 15412 25050
rect 15436 24998 15466 25050
rect 15466 24998 15478 25050
rect 15478 24998 15492 25050
rect 15516 24998 15530 25050
rect 15530 24998 15542 25050
rect 15542 24998 15572 25050
rect 15596 24998 15606 25050
rect 15606 24998 15652 25050
rect 15356 24996 15412 24998
rect 15436 24996 15492 24998
rect 15516 24996 15572 24998
rect 15596 24996 15652 24998
rect 20156 25050 20212 25052
rect 20236 25050 20292 25052
rect 20316 25050 20372 25052
rect 20396 25050 20452 25052
rect 20156 24998 20202 25050
rect 20202 24998 20212 25050
rect 20236 24998 20266 25050
rect 20266 24998 20278 25050
rect 20278 24998 20292 25050
rect 20316 24998 20330 25050
rect 20330 24998 20342 25050
rect 20342 24998 20372 25050
rect 20396 24998 20406 25050
rect 20406 24998 20452 25050
rect 20156 24996 20212 24998
rect 20236 24996 20292 24998
rect 20316 24996 20372 24998
rect 20396 24996 20452 24998
rect 24956 25050 25012 25052
rect 25036 25050 25092 25052
rect 25116 25050 25172 25052
rect 25196 25050 25252 25052
rect 24956 24998 25002 25050
rect 25002 24998 25012 25050
rect 25036 24998 25066 25050
rect 25066 24998 25078 25050
rect 25078 24998 25092 25050
rect 25116 24998 25130 25050
rect 25130 24998 25142 25050
rect 25142 24998 25172 25050
rect 25196 24998 25206 25050
rect 25206 24998 25252 25050
rect 24956 24996 25012 24998
rect 25036 24996 25092 24998
rect 25116 24996 25172 24998
rect 25196 24996 25252 24998
rect 3356 24506 3412 24508
rect 3436 24506 3492 24508
rect 3516 24506 3572 24508
rect 3596 24506 3652 24508
rect 3356 24454 3402 24506
rect 3402 24454 3412 24506
rect 3436 24454 3466 24506
rect 3466 24454 3478 24506
rect 3478 24454 3492 24506
rect 3516 24454 3530 24506
rect 3530 24454 3542 24506
rect 3542 24454 3572 24506
rect 3596 24454 3606 24506
rect 3606 24454 3652 24506
rect 3356 24452 3412 24454
rect 3436 24452 3492 24454
rect 3516 24452 3572 24454
rect 3596 24452 3652 24454
rect 8156 24506 8212 24508
rect 8236 24506 8292 24508
rect 8316 24506 8372 24508
rect 8396 24506 8452 24508
rect 8156 24454 8202 24506
rect 8202 24454 8212 24506
rect 8236 24454 8266 24506
rect 8266 24454 8278 24506
rect 8278 24454 8292 24506
rect 8316 24454 8330 24506
rect 8330 24454 8342 24506
rect 8342 24454 8372 24506
rect 8396 24454 8406 24506
rect 8406 24454 8452 24506
rect 8156 24452 8212 24454
rect 8236 24452 8292 24454
rect 8316 24452 8372 24454
rect 8396 24452 8452 24454
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 17756 24506 17812 24508
rect 17836 24506 17892 24508
rect 17916 24506 17972 24508
rect 17996 24506 18052 24508
rect 17756 24454 17802 24506
rect 17802 24454 17812 24506
rect 17836 24454 17866 24506
rect 17866 24454 17878 24506
rect 17878 24454 17892 24506
rect 17916 24454 17930 24506
rect 17930 24454 17942 24506
rect 17942 24454 17972 24506
rect 17996 24454 18006 24506
rect 18006 24454 18052 24506
rect 17756 24452 17812 24454
rect 17836 24452 17892 24454
rect 17916 24452 17972 24454
rect 17996 24452 18052 24454
rect 22556 24506 22612 24508
rect 22636 24506 22692 24508
rect 22716 24506 22772 24508
rect 22796 24506 22852 24508
rect 22556 24454 22602 24506
rect 22602 24454 22612 24506
rect 22636 24454 22666 24506
rect 22666 24454 22678 24506
rect 22678 24454 22692 24506
rect 22716 24454 22730 24506
rect 22730 24454 22742 24506
rect 22742 24454 22772 24506
rect 22796 24454 22806 24506
rect 22806 24454 22852 24506
rect 22556 24452 22612 24454
rect 22636 24452 22692 24454
rect 22716 24452 22772 24454
rect 22796 24452 22852 24454
rect 27356 24506 27412 24508
rect 27436 24506 27492 24508
rect 27516 24506 27572 24508
rect 27596 24506 27652 24508
rect 27356 24454 27402 24506
rect 27402 24454 27412 24506
rect 27436 24454 27466 24506
rect 27466 24454 27478 24506
rect 27478 24454 27492 24506
rect 27516 24454 27530 24506
rect 27530 24454 27542 24506
rect 27542 24454 27572 24506
rect 27596 24454 27606 24506
rect 27606 24454 27652 24506
rect 27356 24452 27412 24454
rect 27436 24452 27492 24454
rect 27516 24452 27572 24454
rect 27596 24452 27652 24454
rect 5756 23962 5812 23964
rect 5836 23962 5892 23964
rect 5916 23962 5972 23964
rect 5996 23962 6052 23964
rect 5756 23910 5802 23962
rect 5802 23910 5812 23962
rect 5836 23910 5866 23962
rect 5866 23910 5878 23962
rect 5878 23910 5892 23962
rect 5916 23910 5930 23962
rect 5930 23910 5942 23962
rect 5942 23910 5972 23962
rect 5996 23910 6006 23962
rect 6006 23910 6052 23962
rect 5756 23908 5812 23910
rect 5836 23908 5892 23910
rect 5916 23908 5972 23910
rect 5996 23908 6052 23910
rect 10556 23962 10612 23964
rect 10636 23962 10692 23964
rect 10716 23962 10772 23964
rect 10796 23962 10852 23964
rect 10556 23910 10602 23962
rect 10602 23910 10612 23962
rect 10636 23910 10666 23962
rect 10666 23910 10678 23962
rect 10678 23910 10692 23962
rect 10716 23910 10730 23962
rect 10730 23910 10742 23962
rect 10742 23910 10772 23962
rect 10796 23910 10806 23962
rect 10806 23910 10852 23962
rect 10556 23908 10612 23910
rect 10636 23908 10692 23910
rect 10716 23908 10772 23910
rect 10796 23908 10852 23910
rect 15356 23962 15412 23964
rect 15436 23962 15492 23964
rect 15516 23962 15572 23964
rect 15596 23962 15652 23964
rect 15356 23910 15402 23962
rect 15402 23910 15412 23962
rect 15436 23910 15466 23962
rect 15466 23910 15478 23962
rect 15478 23910 15492 23962
rect 15516 23910 15530 23962
rect 15530 23910 15542 23962
rect 15542 23910 15572 23962
rect 15596 23910 15606 23962
rect 15606 23910 15652 23962
rect 15356 23908 15412 23910
rect 15436 23908 15492 23910
rect 15516 23908 15572 23910
rect 15596 23908 15652 23910
rect 20156 23962 20212 23964
rect 20236 23962 20292 23964
rect 20316 23962 20372 23964
rect 20396 23962 20452 23964
rect 20156 23910 20202 23962
rect 20202 23910 20212 23962
rect 20236 23910 20266 23962
rect 20266 23910 20278 23962
rect 20278 23910 20292 23962
rect 20316 23910 20330 23962
rect 20330 23910 20342 23962
rect 20342 23910 20372 23962
rect 20396 23910 20406 23962
rect 20406 23910 20452 23962
rect 20156 23908 20212 23910
rect 20236 23908 20292 23910
rect 20316 23908 20372 23910
rect 20396 23908 20452 23910
rect 24956 23962 25012 23964
rect 25036 23962 25092 23964
rect 25116 23962 25172 23964
rect 25196 23962 25252 23964
rect 24956 23910 25002 23962
rect 25002 23910 25012 23962
rect 25036 23910 25066 23962
rect 25066 23910 25078 23962
rect 25078 23910 25092 23962
rect 25116 23910 25130 23962
rect 25130 23910 25142 23962
rect 25142 23910 25172 23962
rect 25196 23910 25206 23962
rect 25206 23910 25252 23962
rect 24956 23908 25012 23910
rect 25036 23908 25092 23910
rect 25116 23908 25172 23910
rect 25196 23908 25252 23910
rect 3356 23418 3412 23420
rect 3436 23418 3492 23420
rect 3516 23418 3572 23420
rect 3596 23418 3652 23420
rect 3356 23366 3402 23418
rect 3402 23366 3412 23418
rect 3436 23366 3466 23418
rect 3466 23366 3478 23418
rect 3478 23366 3492 23418
rect 3516 23366 3530 23418
rect 3530 23366 3542 23418
rect 3542 23366 3572 23418
rect 3596 23366 3606 23418
rect 3606 23366 3652 23418
rect 3356 23364 3412 23366
rect 3436 23364 3492 23366
rect 3516 23364 3572 23366
rect 3596 23364 3652 23366
rect 8156 23418 8212 23420
rect 8236 23418 8292 23420
rect 8316 23418 8372 23420
rect 8396 23418 8452 23420
rect 8156 23366 8202 23418
rect 8202 23366 8212 23418
rect 8236 23366 8266 23418
rect 8266 23366 8278 23418
rect 8278 23366 8292 23418
rect 8316 23366 8330 23418
rect 8330 23366 8342 23418
rect 8342 23366 8372 23418
rect 8396 23366 8406 23418
rect 8406 23366 8452 23418
rect 8156 23364 8212 23366
rect 8236 23364 8292 23366
rect 8316 23364 8372 23366
rect 8396 23364 8452 23366
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 17756 23418 17812 23420
rect 17836 23418 17892 23420
rect 17916 23418 17972 23420
rect 17996 23418 18052 23420
rect 17756 23366 17802 23418
rect 17802 23366 17812 23418
rect 17836 23366 17866 23418
rect 17866 23366 17878 23418
rect 17878 23366 17892 23418
rect 17916 23366 17930 23418
rect 17930 23366 17942 23418
rect 17942 23366 17972 23418
rect 17996 23366 18006 23418
rect 18006 23366 18052 23418
rect 17756 23364 17812 23366
rect 17836 23364 17892 23366
rect 17916 23364 17972 23366
rect 17996 23364 18052 23366
rect 22556 23418 22612 23420
rect 22636 23418 22692 23420
rect 22716 23418 22772 23420
rect 22796 23418 22852 23420
rect 22556 23366 22602 23418
rect 22602 23366 22612 23418
rect 22636 23366 22666 23418
rect 22666 23366 22678 23418
rect 22678 23366 22692 23418
rect 22716 23366 22730 23418
rect 22730 23366 22742 23418
rect 22742 23366 22772 23418
rect 22796 23366 22806 23418
rect 22806 23366 22852 23418
rect 22556 23364 22612 23366
rect 22636 23364 22692 23366
rect 22716 23364 22772 23366
rect 22796 23364 22852 23366
rect 5756 22874 5812 22876
rect 5836 22874 5892 22876
rect 5916 22874 5972 22876
rect 5996 22874 6052 22876
rect 5756 22822 5802 22874
rect 5802 22822 5812 22874
rect 5836 22822 5866 22874
rect 5866 22822 5878 22874
rect 5878 22822 5892 22874
rect 5916 22822 5930 22874
rect 5930 22822 5942 22874
rect 5942 22822 5972 22874
rect 5996 22822 6006 22874
rect 6006 22822 6052 22874
rect 5756 22820 5812 22822
rect 5836 22820 5892 22822
rect 5916 22820 5972 22822
rect 5996 22820 6052 22822
rect 10556 22874 10612 22876
rect 10636 22874 10692 22876
rect 10716 22874 10772 22876
rect 10796 22874 10852 22876
rect 10556 22822 10602 22874
rect 10602 22822 10612 22874
rect 10636 22822 10666 22874
rect 10666 22822 10678 22874
rect 10678 22822 10692 22874
rect 10716 22822 10730 22874
rect 10730 22822 10742 22874
rect 10742 22822 10772 22874
rect 10796 22822 10806 22874
rect 10806 22822 10852 22874
rect 10556 22820 10612 22822
rect 10636 22820 10692 22822
rect 10716 22820 10772 22822
rect 10796 22820 10852 22822
rect 15356 22874 15412 22876
rect 15436 22874 15492 22876
rect 15516 22874 15572 22876
rect 15596 22874 15652 22876
rect 15356 22822 15402 22874
rect 15402 22822 15412 22874
rect 15436 22822 15466 22874
rect 15466 22822 15478 22874
rect 15478 22822 15492 22874
rect 15516 22822 15530 22874
rect 15530 22822 15542 22874
rect 15542 22822 15572 22874
rect 15596 22822 15606 22874
rect 15606 22822 15652 22874
rect 15356 22820 15412 22822
rect 15436 22820 15492 22822
rect 15516 22820 15572 22822
rect 15596 22820 15652 22822
rect 20156 22874 20212 22876
rect 20236 22874 20292 22876
rect 20316 22874 20372 22876
rect 20396 22874 20452 22876
rect 20156 22822 20202 22874
rect 20202 22822 20212 22874
rect 20236 22822 20266 22874
rect 20266 22822 20278 22874
rect 20278 22822 20292 22874
rect 20316 22822 20330 22874
rect 20330 22822 20342 22874
rect 20342 22822 20372 22874
rect 20396 22822 20406 22874
rect 20406 22822 20452 22874
rect 20156 22820 20212 22822
rect 20236 22820 20292 22822
rect 20316 22820 20372 22822
rect 20396 22820 20452 22822
rect 27356 23418 27412 23420
rect 27436 23418 27492 23420
rect 27516 23418 27572 23420
rect 27596 23418 27652 23420
rect 27356 23366 27402 23418
rect 27402 23366 27412 23418
rect 27436 23366 27466 23418
rect 27466 23366 27478 23418
rect 27478 23366 27492 23418
rect 27516 23366 27530 23418
rect 27530 23366 27542 23418
rect 27542 23366 27572 23418
rect 27596 23366 27606 23418
rect 27606 23366 27652 23418
rect 27356 23364 27412 23366
rect 27436 23364 27492 23366
rect 27516 23364 27572 23366
rect 27596 23364 27652 23366
rect 24956 22874 25012 22876
rect 25036 22874 25092 22876
rect 25116 22874 25172 22876
rect 25196 22874 25252 22876
rect 24956 22822 25002 22874
rect 25002 22822 25012 22874
rect 25036 22822 25066 22874
rect 25066 22822 25078 22874
rect 25078 22822 25092 22874
rect 25116 22822 25130 22874
rect 25130 22822 25142 22874
rect 25142 22822 25172 22874
rect 25196 22822 25206 22874
rect 25206 22822 25252 22874
rect 24956 22820 25012 22822
rect 25036 22820 25092 22822
rect 25116 22820 25172 22822
rect 25196 22820 25252 22822
rect 3356 22330 3412 22332
rect 3436 22330 3492 22332
rect 3516 22330 3572 22332
rect 3596 22330 3652 22332
rect 3356 22278 3402 22330
rect 3402 22278 3412 22330
rect 3436 22278 3466 22330
rect 3466 22278 3478 22330
rect 3478 22278 3492 22330
rect 3516 22278 3530 22330
rect 3530 22278 3542 22330
rect 3542 22278 3572 22330
rect 3596 22278 3606 22330
rect 3606 22278 3652 22330
rect 3356 22276 3412 22278
rect 3436 22276 3492 22278
rect 3516 22276 3572 22278
rect 3596 22276 3652 22278
rect 8156 22330 8212 22332
rect 8236 22330 8292 22332
rect 8316 22330 8372 22332
rect 8396 22330 8452 22332
rect 8156 22278 8202 22330
rect 8202 22278 8212 22330
rect 8236 22278 8266 22330
rect 8266 22278 8278 22330
rect 8278 22278 8292 22330
rect 8316 22278 8330 22330
rect 8330 22278 8342 22330
rect 8342 22278 8372 22330
rect 8396 22278 8406 22330
rect 8406 22278 8452 22330
rect 8156 22276 8212 22278
rect 8236 22276 8292 22278
rect 8316 22276 8372 22278
rect 8396 22276 8452 22278
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 17756 22330 17812 22332
rect 17836 22330 17892 22332
rect 17916 22330 17972 22332
rect 17996 22330 18052 22332
rect 17756 22278 17802 22330
rect 17802 22278 17812 22330
rect 17836 22278 17866 22330
rect 17866 22278 17878 22330
rect 17878 22278 17892 22330
rect 17916 22278 17930 22330
rect 17930 22278 17942 22330
rect 17942 22278 17972 22330
rect 17996 22278 18006 22330
rect 18006 22278 18052 22330
rect 17756 22276 17812 22278
rect 17836 22276 17892 22278
rect 17916 22276 17972 22278
rect 17996 22276 18052 22278
rect 22556 22330 22612 22332
rect 22636 22330 22692 22332
rect 22716 22330 22772 22332
rect 22796 22330 22852 22332
rect 22556 22278 22602 22330
rect 22602 22278 22612 22330
rect 22636 22278 22666 22330
rect 22666 22278 22678 22330
rect 22678 22278 22692 22330
rect 22716 22278 22730 22330
rect 22730 22278 22742 22330
rect 22742 22278 22772 22330
rect 22796 22278 22806 22330
rect 22806 22278 22852 22330
rect 22556 22276 22612 22278
rect 22636 22276 22692 22278
rect 22716 22276 22772 22278
rect 22796 22276 22852 22278
rect 5756 21786 5812 21788
rect 5836 21786 5892 21788
rect 5916 21786 5972 21788
rect 5996 21786 6052 21788
rect 5756 21734 5802 21786
rect 5802 21734 5812 21786
rect 5836 21734 5866 21786
rect 5866 21734 5878 21786
rect 5878 21734 5892 21786
rect 5916 21734 5930 21786
rect 5930 21734 5942 21786
rect 5942 21734 5972 21786
rect 5996 21734 6006 21786
rect 6006 21734 6052 21786
rect 5756 21732 5812 21734
rect 5836 21732 5892 21734
rect 5916 21732 5972 21734
rect 5996 21732 6052 21734
rect 10556 21786 10612 21788
rect 10636 21786 10692 21788
rect 10716 21786 10772 21788
rect 10796 21786 10852 21788
rect 10556 21734 10602 21786
rect 10602 21734 10612 21786
rect 10636 21734 10666 21786
rect 10666 21734 10678 21786
rect 10678 21734 10692 21786
rect 10716 21734 10730 21786
rect 10730 21734 10742 21786
rect 10742 21734 10772 21786
rect 10796 21734 10806 21786
rect 10806 21734 10852 21786
rect 10556 21732 10612 21734
rect 10636 21732 10692 21734
rect 10716 21732 10772 21734
rect 10796 21732 10852 21734
rect 15356 21786 15412 21788
rect 15436 21786 15492 21788
rect 15516 21786 15572 21788
rect 15596 21786 15652 21788
rect 15356 21734 15402 21786
rect 15402 21734 15412 21786
rect 15436 21734 15466 21786
rect 15466 21734 15478 21786
rect 15478 21734 15492 21786
rect 15516 21734 15530 21786
rect 15530 21734 15542 21786
rect 15542 21734 15572 21786
rect 15596 21734 15606 21786
rect 15606 21734 15652 21786
rect 15356 21732 15412 21734
rect 15436 21732 15492 21734
rect 15516 21732 15572 21734
rect 15596 21732 15652 21734
rect 3356 21242 3412 21244
rect 3436 21242 3492 21244
rect 3516 21242 3572 21244
rect 3596 21242 3652 21244
rect 3356 21190 3402 21242
rect 3402 21190 3412 21242
rect 3436 21190 3466 21242
rect 3466 21190 3478 21242
rect 3478 21190 3492 21242
rect 3516 21190 3530 21242
rect 3530 21190 3542 21242
rect 3542 21190 3572 21242
rect 3596 21190 3606 21242
rect 3606 21190 3652 21242
rect 3356 21188 3412 21190
rect 3436 21188 3492 21190
rect 3516 21188 3572 21190
rect 3596 21188 3652 21190
rect 8156 21242 8212 21244
rect 8236 21242 8292 21244
rect 8316 21242 8372 21244
rect 8396 21242 8452 21244
rect 8156 21190 8202 21242
rect 8202 21190 8212 21242
rect 8236 21190 8266 21242
rect 8266 21190 8278 21242
rect 8278 21190 8292 21242
rect 8316 21190 8330 21242
rect 8330 21190 8342 21242
rect 8342 21190 8372 21242
rect 8396 21190 8406 21242
rect 8406 21190 8452 21242
rect 8156 21188 8212 21190
rect 8236 21188 8292 21190
rect 8316 21188 8372 21190
rect 8396 21188 8452 21190
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 17756 21242 17812 21244
rect 17836 21242 17892 21244
rect 17916 21242 17972 21244
rect 17996 21242 18052 21244
rect 17756 21190 17802 21242
rect 17802 21190 17812 21242
rect 17836 21190 17866 21242
rect 17866 21190 17878 21242
rect 17878 21190 17892 21242
rect 17916 21190 17930 21242
rect 17930 21190 17942 21242
rect 17942 21190 17972 21242
rect 17996 21190 18006 21242
rect 18006 21190 18052 21242
rect 17756 21188 17812 21190
rect 17836 21188 17892 21190
rect 17916 21188 17972 21190
rect 17996 21188 18052 21190
rect 3356 20154 3412 20156
rect 3436 20154 3492 20156
rect 3516 20154 3572 20156
rect 3596 20154 3652 20156
rect 3356 20102 3402 20154
rect 3402 20102 3412 20154
rect 3436 20102 3466 20154
rect 3466 20102 3478 20154
rect 3478 20102 3492 20154
rect 3516 20102 3530 20154
rect 3530 20102 3542 20154
rect 3542 20102 3572 20154
rect 3596 20102 3606 20154
rect 3606 20102 3652 20154
rect 3356 20100 3412 20102
rect 3436 20100 3492 20102
rect 3516 20100 3572 20102
rect 3596 20100 3652 20102
rect 3356 19066 3412 19068
rect 3436 19066 3492 19068
rect 3516 19066 3572 19068
rect 3596 19066 3652 19068
rect 3356 19014 3402 19066
rect 3402 19014 3412 19066
rect 3436 19014 3466 19066
rect 3466 19014 3478 19066
rect 3478 19014 3492 19066
rect 3516 19014 3530 19066
rect 3530 19014 3542 19066
rect 3542 19014 3572 19066
rect 3596 19014 3606 19066
rect 3606 19014 3652 19066
rect 3356 19012 3412 19014
rect 3436 19012 3492 19014
rect 3516 19012 3572 19014
rect 3596 19012 3652 19014
rect 1582 17332 1638 17368
rect 3356 17978 3412 17980
rect 3436 17978 3492 17980
rect 3516 17978 3572 17980
rect 3596 17978 3652 17980
rect 3356 17926 3402 17978
rect 3402 17926 3412 17978
rect 3436 17926 3466 17978
rect 3466 17926 3478 17978
rect 3478 17926 3492 17978
rect 3516 17926 3530 17978
rect 3530 17926 3542 17978
rect 3542 17926 3572 17978
rect 3596 17926 3606 17978
rect 3606 17926 3652 17978
rect 3356 17924 3412 17926
rect 3436 17924 3492 17926
rect 3516 17924 3572 17926
rect 3596 17924 3652 17926
rect 1582 17312 1584 17332
rect 1584 17312 1636 17332
rect 1636 17312 1638 17332
rect 5756 20698 5812 20700
rect 5836 20698 5892 20700
rect 5916 20698 5972 20700
rect 5996 20698 6052 20700
rect 5756 20646 5802 20698
rect 5802 20646 5812 20698
rect 5836 20646 5866 20698
rect 5866 20646 5878 20698
rect 5878 20646 5892 20698
rect 5916 20646 5930 20698
rect 5930 20646 5942 20698
rect 5942 20646 5972 20698
rect 5996 20646 6006 20698
rect 6006 20646 6052 20698
rect 5756 20644 5812 20646
rect 5836 20644 5892 20646
rect 5916 20644 5972 20646
rect 5996 20644 6052 20646
rect 5756 19610 5812 19612
rect 5836 19610 5892 19612
rect 5916 19610 5972 19612
rect 5996 19610 6052 19612
rect 5756 19558 5802 19610
rect 5802 19558 5812 19610
rect 5836 19558 5866 19610
rect 5866 19558 5878 19610
rect 5878 19558 5892 19610
rect 5916 19558 5930 19610
rect 5930 19558 5942 19610
rect 5942 19558 5972 19610
rect 5996 19558 6006 19610
rect 6006 19558 6052 19610
rect 5756 19556 5812 19558
rect 5836 19556 5892 19558
rect 5916 19556 5972 19558
rect 5996 19556 6052 19558
rect 10556 20698 10612 20700
rect 10636 20698 10692 20700
rect 10716 20698 10772 20700
rect 10796 20698 10852 20700
rect 10556 20646 10602 20698
rect 10602 20646 10612 20698
rect 10636 20646 10666 20698
rect 10666 20646 10678 20698
rect 10678 20646 10692 20698
rect 10716 20646 10730 20698
rect 10730 20646 10742 20698
rect 10742 20646 10772 20698
rect 10796 20646 10806 20698
rect 10806 20646 10852 20698
rect 10556 20644 10612 20646
rect 10636 20644 10692 20646
rect 10716 20644 10772 20646
rect 10796 20644 10852 20646
rect 15356 20698 15412 20700
rect 15436 20698 15492 20700
rect 15516 20698 15572 20700
rect 15596 20698 15652 20700
rect 15356 20646 15402 20698
rect 15402 20646 15412 20698
rect 15436 20646 15466 20698
rect 15466 20646 15478 20698
rect 15478 20646 15492 20698
rect 15516 20646 15530 20698
rect 15530 20646 15542 20698
rect 15542 20646 15572 20698
rect 15596 20646 15606 20698
rect 15606 20646 15652 20698
rect 15356 20644 15412 20646
rect 15436 20644 15492 20646
rect 15516 20644 15572 20646
rect 15596 20644 15652 20646
rect 8156 20154 8212 20156
rect 8236 20154 8292 20156
rect 8316 20154 8372 20156
rect 8396 20154 8452 20156
rect 8156 20102 8202 20154
rect 8202 20102 8212 20154
rect 8236 20102 8266 20154
rect 8266 20102 8278 20154
rect 8278 20102 8292 20154
rect 8316 20102 8330 20154
rect 8330 20102 8342 20154
rect 8342 20102 8372 20154
rect 8396 20102 8406 20154
rect 8406 20102 8452 20154
rect 8156 20100 8212 20102
rect 8236 20100 8292 20102
rect 8316 20100 8372 20102
rect 8396 20100 8452 20102
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 10556 19610 10612 19612
rect 10636 19610 10692 19612
rect 10716 19610 10772 19612
rect 10796 19610 10852 19612
rect 10556 19558 10602 19610
rect 10602 19558 10612 19610
rect 10636 19558 10666 19610
rect 10666 19558 10678 19610
rect 10678 19558 10692 19610
rect 10716 19558 10730 19610
rect 10730 19558 10742 19610
rect 10742 19558 10772 19610
rect 10796 19558 10806 19610
rect 10806 19558 10852 19610
rect 10556 19556 10612 19558
rect 10636 19556 10692 19558
rect 10716 19556 10772 19558
rect 10796 19556 10852 19558
rect 15356 19610 15412 19612
rect 15436 19610 15492 19612
rect 15516 19610 15572 19612
rect 15596 19610 15652 19612
rect 15356 19558 15402 19610
rect 15402 19558 15412 19610
rect 15436 19558 15466 19610
rect 15466 19558 15478 19610
rect 15478 19558 15492 19610
rect 15516 19558 15530 19610
rect 15530 19558 15542 19610
rect 15542 19558 15572 19610
rect 15596 19558 15606 19610
rect 15606 19558 15652 19610
rect 15356 19556 15412 19558
rect 15436 19556 15492 19558
rect 15516 19556 15572 19558
rect 15596 19556 15652 19558
rect 17756 20154 17812 20156
rect 17836 20154 17892 20156
rect 17916 20154 17972 20156
rect 17996 20154 18052 20156
rect 17756 20102 17802 20154
rect 17802 20102 17812 20154
rect 17836 20102 17866 20154
rect 17866 20102 17878 20154
rect 17878 20102 17892 20154
rect 17916 20102 17930 20154
rect 17930 20102 17942 20154
rect 17942 20102 17972 20154
rect 17996 20102 18006 20154
rect 18006 20102 18052 20154
rect 17756 20100 17812 20102
rect 17836 20100 17892 20102
rect 17916 20100 17972 20102
rect 17996 20100 18052 20102
rect 8156 19066 8212 19068
rect 8236 19066 8292 19068
rect 8316 19066 8372 19068
rect 8396 19066 8452 19068
rect 8156 19014 8202 19066
rect 8202 19014 8212 19066
rect 8236 19014 8266 19066
rect 8266 19014 8278 19066
rect 8278 19014 8292 19066
rect 8316 19014 8330 19066
rect 8330 19014 8342 19066
rect 8342 19014 8372 19066
rect 8396 19014 8406 19066
rect 8406 19014 8452 19066
rect 8156 19012 8212 19014
rect 8236 19012 8292 19014
rect 8316 19012 8372 19014
rect 8396 19012 8452 19014
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 3356 16890 3412 16892
rect 3436 16890 3492 16892
rect 3516 16890 3572 16892
rect 3596 16890 3652 16892
rect 3356 16838 3402 16890
rect 3402 16838 3412 16890
rect 3436 16838 3466 16890
rect 3466 16838 3478 16890
rect 3478 16838 3492 16890
rect 3516 16838 3530 16890
rect 3530 16838 3542 16890
rect 3542 16838 3572 16890
rect 3596 16838 3606 16890
rect 3606 16838 3652 16890
rect 3356 16836 3412 16838
rect 3436 16836 3492 16838
rect 3516 16836 3572 16838
rect 3596 16836 3652 16838
rect 3356 15802 3412 15804
rect 3436 15802 3492 15804
rect 3516 15802 3572 15804
rect 3596 15802 3652 15804
rect 3356 15750 3402 15802
rect 3402 15750 3412 15802
rect 3436 15750 3466 15802
rect 3466 15750 3478 15802
rect 3478 15750 3492 15802
rect 3516 15750 3530 15802
rect 3530 15750 3542 15802
rect 3542 15750 3572 15802
rect 3596 15750 3606 15802
rect 3606 15750 3652 15802
rect 3356 15748 3412 15750
rect 3436 15748 3492 15750
rect 3516 15748 3572 15750
rect 3596 15748 3652 15750
rect 5756 18522 5812 18524
rect 5836 18522 5892 18524
rect 5916 18522 5972 18524
rect 5996 18522 6052 18524
rect 5756 18470 5802 18522
rect 5802 18470 5812 18522
rect 5836 18470 5866 18522
rect 5866 18470 5878 18522
rect 5878 18470 5892 18522
rect 5916 18470 5930 18522
rect 5930 18470 5942 18522
rect 5942 18470 5972 18522
rect 5996 18470 6006 18522
rect 6006 18470 6052 18522
rect 5756 18468 5812 18470
rect 5836 18468 5892 18470
rect 5916 18468 5972 18470
rect 5996 18468 6052 18470
rect 10556 18522 10612 18524
rect 10636 18522 10692 18524
rect 10716 18522 10772 18524
rect 10796 18522 10852 18524
rect 10556 18470 10602 18522
rect 10602 18470 10612 18522
rect 10636 18470 10666 18522
rect 10666 18470 10678 18522
rect 10678 18470 10692 18522
rect 10716 18470 10730 18522
rect 10730 18470 10742 18522
rect 10742 18470 10772 18522
rect 10796 18470 10806 18522
rect 10806 18470 10852 18522
rect 10556 18468 10612 18470
rect 10636 18468 10692 18470
rect 10716 18468 10772 18470
rect 10796 18468 10852 18470
rect 15356 18522 15412 18524
rect 15436 18522 15492 18524
rect 15516 18522 15572 18524
rect 15596 18522 15652 18524
rect 15356 18470 15402 18522
rect 15402 18470 15412 18522
rect 15436 18470 15466 18522
rect 15466 18470 15478 18522
rect 15478 18470 15492 18522
rect 15516 18470 15530 18522
rect 15530 18470 15542 18522
rect 15542 18470 15572 18522
rect 15596 18470 15606 18522
rect 15606 18470 15652 18522
rect 15356 18468 15412 18470
rect 15436 18468 15492 18470
rect 15516 18468 15572 18470
rect 15596 18468 15652 18470
rect 1490 12436 1546 12472
rect 1490 12416 1492 12436
rect 1492 12416 1544 12436
rect 1544 12416 1546 12436
rect 3356 14714 3412 14716
rect 3436 14714 3492 14716
rect 3516 14714 3572 14716
rect 3596 14714 3652 14716
rect 3356 14662 3402 14714
rect 3402 14662 3412 14714
rect 3436 14662 3466 14714
rect 3466 14662 3478 14714
rect 3478 14662 3492 14714
rect 3516 14662 3530 14714
rect 3530 14662 3542 14714
rect 3542 14662 3572 14714
rect 3596 14662 3606 14714
rect 3606 14662 3652 14714
rect 3356 14660 3412 14662
rect 3436 14660 3492 14662
rect 3516 14660 3572 14662
rect 3596 14660 3652 14662
rect 5756 17434 5812 17436
rect 5836 17434 5892 17436
rect 5916 17434 5972 17436
rect 5996 17434 6052 17436
rect 5756 17382 5802 17434
rect 5802 17382 5812 17434
rect 5836 17382 5866 17434
rect 5866 17382 5878 17434
rect 5878 17382 5892 17434
rect 5916 17382 5930 17434
rect 5930 17382 5942 17434
rect 5942 17382 5972 17434
rect 5996 17382 6006 17434
rect 6006 17382 6052 17434
rect 5756 17380 5812 17382
rect 5836 17380 5892 17382
rect 5916 17380 5972 17382
rect 5996 17380 6052 17382
rect 3356 13626 3412 13628
rect 3436 13626 3492 13628
rect 3516 13626 3572 13628
rect 3596 13626 3652 13628
rect 3356 13574 3402 13626
rect 3402 13574 3412 13626
rect 3436 13574 3466 13626
rect 3466 13574 3478 13626
rect 3478 13574 3492 13626
rect 3516 13574 3530 13626
rect 3530 13574 3542 13626
rect 3542 13574 3572 13626
rect 3596 13574 3606 13626
rect 3606 13574 3652 13626
rect 3356 13572 3412 13574
rect 3436 13572 3492 13574
rect 3516 13572 3572 13574
rect 3596 13572 3652 13574
rect 3356 12538 3412 12540
rect 3436 12538 3492 12540
rect 3516 12538 3572 12540
rect 3596 12538 3652 12540
rect 3356 12486 3402 12538
rect 3402 12486 3412 12538
rect 3436 12486 3466 12538
rect 3466 12486 3478 12538
rect 3478 12486 3492 12538
rect 3516 12486 3530 12538
rect 3530 12486 3542 12538
rect 3542 12486 3572 12538
rect 3596 12486 3606 12538
rect 3606 12486 3652 12538
rect 3356 12484 3412 12486
rect 3436 12484 3492 12486
rect 3516 12484 3572 12486
rect 3596 12484 3652 12486
rect 5756 16346 5812 16348
rect 5836 16346 5892 16348
rect 5916 16346 5972 16348
rect 5996 16346 6052 16348
rect 5756 16294 5802 16346
rect 5802 16294 5812 16346
rect 5836 16294 5866 16346
rect 5866 16294 5878 16346
rect 5878 16294 5892 16346
rect 5916 16294 5930 16346
rect 5930 16294 5942 16346
rect 5942 16294 5972 16346
rect 5996 16294 6006 16346
rect 6006 16294 6052 16346
rect 5756 16292 5812 16294
rect 5836 16292 5892 16294
rect 5916 16292 5972 16294
rect 5996 16292 6052 16294
rect 5756 15258 5812 15260
rect 5836 15258 5892 15260
rect 5916 15258 5972 15260
rect 5996 15258 6052 15260
rect 5756 15206 5802 15258
rect 5802 15206 5812 15258
rect 5836 15206 5866 15258
rect 5866 15206 5878 15258
rect 5878 15206 5892 15258
rect 5916 15206 5930 15258
rect 5930 15206 5942 15258
rect 5942 15206 5972 15258
rect 5996 15206 6006 15258
rect 6006 15206 6052 15258
rect 5756 15204 5812 15206
rect 5836 15204 5892 15206
rect 5916 15204 5972 15206
rect 5996 15204 6052 15206
rect 8156 17978 8212 17980
rect 8236 17978 8292 17980
rect 8316 17978 8372 17980
rect 8396 17978 8452 17980
rect 8156 17926 8202 17978
rect 8202 17926 8212 17978
rect 8236 17926 8266 17978
rect 8266 17926 8278 17978
rect 8278 17926 8292 17978
rect 8316 17926 8330 17978
rect 8330 17926 8342 17978
rect 8342 17926 8372 17978
rect 8396 17926 8406 17978
rect 8406 17926 8452 17978
rect 8156 17924 8212 17926
rect 8236 17924 8292 17926
rect 8316 17924 8372 17926
rect 8396 17924 8452 17926
rect 8156 16890 8212 16892
rect 8236 16890 8292 16892
rect 8316 16890 8372 16892
rect 8396 16890 8452 16892
rect 8156 16838 8202 16890
rect 8202 16838 8212 16890
rect 8236 16838 8266 16890
rect 8266 16838 8278 16890
rect 8278 16838 8292 16890
rect 8316 16838 8330 16890
rect 8330 16838 8342 16890
rect 8342 16838 8372 16890
rect 8396 16838 8406 16890
rect 8406 16838 8452 16890
rect 8156 16836 8212 16838
rect 8236 16836 8292 16838
rect 8316 16836 8372 16838
rect 8396 16836 8452 16838
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 10556 17434 10612 17436
rect 10636 17434 10692 17436
rect 10716 17434 10772 17436
rect 10796 17434 10852 17436
rect 10556 17382 10602 17434
rect 10602 17382 10612 17434
rect 10636 17382 10666 17434
rect 10666 17382 10678 17434
rect 10678 17382 10692 17434
rect 10716 17382 10730 17434
rect 10730 17382 10742 17434
rect 10742 17382 10772 17434
rect 10796 17382 10806 17434
rect 10806 17382 10852 17434
rect 10556 17380 10612 17382
rect 10636 17380 10692 17382
rect 10716 17380 10772 17382
rect 10796 17380 10852 17382
rect 15356 17434 15412 17436
rect 15436 17434 15492 17436
rect 15516 17434 15572 17436
rect 15596 17434 15652 17436
rect 15356 17382 15402 17434
rect 15402 17382 15412 17434
rect 15436 17382 15466 17434
rect 15466 17382 15478 17434
rect 15478 17382 15492 17434
rect 15516 17382 15530 17434
rect 15530 17382 15542 17434
rect 15542 17382 15572 17434
rect 15596 17382 15606 17434
rect 15606 17382 15652 17434
rect 15356 17380 15412 17382
rect 15436 17380 15492 17382
rect 15516 17380 15572 17382
rect 15596 17380 15652 17382
rect 8156 15802 8212 15804
rect 8236 15802 8292 15804
rect 8316 15802 8372 15804
rect 8396 15802 8452 15804
rect 8156 15750 8202 15802
rect 8202 15750 8212 15802
rect 8236 15750 8266 15802
rect 8266 15750 8278 15802
rect 8278 15750 8292 15802
rect 8316 15750 8330 15802
rect 8330 15750 8342 15802
rect 8342 15750 8372 15802
rect 8396 15750 8406 15802
rect 8406 15750 8452 15802
rect 8156 15748 8212 15750
rect 8236 15748 8292 15750
rect 8316 15748 8372 15750
rect 8396 15748 8452 15750
rect 10556 16346 10612 16348
rect 10636 16346 10692 16348
rect 10716 16346 10772 16348
rect 10796 16346 10852 16348
rect 10556 16294 10602 16346
rect 10602 16294 10612 16346
rect 10636 16294 10666 16346
rect 10666 16294 10678 16346
rect 10678 16294 10692 16346
rect 10716 16294 10730 16346
rect 10730 16294 10742 16346
rect 10742 16294 10772 16346
rect 10796 16294 10806 16346
rect 10806 16294 10852 16346
rect 10556 16292 10612 16294
rect 10636 16292 10692 16294
rect 10716 16292 10772 16294
rect 10796 16292 10852 16294
rect 3356 11450 3412 11452
rect 3436 11450 3492 11452
rect 3516 11450 3572 11452
rect 3596 11450 3652 11452
rect 3356 11398 3402 11450
rect 3402 11398 3412 11450
rect 3436 11398 3466 11450
rect 3466 11398 3478 11450
rect 3478 11398 3492 11450
rect 3516 11398 3530 11450
rect 3530 11398 3542 11450
rect 3542 11398 3572 11450
rect 3596 11398 3606 11450
rect 3606 11398 3652 11450
rect 3356 11396 3412 11398
rect 3436 11396 3492 11398
rect 3516 11396 3572 11398
rect 3596 11396 3652 11398
rect 3356 10362 3412 10364
rect 3436 10362 3492 10364
rect 3516 10362 3572 10364
rect 3596 10362 3652 10364
rect 3356 10310 3402 10362
rect 3402 10310 3412 10362
rect 3436 10310 3466 10362
rect 3466 10310 3478 10362
rect 3478 10310 3492 10362
rect 3516 10310 3530 10362
rect 3530 10310 3542 10362
rect 3542 10310 3572 10362
rect 3596 10310 3606 10362
rect 3606 10310 3652 10362
rect 3356 10308 3412 10310
rect 3436 10308 3492 10310
rect 3516 10308 3572 10310
rect 3596 10308 3652 10310
rect 3356 9274 3412 9276
rect 3436 9274 3492 9276
rect 3516 9274 3572 9276
rect 3596 9274 3652 9276
rect 3356 9222 3402 9274
rect 3402 9222 3412 9274
rect 3436 9222 3466 9274
rect 3466 9222 3478 9274
rect 3478 9222 3492 9274
rect 3516 9222 3530 9274
rect 3530 9222 3542 9274
rect 3542 9222 3572 9274
rect 3596 9222 3606 9274
rect 3606 9222 3652 9274
rect 3356 9220 3412 9222
rect 3436 9220 3492 9222
rect 3516 9220 3572 9222
rect 3596 9220 3652 9222
rect 1582 7540 1638 7576
rect 1582 7520 1584 7540
rect 1584 7520 1636 7540
rect 1636 7520 1638 7540
rect 3356 8186 3412 8188
rect 3436 8186 3492 8188
rect 3516 8186 3572 8188
rect 3596 8186 3652 8188
rect 3356 8134 3402 8186
rect 3402 8134 3412 8186
rect 3436 8134 3466 8186
rect 3466 8134 3478 8186
rect 3478 8134 3492 8186
rect 3516 8134 3530 8186
rect 3530 8134 3542 8186
rect 3542 8134 3572 8186
rect 3596 8134 3606 8186
rect 3606 8134 3652 8186
rect 3356 8132 3412 8134
rect 3436 8132 3492 8134
rect 3516 8132 3572 8134
rect 3596 8132 3652 8134
rect 5756 14170 5812 14172
rect 5836 14170 5892 14172
rect 5916 14170 5972 14172
rect 5996 14170 6052 14172
rect 5756 14118 5802 14170
rect 5802 14118 5812 14170
rect 5836 14118 5866 14170
rect 5866 14118 5878 14170
rect 5878 14118 5892 14170
rect 5916 14118 5930 14170
rect 5930 14118 5942 14170
rect 5942 14118 5972 14170
rect 5996 14118 6006 14170
rect 6006 14118 6052 14170
rect 5756 14116 5812 14118
rect 5836 14116 5892 14118
rect 5916 14116 5972 14118
rect 5996 14116 6052 14118
rect 8156 14714 8212 14716
rect 8236 14714 8292 14716
rect 8316 14714 8372 14716
rect 8396 14714 8452 14716
rect 8156 14662 8202 14714
rect 8202 14662 8212 14714
rect 8236 14662 8266 14714
rect 8266 14662 8278 14714
rect 8278 14662 8292 14714
rect 8316 14662 8330 14714
rect 8330 14662 8342 14714
rect 8342 14662 8372 14714
rect 8396 14662 8406 14714
rect 8406 14662 8452 14714
rect 8156 14660 8212 14662
rect 8236 14660 8292 14662
rect 8316 14660 8372 14662
rect 8396 14660 8452 14662
rect 5756 13082 5812 13084
rect 5836 13082 5892 13084
rect 5916 13082 5972 13084
rect 5996 13082 6052 13084
rect 5756 13030 5802 13082
rect 5802 13030 5812 13082
rect 5836 13030 5866 13082
rect 5866 13030 5878 13082
rect 5878 13030 5892 13082
rect 5916 13030 5930 13082
rect 5930 13030 5942 13082
rect 5942 13030 5972 13082
rect 5996 13030 6006 13082
rect 6006 13030 6052 13082
rect 5756 13028 5812 13030
rect 5836 13028 5892 13030
rect 5916 13028 5972 13030
rect 5996 13028 6052 13030
rect 5756 11994 5812 11996
rect 5836 11994 5892 11996
rect 5916 11994 5972 11996
rect 5996 11994 6052 11996
rect 5756 11942 5802 11994
rect 5802 11942 5812 11994
rect 5836 11942 5866 11994
rect 5866 11942 5878 11994
rect 5878 11942 5892 11994
rect 5916 11942 5930 11994
rect 5930 11942 5942 11994
rect 5942 11942 5972 11994
rect 5996 11942 6006 11994
rect 6006 11942 6052 11994
rect 5756 11940 5812 11942
rect 5836 11940 5892 11942
rect 5916 11940 5972 11942
rect 5996 11940 6052 11942
rect 5756 10906 5812 10908
rect 5836 10906 5892 10908
rect 5916 10906 5972 10908
rect 5996 10906 6052 10908
rect 5756 10854 5802 10906
rect 5802 10854 5812 10906
rect 5836 10854 5866 10906
rect 5866 10854 5878 10906
rect 5878 10854 5892 10906
rect 5916 10854 5930 10906
rect 5930 10854 5942 10906
rect 5942 10854 5972 10906
rect 5996 10854 6006 10906
rect 6006 10854 6052 10906
rect 5756 10852 5812 10854
rect 5836 10852 5892 10854
rect 5916 10852 5972 10854
rect 5996 10852 6052 10854
rect 5756 9818 5812 9820
rect 5836 9818 5892 9820
rect 5916 9818 5972 9820
rect 5996 9818 6052 9820
rect 5756 9766 5802 9818
rect 5802 9766 5812 9818
rect 5836 9766 5866 9818
rect 5866 9766 5878 9818
rect 5878 9766 5892 9818
rect 5916 9766 5930 9818
rect 5930 9766 5942 9818
rect 5942 9766 5972 9818
rect 5996 9766 6006 9818
rect 6006 9766 6052 9818
rect 5756 9764 5812 9766
rect 5836 9764 5892 9766
rect 5916 9764 5972 9766
rect 5996 9764 6052 9766
rect 8156 13626 8212 13628
rect 8236 13626 8292 13628
rect 8316 13626 8372 13628
rect 8396 13626 8452 13628
rect 8156 13574 8202 13626
rect 8202 13574 8212 13626
rect 8236 13574 8266 13626
rect 8266 13574 8278 13626
rect 8278 13574 8292 13626
rect 8316 13574 8330 13626
rect 8330 13574 8342 13626
rect 8342 13574 8372 13626
rect 8396 13574 8406 13626
rect 8406 13574 8452 13626
rect 8156 13572 8212 13574
rect 8236 13572 8292 13574
rect 8316 13572 8372 13574
rect 8396 13572 8452 13574
rect 10556 15258 10612 15260
rect 10636 15258 10692 15260
rect 10716 15258 10772 15260
rect 10796 15258 10852 15260
rect 10556 15206 10602 15258
rect 10602 15206 10612 15258
rect 10636 15206 10666 15258
rect 10666 15206 10678 15258
rect 10678 15206 10692 15258
rect 10716 15206 10730 15258
rect 10730 15206 10742 15258
rect 10742 15206 10772 15258
rect 10796 15206 10806 15258
rect 10806 15206 10852 15258
rect 10556 15204 10612 15206
rect 10636 15204 10692 15206
rect 10716 15204 10772 15206
rect 10796 15204 10852 15206
rect 10556 14170 10612 14172
rect 10636 14170 10692 14172
rect 10716 14170 10772 14172
rect 10796 14170 10852 14172
rect 10556 14118 10602 14170
rect 10602 14118 10612 14170
rect 10636 14118 10666 14170
rect 10666 14118 10678 14170
rect 10678 14118 10692 14170
rect 10716 14118 10730 14170
rect 10730 14118 10742 14170
rect 10742 14118 10772 14170
rect 10796 14118 10806 14170
rect 10806 14118 10852 14170
rect 10556 14116 10612 14118
rect 10636 14116 10692 14118
rect 10716 14116 10772 14118
rect 10796 14116 10852 14118
rect 8156 12538 8212 12540
rect 8236 12538 8292 12540
rect 8316 12538 8372 12540
rect 8396 12538 8452 12540
rect 8156 12486 8202 12538
rect 8202 12486 8212 12538
rect 8236 12486 8266 12538
rect 8266 12486 8278 12538
rect 8278 12486 8292 12538
rect 8316 12486 8330 12538
rect 8330 12486 8342 12538
rect 8342 12486 8372 12538
rect 8396 12486 8406 12538
rect 8406 12486 8452 12538
rect 8156 12484 8212 12486
rect 8236 12484 8292 12486
rect 8316 12484 8372 12486
rect 8396 12484 8452 12486
rect 8156 11450 8212 11452
rect 8236 11450 8292 11452
rect 8316 11450 8372 11452
rect 8396 11450 8452 11452
rect 8156 11398 8202 11450
rect 8202 11398 8212 11450
rect 8236 11398 8266 11450
rect 8266 11398 8278 11450
rect 8278 11398 8292 11450
rect 8316 11398 8330 11450
rect 8330 11398 8342 11450
rect 8342 11398 8372 11450
rect 8396 11398 8406 11450
rect 8406 11398 8452 11450
rect 8156 11396 8212 11398
rect 8236 11396 8292 11398
rect 8316 11396 8372 11398
rect 8396 11396 8452 11398
rect 8156 10362 8212 10364
rect 8236 10362 8292 10364
rect 8316 10362 8372 10364
rect 8396 10362 8452 10364
rect 8156 10310 8202 10362
rect 8202 10310 8212 10362
rect 8236 10310 8266 10362
rect 8266 10310 8278 10362
rect 8278 10310 8292 10362
rect 8316 10310 8330 10362
rect 8330 10310 8342 10362
rect 8342 10310 8372 10362
rect 8396 10310 8406 10362
rect 8406 10310 8452 10362
rect 8156 10308 8212 10310
rect 8236 10308 8292 10310
rect 8316 10308 8372 10310
rect 8396 10308 8452 10310
rect 8156 9274 8212 9276
rect 8236 9274 8292 9276
rect 8316 9274 8372 9276
rect 8396 9274 8452 9276
rect 8156 9222 8202 9274
rect 8202 9222 8212 9274
rect 8236 9222 8266 9274
rect 8266 9222 8278 9274
rect 8278 9222 8292 9274
rect 8316 9222 8330 9274
rect 8330 9222 8342 9274
rect 8342 9222 8372 9274
rect 8396 9222 8406 9274
rect 8406 9222 8452 9274
rect 8156 9220 8212 9222
rect 8236 9220 8292 9222
rect 8316 9220 8372 9222
rect 8396 9220 8452 9222
rect 5756 8730 5812 8732
rect 5836 8730 5892 8732
rect 5916 8730 5972 8732
rect 5996 8730 6052 8732
rect 5756 8678 5802 8730
rect 5802 8678 5812 8730
rect 5836 8678 5866 8730
rect 5866 8678 5878 8730
rect 5878 8678 5892 8730
rect 5916 8678 5930 8730
rect 5930 8678 5942 8730
rect 5942 8678 5972 8730
rect 5996 8678 6006 8730
rect 6006 8678 6052 8730
rect 5756 8676 5812 8678
rect 5836 8676 5892 8678
rect 5916 8676 5972 8678
rect 5996 8676 6052 8678
rect 10556 13082 10612 13084
rect 10636 13082 10692 13084
rect 10716 13082 10772 13084
rect 10796 13082 10852 13084
rect 10556 13030 10602 13082
rect 10602 13030 10612 13082
rect 10636 13030 10666 13082
rect 10666 13030 10678 13082
rect 10678 13030 10692 13082
rect 10716 13030 10730 13082
rect 10730 13030 10742 13082
rect 10742 13030 10772 13082
rect 10796 13030 10806 13082
rect 10806 13030 10852 13082
rect 10556 13028 10612 13030
rect 10636 13028 10692 13030
rect 10716 13028 10772 13030
rect 10796 13028 10852 13030
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 15356 16346 15412 16348
rect 15436 16346 15492 16348
rect 15516 16346 15572 16348
rect 15596 16346 15652 16348
rect 15356 16294 15402 16346
rect 15402 16294 15412 16346
rect 15436 16294 15466 16346
rect 15466 16294 15478 16346
rect 15478 16294 15492 16346
rect 15516 16294 15530 16346
rect 15530 16294 15542 16346
rect 15542 16294 15572 16346
rect 15596 16294 15606 16346
rect 15606 16294 15652 16346
rect 15356 16292 15412 16294
rect 15436 16292 15492 16294
rect 15516 16292 15572 16294
rect 15596 16292 15652 16294
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 15356 15258 15412 15260
rect 15436 15258 15492 15260
rect 15516 15258 15572 15260
rect 15596 15258 15652 15260
rect 15356 15206 15402 15258
rect 15402 15206 15412 15258
rect 15436 15206 15466 15258
rect 15466 15206 15478 15258
rect 15478 15206 15492 15258
rect 15516 15206 15530 15258
rect 15530 15206 15542 15258
rect 15542 15206 15572 15258
rect 15596 15206 15606 15258
rect 15606 15206 15652 15258
rect 15356 15204 15412 15206
rect 15436 15204 15492 15206
rect 15516 15204 15572 15206
rect 15596 15204 15652 15206
rect 15356 14170 15412 14172
rect 15436 14170 15492 14172
rect 15516 14170 15572 14172
rect 15596 14170 15652 14172
rect 15356 14118 15402 14170
rect 15402 14118 15412 14170
rect 15436 14118 15466 14170
rect 15466 14118 15478 14170
rect 15478 14118 15492 14170
rect 15516 14118 15530 14170
rect 15530 14118 15542 14170
rect 15542 14118 15572 14170
rect 15596 14118 15606 14170
rect 15606 14118 15652 14170
rect 15356 14116 15412 14118
rect 15436 14116 15492 14118
rect 15516 14116 15572 14118
rect 15596 14116 15652 14118
rect 3356 7098 3412 7100
rect 3436 7098 3492 7100
rect 3516 7098 3572 7100
rect 3596 7098 3652 7100
rect 3356 7046 3402 7098
rect 3402 7046 3412 7098
rect 3436 7046 3466 7098
rect 3466 7046 3478 7098
rect 3478 7046 3492 7098
rect 3516 7046 3530 7098
rect 3530 7046 3542 7098
rect 3542 7046 3572 7098
rect 3596 7046 3606 7098
rect 3606 7046 3652 7098
rect 3356 7044 3412 7046
rect 3436 7044 3492 7046
rect 3516 7044 3572 7046
rect 3596 7044 3652 7046
rect 3356 6010 3412 6012
rect 3436 6010 3492 6012
rect 3516 6010 3572 6012
rect 3596 6010 3652 6012
rect 3356 5958 3402 6010
rect 3402 5958 3412 6010
rect 3436 5958 3466 6010
rect 3466 5958 3478 6010
rect 3478 5958 3492 6010
rect 3516 5958 3530 6010
rect 3530 5958 3542 6010
rect 3542 5958 3572 6010
rect 3596 5958 3606 6010
rect 3606 5958 3652 6010
rect 3356 5956 3412 5958
rect 3436 5956 3492 5958
rect 3516 5956 3572 5958
rect 3596 5956 3652 5958
rect 3356 4922 3412 4924
rect 3436 4922 3492 4924
rect 3516 4922 3572 4924
rect 3596 4922 3652 4924
rect 3356 4870 3402 4922
rect 3402 4870 3412 4922
rect 3436 4870 3466 4922
rect 3466 4870 3478 4922
rect 3478 4870 3492 4922
rect 3516 4870 3530 4922
rect 3530 4870 3542 4922
rect 3542 4870 3572 4922
rect 3596 4870 3606 4922
rect 3606 4870 3652 4922
rect 3356 4868 3412 4870
rect 3436 4868 3492 4870
rect 3516 4868 3572 4870
rect 3596 4868 3652 4870
rect 3356 3834 3412 3836
rect 3436 3834 3492 3836
rect 3516 3834 3572 3836
rect 3596 3834 3652 3836
rect 3356 3782 3402 3834
rect 3402 3782 3412 3834
rect 3436 3782 3466 3834
rect 3466 3782 3478 3834
rect 3478 3782 3492 3834
rect 3516 3782 3530 3834
rect 3530 3782 3542 3834
rect 3542 3782 3572 3834
rect 3596 3782 3606 3834
rect 3606 3782 3652 3834
rect 3356 3780 3412 3782
rect 3436 3780 3492 3782
rect 3516 3780 3572 3782
rect 3596 3780 3652 3782
rect 3356 2746 3412 2748
rect 3436 2746 3492 2748
rect 3516 2746 3572 2748
rect 3596 2746 3652 2748
rect 3356 2694 3402 2746
rect 3402 2694 3412 2746
rect 3436 2694 3466 2746
rect 3466 2694 3478 2746
rect 3478 2694 3492 2746
rect 3516 2694 3530 2746
rect 3530 2694 3542 2746
rect 3542 2694 3572 2746
rect 3596 2694 3606 2746
rect 3606 2694 3652 2746
rect 3356 2692 3412 2694
rect 3436 2692 3492 2694
rect 3516 2692 3572 2694
rect 3596 2692 3652 2694
rect 1582 2624 1638 2680
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 8316 8186 8372 8188
rect 8396 8186 8452 8188
rect 8156 8134 8202 8186
rect 8202 8134 8212 8186
rect 8236 8134 8266 8186
rect 8266 8134 8278 8186
rect 8278 8134 8292 8186
rect 8316 8134 8330 8186
rect 8330 8134 8342 8186
rect 8342 8134 8372 8186
rect 8396 8134 8406 8186
rect 8406 8134 8452 8186
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 8316 8132 8372 8134
rect 8396 8132 8452 8134
rect 5756 7642 5812 7644
rect 5836 7642 5892 7644
rect 5916 7642 5972 7644
rect 5996 7642 6052 7644
rect 5756 7590 5802 7642
rect 5802 7590 5812 7642
rect 5836 7590 5866 7642
rect 5866 7590 5878 7642
rect 5878 7590 5892 7642
rect 5916 7590 5930 7642
rect 5930 7590 5942 7642
rect 5942 7590 5972 7642
rect 5996 7590 6006 7642
rect 6006 7590 6052 7642
rect 5756 7588 5812 7590
rect 5836 7588 5892 7590
rect 5916 7588 5972 7590
rect 5996 7588 6052 7590
rect 5756 6554 5812 6556
rect 5836 6554 5892 6556
rect 5916 6554 5972 6556
rect 5996 6554 6052 6556
rect 5756 6502 5802 6554
rect 5802 6502 5812 6554
rect 5836 6502 5866 6554
rect 5866 6502 5878 6554
rect 5878 6502 5892 6554
rect 5916 6502 5930 6554
rect 5930 6502 5942 6554
rect 5942 6502 5972 6554
rect 5996 6502 6006 6554
rect 6006 6502 6052 6554
rect 5756 6500 5812 6502
rect 5836 6500 5892 6502
rect 5916 6500 5972 6502
rect 5996 6500 6052 6502
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 8316 7098 8372 7100
rect 8396 7098 8452 7100
rect 8156 7046 8202 7098
rect 8202 7046 8212 7098
rect 8236 7046 8266 7098
rect 8266 7046 8278 7098
rect 8278 7046 8292 7098
rect 8316 7046 8330 7098
rect 8330 7046 8342 7098
rect 8342 7046 8372 7098
rect 8396 7046 8406 7098
rect 8406 7046 8452 7098
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 8316 7044 8372 7046
rect 8396 7044 8452 7046
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 8316 6010 8372 6012
rect 8396 6010 8452 6012
rect 8156 5958 8202 6010
rect 8202 5958 8212 6010
rect 8236 5958 8266 6010
rect 8266 5958 8278 6010
rect 8278 5958 8292 6010
rect 8316 5958 8330 6010
rect 8330 5958 8342 6010
rect 8342 5958 8372 6010
rect 8396 5958 8406 6010
rect 8406 5958 8452 6010
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 8316 5956 8372 5958
rect 8396 5956 8452 5958
rect 5756 5466 5812 5468
rect 5836 5466 5892 5468
rect 5916 5466 5972 5468
rect 5996 5466 6052 5468
rect 5756 5414 5802 5466
rect 5802 5414 5812 5466
rect 5836 5414 5866 5466
rect 5866 5414 5878 5466
rect 5878 5414 5892 5466
rect 5916 5414 5930 5466
rect 5930 5414 5942 5466
rect 5942 5414 5972 5466
rect 5996 5414 6006 5466
rect 6006 5414 6052 5466
rect 5756 5412 5812 5414
rect 5836 5412 5892 5414
rect 5916 5412 5972 5414
rect 5996 5412 6052 5414
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 8316 4922 8372 4924
rect 8396 4922 8452 4924
rect 8156 4870 8202 4922
rect 8202 4870 8212 4922
rect 8236 4870 8266 4922
rect 8266 4870 8278 4922
rect 8278 4870 8292 4922
rect 8316 4870 8330 4922
rect 8330 4870 8342 4922
rect 8342 4870 8372 4922
rect 8396 4870 8406 4922
rect 8406 4870 8452 4922
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 8316 4868 8372 4870
rect 8396 4868 8452 4870
rect 5756 4378 5812 4380
rect 5836 4378 5892 4380
rect 5916 4378 5972 4380
rect 5996 4378 6052 4380
rect 5756 4326 5802 4378
rect 5802 4326 5812 4378
rect 5836 4326 5866 4378
rect 5866 4326 5878 4378
rect 5878 4326 5892 4378
rect 5916 4326 5930 4378
rect 5930 4326 5942 4378
rect 5942 4326 5972 4378
rect 5996 4326 6006 4378
rect 6006 4326 6052 4378
rect 5756 4324 5812 4326
rect 5836 4324 5892 4326
rect 5916 4324 5972 4326
rect 5996 4324 6052 4326
rect 10556 11994 10612 11996
rect 10636 11994 10692 11996
rect 10716 11994 10772 11996
rect 10796 11994 10852 11996
rect 10556 11942 10602 11994
rect 10602 11942 10612 11994
rect 10636 11942 10666 11994
rect 10666 11942 10678 11994
rect 10678 11942 10692 11994
rect 10716 11942 10730 11994
rect 10730 11942 10742 11994
rect 10742 11942 10772 11994
rect 10796 11942 10806 11994
rect 10806 11942 10852 11994
rect 10556 11940 10612 11942
rect 10636 11940 10692 11942
rect 10716 11940 10772 11942
rect 10796 11940 10852 11942
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 10556 10906 10612 10908
rect 10636 10906 10692 10908
rect 10716 10906 10772 10908
rect 10796 10906 10852 10908
rect 10556 10854 10602 10906
rect 10602 10854 10612 10906
rect 10636 10854 10666 10906
rect 10666 10854 10678 10906
rect 10678 10854 10692 10906
rect 10716 10854 10730 10906
rect 10730 10854 10742 10906
rect 10742 10854 10772 10906
rect 10796 10854 10806 10906
rect 10806 10854 10852 10906
rect 10556 10852 10612 10854
rect 10636 10852 10692 10854
rect 10716 10852 10772 10854
rect 10796 10852 10852 10854
rect 10556 9818 10612 9820
rect 10636 9818 10692 9820
rect 10716 9818 10772 9820
rect 10796 9818 10852 9820
rect 10556 9766 10602 9818
rect 10602 9766 10612 9818
rect 10636 9766 10666 9818
rect 10666 9766 10678 9818
rect 10678 9766 10692 9818
rect 10716 9766 10730 9818
rect 10730 9766 10742 9818
rect 10742 9766 10772 9818
rect 10796 9766 10806 9818
rect 10806 9766 10852 9818
rect 10556 9764 10612 9766
rect 10636 9764 10692 9766
rect 10716 9764 10772 9766
rect 10796 9764 10852 9766
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 10556 8730 10612 8732
rect 10636 8730 10692 8732
rect 10716 8730 10772 8732
rect 10796 8730 10852 8732
rect 10556 8678 10602 8730
rect 10602 8678 10612 8730
rect 10636 8678 10666 8730
rect 10666 8678 10678 8730
rect 10678 8678 10692 8730
rect 10716 8678 10730 8730
rect 10730 8678 10742 8730
rect 10742 8678 10772 8730
rect 10796 8678 10806 8730
rect 10806 8678 10852 8730
rect 10556 8676 10612 8678
rect 10636 8676 10692 8678
rect 10716 8676 10772 8678
rect 10796 8676 10852 8678
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 10556 7642 10612 7644
rect 10636 7642 10692 7644
rect 10716 7642 10772 7644
rect 10796 7642 10852 7644
rect 10556 7590 10602 7642
rect 10602 7590 10612 7642
rect 10636 7590 10666 7642
rect 10666 7590 10678 7642
rect 10678 7590 10692 7642
rect 10716 7590 10730 7642
rect 10730 7590 10742 7642
rect 10742 7590 10772 7642
rect 10796 7590 10806 7642
rect 10806 7590 10852 7642
rect 10556 7588 10612 7590
rect 10636 7588 10692 7590
rect 10716 7588 10772 7590
rect 10796 7588 10852 7590
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 10556 6554 10612 6556
rect 10636 6554 10692 6556
rect 10716 6554 10772 6556
rect 10796 6554 10852 6556
rect 10556 6502 10602 6554
rect 10602 6502 10612 6554
rect 10636 6502 10666 6554
rect 10666 6502 10678 6554
rect 10678 6502 10692 6554
rect 10716 6502 10730 6554
rect 10730 6502 10742 6554
rect 10742 6502 10772 6554
rect 10796 6502 10806 6554
rect 10806 6502 10852 6554
rect 10556 6500 10612 6502
rect 10636 6500 10692 6502
rect 10716 6500 10772 6502
rect 10796 6500 10852 6502
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 10556 5466 10612 5468
rect 10636 5466 10692 5468
rect 10716 5466 10772 5468
rect 10796 5466 10852 5468
rect 10556 5414 10602 5466
rect 10602 5414 10612 5466
rect 10636 5414 10666 5466
rect 10666 5414 10678 5466
rect 10678 5414 10692 5466
rect 10716 5414 10730 5466
rect 10730 5414 10742 5466
rect 10742 5414 10772 5466
rect 10796 5414 10806 5466
rect 10806 5414 10852 5466
rect 10556 5412 10612 5414
rect 10636 5412 10692 5414
rect 10716 5412 10772 5414
rect 10796 5412 10852 5414
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 10556 4378 10612 4380
rect 10636 4378 10692 4380
rect 10716 4378 10772 4380
rect 10796 4378 10852 4380
rect 10556 4326 10602 4378
rect 10602 4326 10612 4378
rect 10636 4326 10666 4378
rect 10666 4326 10678 4378
rect 10678 4326 10692 4378
rect 10716 4326 10730 4378
rect 10730 4326 10742 4378
rect 10742 4326 10772 4378
rect 10796 4326 10806 4378
rect 10806 4326 10852 4378
rect 10556 4324 10612 4326
rect 10636 4324 10692 4326
rect 10716 4324 10772 4326
rect 10796 4324 10852 4326
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 8316 3834 8372 3836
rect 8396 3834 8452 3836
rect 8156 3782 8202 3834
rect 8202 3782 8212 3834
rect 8236 3782 8266 3834
rect 8266 3782 8278 3834
rect 8278 3782 8292 3834
rect 8316 3782 8330 3834
rect 8330 3782 8342 3834
rect 8342 3782 8372 3834
rect 8396 3782 8406 3834
rect 8406 3782 8452 3834
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 8316 3780 8372 3782
rect 8396 3780 8452 3782
rect 5756 3290 5812 3292
rect 5836 3290 5892 3292
rect 5916 3290 5972 3292
rect 5996 3290 6052 3292
rect 5756 3238 5802 3290
rect 5802 3238 5812 3290
rect 5836 3238 5866 3290
rect 5866 3238 5878 3290
rect 5878 3238 5892 3290
rect 5916 3238 5930 3290
rect 5930 3238 5942 3290
rect 5942 3238 5972 3290
rect 5996 3238 6006 3290
rect 6006 3238 6052 3290
rect 5756 3236 5812 3238
rect 5836 3236 5892 3238
rect 5916 3236 5972 3238
rect 5996 3236 6052 3238
rect 10556 3290 10612 3292
rect 10636 3290 10692 3292
rect 10716 3290 10772 3292
rect 10796 3290 10852 3292
rect 10556 3238 10602 3290
rect 10602 3238 10612 3290
rect 10636 3238 10666 3290
rect 10666 3238 10678 3290
rect 10678 3238 10692 3290
rect 10716 3238 10730 3290
rect 10730 3238 10742 3290
rect 10742 3238 10772 3290
rect 10796 3238 10806 3290
rect 10806 3238 10852 3290
rect 10556 3236 10612 3238
rect 10636 3236 10692 3238
rect 10716 3236 10772 3238
rect 10796 3236 10852 3238
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 8316 2746 8372 2748
rect 8396 2746 8452 2748
rect 8156 2694 8202 2746
rect 8202 2694 8212 2746
rect 8236 2694 8266 2746
rect 8266 2694 8278 2746
rect 8278 2694 8292 2746
rect 8316 2694 8330 2746
rect 8330 2694 8342 2746
rect 8342 2694 8372 2746
rect 8396 2694 8406 2746
rect 8406 2694 8452 2746
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 8316 2692 8372 2694
rect 8396 2692 8452 2694
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 15356 13082 15412 13084
rect 15436 13082 15492 13084
rect 15516 13082 15572 13084
rect 15596 13082 15652 13084
rect 15356 13030 15402 13082
rect 15402 13030 15412 13082
rect 15436 13030 15466 13082
rect 15466 13030 15478 13082
rect 15478 13030 15492 13082
rect 15516 13030 15530 13082
rect 15530 13030 15542 13082
rect 15542 13030 15572 13082
rect 15596 13030 15606 13082
rect 15606 13030 15652 13082
rect 15356 13028 15412 13030
rect 15436 13028 15492 13030
rect 15516 13028 15572 13030
rect 15596 13028 15652 13030
rect 15356 11994 15412 11996
rect 15436 11994 15492 11996
rect 15516 11994 15572 11996
rect 15596 11994 15652 11996
rect 15356 11942 15402 11994
rect 15402 11942 15412 11994
rect 15436 11942 15466 11994
rect 15466 11942 15478 11994
rect 15478 11942 15492 11994
rect 15516 11942 15530 11994
rect 15530 11942 15542 11994
rect 15542 11942 15572 11994
rect 15596 11942 15606 11994
rect 15606 11942 15652 11994
rect 15356 11940 15412 11942
rect 15436 11940 15492 11942
rect 15516 11940 15572 11942
rect 15596 11940 15652 11942
rect 15356 10906 15412 10908
rect 15436 10906 15492 10908
rect 15516 10906 15572 10908
rect 15596 10906 15652 10908
rect 15356 10854 15402 10906
rect 15402 10854 15412 10906
rect 15436 10854 15466 10906
rect 15466 10854 15478 10906
rect 15478 10854 15492 10906
rect 15516 10854 15530 10906
rect 15530 10854 15542 10906
rect 15542 10854 15572 10906
rect 15596 10854 15606 10906
rect 15606 10854 15652 10906
rect 15356 10852 15412 10854
rect 15436 10852 15492 10854
rect 15516 10852 15572 10854
rect 15596 10852 15652 10854
rect 20156 21786 20212 21788
rect 20236 21786 20292 21788
rect 20316 21786 20372 21788
rect 20396 21786 20452 21788
rect 20156 21734 20202 21786
rect 20202 21734 20212 21786
rect 20236 21734 20266 21786
rect 20266 21734 20278 21786
rect 20278 21734 20292 21786
rect 20316 21734 20330 21786
rect 20330 21734 20342 21786
rect 20342 21734 20372 21786
rect 20396 21734 20406 21786
rect 20406 21734 20452 21786
rect 20156 21732 20212 21734
rect 20236 21732 20292 21734
rect 20316 21732 20372 21734
rect 20396 21732 20452 21734
rect 20156 20698 20212 20700
rect 20236 20698 20292 20700
rect 20316 20698 20372 20700
rect 20396 20698 20452 20700
rect 20156 20646 20202 20698
rect 20202 20646 20212 20698
rect 20236 20646 20266 20698
rect 20266 20646 20278 20698
rect 20278 20646 20292 20698
rect 20316 20646 20330 20698
rect 20330 20646 20342 20698
rect 20342 20646 20372 20698
rect 20396 20646 20406 20698
rect 20406 20646 20452 20698
rect 20156 20644 20212 20646
rect 20236 20644 20292 20646
rect 20316 20644 20372 20646
rect 20396 20644 20452 20646
rect 17756 19066 17812 19068
rect 17836 19066 17892 19068
rect 17916 19066 17972 19068
rect 17996 19066 18052 19068
rect 17756 19014 17802 19066
rect 17802 19014 17812 19066
rect 17836 19014 17866 19066
rect 17866 19014 17878 19066
rect 17878 19014 17892 19066
rect 17916 19014 17930 19066
rect 17930 19014 17942 19066
rect 17942 19014 17972 19066
rect 17996 19014 18006 19066
rect 18006 19014 18052 19066
rect 17756 19012 17812 19014
rect 17836 19012 17892 19014
rect 17916 19012 17972 19014
rect 17996 19012 18052 19014
rect 17756 17978 17812 17980
rect 17836 17978 17892 17980
rect 17916 17978 17972 17980
rect 17996 17978 18052 17980
rect 17756 17926 17802 17978
rect 17802 17926 17812 17978
rect 17836 17926 17866 17978
rect 17866 17926 17878 17978
rect 17878 17926 17892 17978
rect 17916 17926 17930 17978
rect 17930 17926 17942 17978
rect 17942 17926 17972 17978
rect 17996 17926 18006 17978
rect 18006 17926 18052 17978
rect 17756 17924 17812 17926
rect 17836 17924 17892 17926
rect 17916 17924 17972 17926
rect 17996 17924 18052 17926
rect 17756 16890 17812 16892
rect 17836 16890 17892 16892
rect 17916 16890 17972 16892
rect 17996 16890 18052 16892
rect 17756 16838 17802 16890
rect 17802 16838 17812 16890
rect 17836 16838 17866 16890
rect 17866 16838 17878 16890
rect 17878 16838 17892 16890
rect 17916 16838 17930 16890
rect 17930 16838 17942 16890
rect 17942 16838 17972 16890
rect 17996 16838 18006 16890
rect 18006 16838 18052 16890
rect 17756 16836 17812 16838
rect 17836 16836 17892 16838
rect 17916 16836 17972 16838
rect 17996 16836 18052 16838
rect 22556 21242 22612 21244
rect 22636 21242 22692 21244
rect 22716 21242 22772 21244
rect 22796 21242 22852 21244
rect 22556 21190 22602 21242
rect 22602 21190 22612 21242
rect 22636 21190 22666 21242
rect 22666 21190 22678 21242
rect 22678 21190 22692 21242
rect 22716 21190 22730 21242
rect 22730 21190 22742 21242
rect 22742 21190 22772 21242
rect 22796 21190 22806 21242
rect 22806 21190 22852 21242
rect 22556 21188 22612 21190
rect 22636 21188 22692 21190
rect 22716 21188 22772 21190
rect 22796 21188 22852 21190
rect 24956 21786 25012 21788
rect 25036 21786 25092 21788
rect 25116 21786 25172 21788
rect 25196 21786 25252 21788
rect 24956 21734 25002 21786
rect 25002 21734 25012 21786
rect 25036 21734 25066 21786
rect 25066 21734 25078 21786
rect 25078 21734 25092 21786
rect 25116 21734 25130 21786
rect 25130 21734 25142 21786
rect 25142 21734 25172 21786
rect 25196 21734 25206 21786
rect 25206 21734 25252 21786
rect 24956 21732 25012 21734
rect 25036 21732 25092 21734
rect 25116 21732 25172 21734
rect 25196 21732 25252 21734
rect 24956 20698 25012 20700
rect 25036 20698 25092 20700
rect 25116 20698 25172 20700
rect 25196 20698 25252 20700
rect 24956 20646 25002 20698
rect 25002 20646 25012 20698
rect 25036 20646 25066 20698
rect 25066 20646 25078 20698
rect 25078 20646 25092 20698
rect 25116 20646 25130 20698
rect 25130 20646 25142 20698
rect 25142 20646 25172 20698
rect 25196 20646 25206 20698
rect 25206 20646 25252 20698
rect 24956 20644 25012 20646
rect 25036 20644 25092 20646
rect 25116 20644 25172 20646
rect 25196 20644 25252 20646
rect 20156 19610 20212 19612
rect 20236 19610 20292 19612
rect 20316 19610 20372 19612
rect 20396 19610 20452 19612
rect 20156 19558 20202 19610
rect 20202 19558 20212 19610
rect 20236 19558 20266 19610
rect 20266 19558 20278 19610
rect 20278 19558 20292 19610
rect 20316 19558 20330 19610
rect 20330 19558 20342 19610
rect 20342 19558 20372 19610
rect 20396 19558 20406 19610
rect 20406 19558 20452 19610
rect 20156 19556 20212 19558
rect 20236 19556 20292 19558
rect 20316 19556 20372 19558
rect 20396 19556 20452 19558
rect 22556 20154 22612 20156
rect 22636 20154 22692 20156
rect 22716 20154 22772 20156
rect 22796 20154 22852 20156
rect 22556 20102 22602 20154
rect 22602 20102 22612 20154
rect 22636 20102 22666 20154
rect 22666 20102 22678 20154
rect 22678 20102 22692 20154
rect 22716 20102 22730 20154
rect 22730 20102 22742 20154
rect 22742 20102 22772 20154
rect 22796 20102 22806 20154
rect 22806 20102 22852 20154
rect 22556 20100 22612 20102
rect 22636 20100 22692 20102
rect 22716 20100 22772 20102
rect 22796 20100 22852 20102
rect 22556 19066 22612 19068
rect 22636 19066 22692 19068
rect 22716 19066 22772 19068
rect 22796 19066 22852 19068
rect 22556 19014 22602 19066
rect 22602 19014 22612 19066
rect 22636 19014 22666 19066
rect 22666 19014 22678 19066
rect 22678 19014 22692 19066
rect 22716 19014 22730 19066
rect 22730 19014 22742 19066
rect 22742 19014 22772 19066
rect 22796 19014 22806 19066
rect 22806 19014 22852 19066
rect 22556 19012 22612 19014
rect 22636 19012 22692 19014
rect 22716 19012 22772 19014
rect 22796 19012 22852 19014
rect 20156 18522 20212 18524
rect 20236 18522 20292 18524
rect 20316 18522 20372 18524
rect 20396 18522 20452 18524
rect 20156 18470 20202 18522
rect 20202 18470 20212 18522
rect 20236 18470 20266 18522
rect 20266 18470 20278 18522
rect 20278 18470 20292 18522
rect 20316 18470 20330 18522
rect 20330 18470 20342 18522
rect 20342 18470 20372 18522
rect 20396 18470 20406 18522
rect 20406 18470 20452 18522
rect 20156 18468 20212 18470
rect 20236 18468 20292 18470
rect 20316 18468 20372 18470
rect 20396 18468 20452 18470
rect 17756 15802 17812 15804
rect 17836 15802 17892 15804
rect 17916 15802 17972 15804
rect 17996 15802 18052 15804
rect 17756 15750 17802 15802
rect 17802 15750 17812 15802
rect 17836 15750 17866 15802
rect 17866 15750 17878 15802
rect 17878 15750 17892 15802
rect 17916 15750 17930 15802
rect 17930 15750 17942 15802
rect 17942 15750 17972 15802
rect 17996 15750 18006 15802
rect 18006 15750 18052 15802
rect 17756 15748 17812 15750
rect 17836 15748 17892 15750
rect 17916 15748 17972 15750
rect 17996 15748 18052 15750
rect 15356 9818 15412 9820
rect 15436 9818 15492 9820
rect 15516 9818 15572 9820
rect 15596 9818 15652 9820
rect 15356 9766 15402 9818
rect 15402 9766 15412 9818
rect 15436 9766 15466 9818
rect 15466 9766 15478 9818
rect 15478 9766 15492 9818
rect 15516 9766 15530 9818
rect 15530 9766 15542 9818
rect 15542 9766 15572 9818
rect 15596 9766 15606 9818
rect 15606 9766 15652 9818
rect 15356 9764 15412 9766
rect 15436 9764 15492 9766
rect 15516 9764 15572 9766
rect 15596 9764 15652 9766
rect 15356 8730 15412 8732
rect 15436 8730 15492 8732
rect 15516 8730 15572 8732
rect 15596 8730 15652 8732
rect 15356 8678 15402 8730
rect 15402 8678 15412 8730
rect 15436 8678 15466 8730
rect 15466 8678 15478 8730
rect 15478 8678 15492 8730
rect 15516 8678 15530 8730
rect 15530 8678 15542 8730
rect 15542 8678 15572 8730
rect 15596 8678 15606 8730
rect 15606 8678 15652 8730
rect 15356 8676 15412 8678
rect 15436 8676 15492 8678
rect 15516 8676 15572 8678
rect 15596 8676 15652 8678
rect 17756 14714 17812 14716
rect 17836 14714 17892 14716
rect 17916 14714 17972 14716
rect 17996 14714 18052 14716
rect 17756 14662 17802 14714
rect 17802 14662 17812 14714
rect 17836 14662 17866 14714
rect 17866 14662 17878 14714
rect 17878 14662 17892 14714
rect 17916 14662 17930 14714
rect 17930 14662 17942 14714
rect 17942 14662 17972 14714
rect 17996 14662 18006 14714
rect 18006 14662 18052 14714
rect 17756 14660 17812 14662
rect 17836 14660 17892 14662
rect 17916 14660 17972 14662
rect 17996 14660 18052 14662
rect 17756 13626 17812 13628
rect 17836 13626 17892 13628
rect 17916 13626 17972 13628
rect 17996 13626 18052 13628
rect 17756 13574 17802 13626
rect 17802 13574 17812 13626
rect 17836 13574 17866 13626
rect 17866 13574 17878 13626
rect 17878 13574 17892 13626
rect 17916 13574 17930 13626
rect 17930 13574 17942 13626
rect 17942 13574 17972 13626
rect 17996 13574 18006 13626
rect 18006 13574 18052 13626
rect 17756 13572 17812 13574
rect 17836 13572 17892 13574
rect 17916 13572 17972 13574
rect 17996 13572 18052 13574
rect 17756 12538 17812 12540
rect 17836 12538 17892 12540
rect 17916 12538 17972 12540
rect 17996 12538 18052 12540
rect 17756 12486 17802 12538
rect 17802 12486 17812 12538
rect 17836 12486 17866 12538
rect 17866 12486 17878 12538
rect 17878 12486 17892 12538
rect 17916 12486 17930 12538
rect 17930 12486 17942 12538
rect 17942 12486 17972 12538
rect 17996 12486 18006 12538
rect 18006 12486 18052 12538
rect 17756 12484 17812 12486
rect 17836 12484 17892 12486
rect 17916 12484 17972 12486
rect 17996 12484 18052 12486
rect 20156 17434 20212 17436
rect 20236 17434 20292 17436
rect 20316 17434 20372 17436
rect 20396 17434 20452 17436
rect 20156 17382 20202 17434
rect 20202 17382 20212 17434
rect 20236 17382 20266 17434
rect 20266 17382 20278 17434
rect 20278 17382 20292 17434
rect 20316 17382 20330 17434
rect 20330 17382 20342 17434
rect 20342 17382 20372 17434
rect 20396 17382 20406 17434
rect 20406 17382 20452 17434
rect 20156 17380 20212 17382
rect 20236 17380 20292 17382
rect 20316 17380 20372 17382
rect 20396 17380 20452 17382
rect 20156 16346 20212 16348
rect 20236 16346 20292 16348
rect 20316 16346 20372 16348
rect 20396 16346 20452 16348
rect 20156 16294 20202 16346
rect 20202 16294 20212 16346
rect 20236 16294 20266 16346
rect 20266 16294 20278 16346
rect 20278 16294 20292 16346
rect 20316 16294 20330 16346
rect 20330 16294 20342 16346
rect 20342 16294 20372 16346
rect 20396 16294 20406 16346
rect 20406 16294 20452 16346
rect 20156 16292 20212 16294
rect 20236 16292 20292 16294
rect 20316 16292 20372 16294
rect 20396 16292 20452 16294
rect 20156 15258 20212 15260
rect 20236 15258 20292 15260
rect 20316 15258 20372 15260
rect 20396 15258 20452 15260
rect 20156 15206 20202 15258
rect 20202 15206 20212 15258
rect 20236 15206 20266 15258
rect 20266 15206 20278 15258
rect 20278 15206 20292 15258
rect 20316 15206 20330 15258
rect 20330 15206 20342 15258
rect 20342 15206 20372 15258
rect 20396 15206 20406 15258
rect 20406 15206 20452 15258
rect 20156 15204 20212 15206
rect 20236 15204 20292 15206
rect 20316 15204 20372 15206
rect 20396 15204 20452 15206
rect 17756 11450 17812 11452
rect 17836 11450 17892 11452
rect 17916 11450 17972 11452
rect 17996 11450 18052 11452
rect 17756 11398 17802 11450
rect 17802 11398 17812 11450
rect 17836 11398 17866 11450
rect 17866 11398 17878 11450
rect 17878 11398 17892 11450
rect 17916 11398 17930 11450
rect 17930 11398 17942 11450
rect 17942 11398 17972 11450
rect 17996 11398 18006 11450
rect 18006 11398 18052 11450
rect 17756 11396 17812 11398
rect 17836 11396 17892 11398
rect 17916 11396 17972 11398
rect 17996 11396 18052 11398
rect 17756 10362 17812 10364
rect 17836 10362 17892 10364
rect 17916 10362 17972 10364
rect 17996 10362 18052 10364
rect 17756 10310 17802 10362
rect 17802 10310 17812 10362
rect 17836 10310 17866 10362
rect 17866 10310 17878 10362
rect 17878 10310 17892 10362
rect 17916 10310 17930 10362
rect 17930 10310 17942 10362
rect 17942 10310 17972 10362
rect 17996 10310 18006 10362
rect 18006 10310 18052 10362
rect 17756 10308 17812 10310
rect 17836 10308 17892 10310
rect 17916 10308 17972 10310
rect 17996 10308 18052 10310
rect 17756 9274 17812 9276
rect 17836 9274 17892 9276
rect 17916 9274 17972 9276
rect 17996 9274 18052 9276
rect 17756 9222 17802 9274
rect 17802 9222 17812 9274
rect 17836 9222 17866 9274
rect 17866 9222 17878 9274
rect 17878 9222 17892 9274
rect 17916 9222 17930 9274
rect 17930 9222 17942 9274
rect 17942 9222 17972 9274
rect 17996 9222 18006 9274
rect 18006 9222 18052 9274
rect 17756 9220 17812 9222
rect 17836 9220 17892 9222
rect 17916 9220 17972 9222
rect 17996 9220 18052 9222
rect 17756 8186 17812 8188
rect 17836 8186 17892 8188
rect 17916 8186 17972 8188
rect 17996 8186 18052 8188
rect 17756 8134 17802 8186
rect 17802 8134 17812 8186
rect 17836 8134 17866 8186
rect 17866 8134 17878 8186
rect 17878 8134 17892 8186
rect 17916 8134 17930 8186
rect 17930 8134 17942 8186
rect 17942 8134 17972 8186
rect 17996 8134 18006 8186
rect 18006 8134 18052 8186
rect 17756 8132 17812 8134
rect 17836 8132 17892 8134
rect 17916 8132 17972 8134
rect 17996 8132 18052 8134
rect 15356 7642 15412 7644
rect 15436 7642 15492 7644
rect 15516 7642 15572 7644
rect 15596 7642 15652 7644
rect 15356 7590 15402 7642
rect 15402 7590 15412 7642
rect 15436 7590 15466 7642
rect 15466 7590 15478 7642
rect 15478 7590 15492 7642
rect 15516 7590 15530 7642
rect 15530 7590 15542 7642
rect 15542 7590 15572 7642
rect 15596 7590 15606 7642
rect 15606 7590 15652 7642
rect 15356 7588 15412 7590
rect 15436 7588 15492 7590
rect 15516 7588 15572 7590
rect 15596 7588 15652 7590
rect 17756 7098 17812 7100
rect 17836 7098 17892 7100
rect 17916 7098 17972 7100
rect 17996 7098 18052 7100
rect 17756 7046 17802 7098
rect 17802 7046 17812 7098
rect 17836 7046 17866 7098
rect 17866 7046 17878 7098
rect 17878 7046 17892 7098
rect 17916 7046 17930 7098
rect 17930 7046 17942 7098
rect 17942 7046 17972 7098
rect 17996 7046 18006 7098
rect 18006 7046 18052 7098
rect 17756 7044 17812 7046
rect 17836 7044 17892 7046
rect 17916 7044 17972 7046
rect 17996 7044 18052 7046
rect 15356 6554 15412 6556
rect 15436 6554 15492 6556
rect 15516 6554 15572 6556
rect 15596 6554 15652 6556
rect 15356 6502 15402 6554
rect 15402 6502 15412 6554
rect 15436 6502 15466 6554
rect 15466 6502 15478 6554
rect 15478 6502 15492 6554
rect 15516 6502 15530 6554
rect 15530 6502 15542 6554
rect 15542 6502 15572 6554
rect 15596 6502 15606 6554
rect 15606 6502 15652 6554
rect 15356 6500 15412 6502
rect 15436 6500 15492 6502
rect 15516 6500 15572 6502
rect 15596 6500 15652 6502
rect 17756 6010 17812 6012
rect 17836 6010 17892 6012
rect 17916 6010 17972 6012
rect 17996 6010 18052 6012
rect 17756 5958 17802 6010
rect 17802 5958 17812 6010
rect 17836 5958 17866 6010
rect 17866 5958 17878 6010
rect 17878 5958 17892 6010
rect 17916 5958 17930 6010
rect 17930 5958 17942 6010
rect 17942 5958 17972 6010
rect 17996 5958 18006 6010
rect 18006 5958 18052 6010
rect 17756 5956 17812 5958
rect 17836 5956 17892 5958
rect 17916 5956 17972 5958
rect 17996 5956 18052 5958
rect 15356 5466 15412 5468
rect 15436 5466 15492 5468
rect 15516 5466 15572 5468
rect 15596 5466 15652 5468
rect 15356 5414 15402 5466
rect 15402 5414 15412 5466
rect 15436 5414 15466 5466
rect 15466 5414 15478 5466
rect 15478 5414 15492 5466
rect 15516 5414 15530 5466
rect 15530 5414 15542 5466
rect 15542 5414 15572 5466
rect 15596 5414 15606 5466
rect 15606 5414 15652 5466
rect 15356 5412 15412 5414
rect 15436 5412 15492 5414
rect 15516 5412 15572 5414
rect 15596 5412 15652 5414
rect 17756 4922 17812 4924
rect 17836 4922 17892 4924
rect 17916 4922 17972 4924
rect 17996 4922 18052 4924
rect 17756 4870 17802 4922
rect 17802 4870 17812 4922
rect 17836 4870 17866 4922
rect 17866 4870 17878 4922
rect 17878 4870 17892 4922
rect 17916 4870 17930 4922
rect 17930 4870 17942 4922
rect 17942 4870 17972 4922
rect 17996 4870 18006 4922
rect 18006 4870 18052 4922
rect 17756 4868 17812 4870
rect 17836 4868 17892 4870
rect 17916 4868 17972 4870
rect 17996 4868 18052 4870
rect 15356 4378 15412 4380
rect 15436 4378 15492 4380
rect 15516 4378 15572 4380
rect 15596 4378 15652 4380
rect 15356 4326 15402 4378
rect 15402 4326 15412 4378
rect 15436 4326 15466 4378
rect 15466 4326 15478 4378
rect 15478 4326 15492 4378
rect 15516 4326 15530 4378
rect 15530 4326 15542 4378
rect 15542 4326 15572 4378
rect 15596 4326 15606 4378
rect 15606 4326 15652 4378
rect 15356 4324 15412 4326
rect 15436 4324 15492 4326
rect 15516 4324 15572 4326
rect 15596 4324 15652 4326
rect 17756 3834 17812 3836
rect 17836 3834 17892 3836
rect 17916 3834 17972 3836
rect 17996 3834 18052 3836
rect 17756 3782 17802 3834
rect 17802 3782 17812 3834
rect 17836 3782 17866 3834
rect 17866 3782 17878 3834
rect 17878 3782 17892 3834
rect 17916 3782 17930 3834
rect 17930 3782 17942 3834
rect 17942 3782 17972 3834
rect 17996 3782 18006 3834
rect 18006 3782 18052 3834
rect 17756 3780 17812 3782
rect 17836 3780 17892 3782
rect 17916 3780 17972 3782
rect 17996 3780 18052 3782
rect 15356 3290 15412 3292
rect 15436 3290 15492 3292
rect 15516 3290 15572 3292
rect 15596 3290 15652 3292
rect 15356 3238 15402 3290
rect 15402 3238 15412 3290
rect 15436 3238 15466 3290
rect 15466 3238 15478 3290
rect 15478 3238 15492 3290
rect 15516 3238 15530 3290
rect 15530 3238 15542 3290
rect 15542 3238 15572 3290
rect 15596 3238 15606 3290
rect 15606 3238 15652 3290
rect 15356 3236 15412 3238
rect 15436 3236 15492 3238
rect 15516 3236 15572 3238
rect 15596 3236 15652 3238
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17756 2746 17812 2748
rect 17836 2746 17892 2748
rect 17916 2746 17972 2748
rect 17996 2746 18052 2748
rect 17756 2694 17802 2746
rect 17802 2694 17812 2746
rect 17836 2694 17866 2746
rect 17866 2694 17878 2746
rect 17878 2694 17892 2746
rect 17916 2694 17930 2746
rect 17930 2694 17942 2746
rect 17942 2694 17972 2746
rect 17996 2694 18006 2746
rect 18006 2694 18052 2746
rect 17756 2692 17812 2694
rect 17836 2692 17892 2694
rect 17916 2692 17972 2694
rect 17996 2692 18052 2694
rect 20156 14170 20212 14172
rect 20236 14170 20292 14172
rect 20316 14170 20372 14172
rect 20396 14170 20452 14172
rect 20156 14118 20202 14170
rect 20202 14118 20212 14170
rect 20236 14118 20266 14170
rect 20266 14118 20278 14170
rect 20278 14118 20292 14170
rect 20316 14118 20330 14170
rect 20330 14118 20342 14170
rect 20342 14118 20372 14170
rect 20396 14118 20406 14170
rect 20406 14118 20452 14170
rect 20156 14116 20212 14118
rect 20236 14116 20292 14118
rect 20316 14116 20372 14118
rect 20396 14116 20452 14118
rect 20156 13082 20212 13084
rect 20236 13082 20292 13084
rect 20316 13082 20372 13084
rect 20396 13082 20452 13084
rect 20156 13030 20202 13082
rect 20202 13030 20212 13082
rect 20236 13030 20266 13082
rect 20266 13030 20278 13082
rect 20278 13030 20292 13082
rect 20316 13030 20330 13082
rect 20330 13030 20342 13082
rect 20342 13030 20372 13082
rect 20396 13030 20406 13082
rect 20406 13030 20452 13082
rect 20156 13028 20212 13030
rect 20236 13028 20292 13030
rect 20316 13028 20372 13030
rect 20396 13028 20452 13030
rect 20156 11994 20212 11996
rect 20236 11994 20292 11996
rect 20316 11994 20372 11996
rect 20396 11994 20452 11996
rect 20156 11942 20202 11994
rect 20202 11942 20212 11994
rect 20236 11942 20266 11994
rect 20266 11942 20278 11994
rect 20278 11942 20292 11994
rect 20316 11942 20330 11994
rect 20330 11942 20342 11994
rect 20342 11942 20372 11994
rect 20396 11942 20406 11994
rect 20406 11942 20452 11994
rect 20156 11940 20212 11942
rect 20236 11940 20292 11942
rect 20316 11940 20372 11942
rect 20396 11940 20452 11942
rect 20156 10906 20212 10908
rect 20236 10906 20292 10908
rect 20316 10906 20372 10908
rect 20396 10906 20452 10908
rect 20156 10854 20202 10906
rect 20202 10854 20212 10906
rect 20236 10854 20266 10906
rect 20266 10854 20278 10906
rect 20278 10854 20292 10906
rect 20316 10854 20330 10906
rect 20330 10854 20342 10906
rect 20342 10854 20372 10906
rect 20396 10854 20406 10906
rect 20406 10854 20452 10906
rect 20156 10852 20212 10854
rect 20236 10852 20292 10854
rect 20316 10852 20372 10854
rect 20396 10852 20452 10854
rect 20156 9818 20212 9820
rect 20236 9818 20292 9820
rect 20316 9818 20372 9820
rect 20396 9818 20452 9820
rect 20156 9766 20202 9818
rect 20202 9766 20212 9818
rect 20236 9766 20266 9818
rect 20266 9766 20278 9818
rect 20278 9766 20292 9818
rect 20316 9766 20330 9818
rect 20330 9766 20342 9818
rect 20342 9766 20372 9818
rect 20396 9766 20406 9818
rect 20406 9766 20452 9818
rect 20156 9764 20212 9766
rect 20236 9764 20292 9766
rect 20316 9764 20372 9766
rect 20396 9764 20452 9766
rect 20156 8730 20212 8732
rect 20236 8730 20292 8732
rect 20316 8730 20372 8732
rect 20396 8730 20452 8732
rect 20156 8678 20202 8730
rect 20202 8678 20212 8730
rect 20236 8678 20266 8730
rect 20266 8678 20278 8730
rect 20278 8678 20292 8730
rect 20316 8678 20330 8730
rect 20330 8678 20342 8730
rect 20342 8678 20372 8730
rect 20396 8678 20406 8730
rect 20406 8678 20452 8730
rect 20156 8676 20212 8678
rect 20236 8676 20292 8678
rect 20316 8676 20372 8678
rect 20396 8676 20452 8678
rect 22556 17978 22612 17980
rect 22636 17978 22692 17980
rect 22716 17978 22772 17980
rect 22796 17978 22852 17980
rect 22556 17926 22602 17978
rect 22602 17926 22612 17978
rect 22636 17926 22666 17978
rect 22666 17926 22678 17978
rect 22678 17926 22692 17978
rect 22716 17926 22730 17978
rect 22730 17926 22742 17978
rect 22742 17926 22772 17978
rect 22796 17926 22806 17978
rect 22806 17926 22852 17978
rect 22556 17924 22612 17926
rect 22636 17924 22692 17926
rect 22716 17924 22772 17926
rect 22796 17924 22852 17926
rect 24956 19610 25012 19612
rect 25036 19610 25092 19612
rect 25116 19610 25172 19612
rect 25196 19610 25252 19612
rect 24956 19558 25002 19610
rect 25002 19558 25012 19610
rect 25036 19558 25066 19610
rect 25066 19558 25078 19610
rect 25078 19558 25092 19610
rect 25116 19558 25130 19610
rect 25130 19558 25142 19610
rect 25142 19558 25172 19610
rect 25196 19558 25206 19610
rect 25206 19558 25252 19610
rect 24956 19556 25012 19558
rect 25036 19556 25092 19558
rect 25116 19556 25172 19558
rect 25196 19556 25252 19558
rect 24956 18522 25012 18524
rect 25036 18522 25092 18524
rect 25116 18522 25172 18524
rect 25196 18522 25252 18524
rect 24956 18470 25002 18522
rect 25002 18470 25012 18522
rect 25036 18470 25066 18522
rect 25066 18470 25078 18522
rect 25078 18470 25092 18522
rect 25116 18470 25130 18522
rect 25130 18470 25142 18522
rect 25142 18470 25172 18522
rect 25196 18470 25206 18522
rect 25206 18470 25252 18522
rect 24956 18468 25012 18470
rect 25036 18468 25092 18470
rect 25116 18468 25172 18470
rect 25196 18468 25252 18470
rect 22556 16890 22612 16892
rect 22636 16890 22692 16892
rect 22716 16890 22772 16892
rect 22796 16890 22852 16892
rect 22556 16838 22602 16890
rect 22602 16838 22612 16890
rect 22636 16838 22666 16890
rect 22666 16838 22678 16890
rect 22678 16838 22692 16890
rect 22716 16838 22730 16890
rect 22730 16838 22742 16890
rect 22742 16838 22772 16890
rect 22796 16838 22806 16890
rect 22806 16838 22852 16890
rect 22556 16836 22612 16838
rect 22636 16836 22692 16838
rect 22716 16836 22772 16838
rect 22796 16836 22852 16838
rect 22556 15802 22612 15804
rect 22636 15802 22692 15804
rect 22716 15802 22772 15804
rect 22796 15802 22852 15804
rect 22556 15750 22602 15802
rect 22602 15750 22612 15802
rect 22636 15750 22666 15802
rect 22666 15750 22678 15802
rect 22678 15750 22692 15802
rect 22716 15750 22730 15802
rect 22730 15750 22742 15802
rect 22742 15750 22772 15802
rect 22796 15750 22806 15802
rect 22806 15750 22852 15802
rect 22556 15748 22612 15750
rect 22636 15748 22692 15750
rect 22716 15748 22772 15750
rect 22796 15748 22852 15750
rect 24956 17434 25012 17436
rect 25036 17434 25092 17436
rect 25116 17434 25172 17436
rect 25196 17434 25252 17436
rect 24956 17382 25002 17434
rect 25002 17382 25012 17434
rect 25036 17382 25066 17434
rect 25066 17382 25078 17434
rect 25078 17382 25092 17434
rect 25116 17382 25130 17434
rect 25130 17382 25142 17434
rect 25142 17382 25172 17434
rect 25196 17382 25206 17434
rect 25206 17382 25252 17434
rect 24956 17380 25012 17382
rect 25036 17380 25092 17382
rect 25116 17380 25172 17382
rect 25196 17380 25252 17382
rect 27356 22330 27412 22332
rect 27436 22330 27492 22332
rect 27516 22330 27572 22332
rect 27596 22330 27652 22332
rect 27356 22278 27402 22330
rect 27402 22278 27412 22330
rect 27436 22278 27466 22330
rect 27466 22278 27478 22330
rect 27478 22278 27492 22330
rect 27516 22278 27530 22330
rect 27530 22278 27542 22330
rect 27542 22278 27572 22330
rect 27596 22278 27606 22330
rect 27606 22278 27652 22330
rect 27356 22276 27412 22278
rect 27436 22276 27492 22278
rect 27516 22276 27572 22278
rect 27596 22276 27652 22278
rect 28354 25880 28410 25936
rect 28354 23468 28356 23488
rect 28356 23468 28408 23488
rect 28408 23468 28410 23488
rect 28354 23432 28410 23468
rect 27356 21242 27412 21244
rect 27436 21242 27492 21244
rect 27516 21242 27572 21244
rect 27596 21242 27652 21244
rect 27356 21190 27402 21242
rect 27402 21190 27412 21242
rect 27436 21190 27466 21242
rect 27466 21190 27478 21242
rect 27478 21190 27492 21242
rect 27516 21190 27530 21242
rect 27530 21190 27542 21242
rect 27542 21190 27572 21242
rect 27596 21190 27606 21242
rect 27606 21190 27652 21242
rect 27356 21188 27412 21190
rect 27436 21188 27492 21190
rect 27516 21188 27572 21190
rect 27596 21188 27652 21190
rect 28354 20984 28410 21040
rect 27356 20154 27412 20156
rect 27436 20154 27492 20156
rect 27516 20154 27572 20156
rect 27596 20154 27652 20156
rect 27356 20102 27402 20154
rect 27402 20102 27412 20154
rect 27436 20102 27466 20154
rect 27466 20102 27478 20154
rect 27478 20102 27492 20154
rect 27516 20102 27530 20154
rect 27530 20102 27542 20154
rect 27542 20102 27572 20154
rect 27596 20102 27606 20154
rect 27606 20102 27652 20154
rect 27356 20100 27412 20102
rect 27436 20100 27492 20102
rect 27516 20100 27572 20102
rect 27596 20100 27652 20102
rect 27356 19066 27412 19068
rect 27436 19066 27492 19068
rect 27516 19066 27572 19068
rect 27596 19066 27652 19068
rect 27356 19014 27402 19066
rect 27402 19014 27412 19066
rect 27436 19014 27466 19066
rect 27466 19014 27478 19066
rect 27478 19014 27492 19066
rect 27516 19014 27530 19066
rect 27530 19014 27542 19066
rect 27542 19014 27572 19066
rect 27596 19014 27606 19066
rect 27606 19014 27652 19066
rect 27356 19012 27412 19014
rect 27436 19012 27492 19014
rect 27516 19012 27572 19014
rect 27596 19012 27652 19014
rect 24956 16346 25012 16348
rect 25036 16346 25092 16348
rect 25116 16346 25172 16348
rect 25196 16346 25252 16348
rect 24956 16294 25002 16346
rect 25002 16294 25012 16346
rect 25036 16294 25066 16346
rect 25066 16294 25078 16346
rect 25078 16294 25092 16346
rect 25116 16294 25130 16346
rect 25130 16294 25142 16346
rect 25142 16294 25172 16346
rect 25196 16294 25206 16346
rect 25206 16294 25252 16346
rect 24956 16292 25012 16294
rect 25036 16292 25092 16294
rect 25116 16292 25172 16294
rect 25196 16292 25252 16294
rect 24956 15258 25012 15260
rect 25036 15258 25092 15260
rect 25116 15258 25172 15260
rect 25196 15258 25252 15260
rect 24956 15206 25002 15258
rect 25002 15206 25012 15258
rect 25036 15206 25066 15258
rect 25066 15206 25078 15258
rect 25078 15206 25092 15258
rect 25116 15206 25130 15258
rect 25130 15206 25142 15258
rect 25142 15206 25172 15258
rect 25196 15206 25206 15258
rect 25206 15206 25252 15258
rect 24956 15204 25012 15206
rect 25036 15204 25092 15206
rect 25116 15204 25172 15206
rect 25196 15204 25252 15206
rect 22556 14714 22612 14716
rect 22636 14714 22692 14716
rect 22716 14714 22772 14716
rect 22796 14714 22852 14716
rect 22556 14662 22602 14714
rect 22602 14662 22612 14714
rect 22636 14662 22666 14714
rect 22666 14662 22678 14714
rect 22678 14662 22692 14714
rect 22716 14662 22730 14714
rect 22730 14662 22742 14714
rect 22742 14662 22772 14714
rect 22796 14662 22806 14714
rect 22806 14662 22852 14714
rect 22556 14660 22612 14662
rect 22636 14660 22692 14662
rect 22716 14660 22772 14662
rect 22796 14660 22852 14662
rect 22556 13626 22612 13628
rect 22636 13626 22692 13628
rect 22716 13626 22772 13628
rect 22796 13626 22852 13628
rect 22556 13574 22602 13626
rect 22602 13574 22612 13626
rect 22636 13574 22666 13626
rect 22666 13574 22678 13626
rect 22678 13574 22692 13626
rect 22716 13574 22730 13626
rect 22730 13574 22742 13626
rect 22742 13574 22772 13626
rect 22796 13574 22806 13626
rect 22806 13574 22852 13626
rect 22556 13572 22612 13574
rect 22636 13572 22692 13574
rect 22716 13572 22772 13574
rect 22796 13572 22852 13574
rect 22556 12538 22612 12540
rect 22636 12538 22692 12540
rect 22716 12538 22772 12540
rect 22796 12538 22852 12540
rect 22556 12486 22602 12538
rect 22602 12486 22612 12538
rect 22636 12486 22666 12538
rect 22666 12486 22678 12538
rect 22678 12486 22692 12538
rect 22716 12486 22730 12538
rect 22730 12486 22742 12538
rect 22742 12486 22772 12538
rect 22796 12486 22806 12538
rect 22806 12486 22852 12538
rect 22556 12484 22612 12486
rect 22636 12484 22692 12486
rect 22716 12484 22772 12486
rect 22796 12484 22852 12486
rect 24956 14170 25012 14172
rect 25036 14170 25092 14172
rect 25116 14170 25172 14172
rect 25196 14170 25252 14172
rect 24956 14118 25002 14170
rect 25002 14118 25012 14170
rect 25036 14118 25066 14170
rect 25066 14118 25078 14170
rect 25078 14118 25092 14170
rect 25116 14118 25130 14170
rect 25130 14118 25142 14170
rect 25142 14118 25172 14170
rect 25196 14118 25206 14170
rect 25206 14118 25252 14170
rect 24956 14116 25012 14118
rect 25036 14116 25092 14118
rect 25116 14116 25172 14118
rect 25196 14116 25252 14118
rect 27356 17978 27412 17980
rect 27436 17978 27492 17980
rect 27516 17978 27572 17980
rect 27596 17978 27652 17980
rect 27356 17926 27402 17978
rect 27402 17926 27412 17978
rect 27436 17926 27466 17978
rect 27466 17926 27478 17978
rect 27478 17926 27492 17978
rect 27516 17926 27530 17978
rect 27530 17926 27542 17978
rect 27542 17926 27572 17978
rect 27596 17926 27606 17978
rect 27606 17926 27652 17978
rect 27356 17924 27412 17926
rect 27436 17924 27492 17926
rect 27516 17924 27572 17926
rect 27596 17924 27652 17926
rect 28354 18572 28356 18592
rect 28356 18572 28408 18592
rect 28408 18572 28410 18592
rect 28354 18536 28410 18572
rect 27356 16890 27412 16892
rect 27436 16890 27492 16892
rect 27516 16890 27572 16892
rect 27596 16890 27652 16892
rect 27356 16838 27402 16890
rect 27402 16838 27412 16890
rect 27436 16838 27466 16890
rect 27466 16838 27478 16890
rect 27478 16838 27492 16890
rect 27516 16838 27530 16890
rect 27530 16838 27542 16890
rect 27542 16838 27572 16890
rect 27596 16838 27606 16890
rect 27606 16838 27652 16890
rect 27356 16836 27412 16838
rect 27436 16836 27492 16838
rect 27516 16836 27572 16838
rect 27596 16836 27652 16838
rect 27356 15802 27412 15804
rect 27436 15802 27492 15804
rect 27516 15802 27572 15804
rect 27596 15802 27652 15804
rect 27356 15750 27402 15802
rect 27402 15750 27412 15802
rect 27436 15750 27466 15802
rect 27466 15750 27478 15802
rect 27478 15750 27492 15802
rect 27516 15750 27530 15802
rect 27530 15750 27542 15802
rect 27542 15750 27572 15802
rect 27596 15750 27606 15802
rect 27606 15750 27652 15802
rect 27356 15748 27412 15750
rect 27436 15748 27492 15750
rect 27516 15748 27572 15750
rect 27596 15748 27652 15750
rect 28354 16088 28410 16144
rect 27356 14714 27412 14716
rect 27436 14714 27492 14716
rect 27516 14714 27572 14716
rect 27596 14714 27652 14716
rect 27356 14662 27402 14714
rect 27402 14662 27412 14714
rect 27436 14662 27466 14714
rect 27466 14662 27478 14714
rect 27478 14662 27492 14714
rect 27516 14662 27530 14714
rect 27530 14662 27542 14714
rect 27542 14662 27572 14714
rect 27596 14662 27606 14714
rect 27606 14662 27652 14714
rect 27356 14660 27412 14662
rect 27436 14660 27492 14662
rect 27516 14660 27572 14662
rect 27596 14660 27652 14662
rect 24956 13082 25012 13084
rect 25036 13082 25092 13084
rect 25116 13082 25172 13084
rect 25196 13082 25252 13084
rect 24956 13030 25002 13082
rect 25002 13030 25012 13082
rect 25036 13030 25066 13082
rect 25066 13030 25078 13082
rect 25078 13030 25092 13082
rect 25116 13030 25130 13082
rect 25130 13030 25142 13082
rect 25142 13030 25172 13082
rect 25196 13030 25206 13082
rect 25206 13030 25252 13082
rect 24956 13028 25012 13030
rect 25036 13028 25092 13030
rect 25116 13028 25172 13030
rect 25196 13028 25252 13030
rect 27356 13626 27412 13628
rect 27436 13626 27492 13628
rect 27516 13626 27572 13628
rect 27596 13626 27652 13628
rect 27356 13574 27402 13626
rect 27402 13574 27412 13626
rect 27436 13574 27466 13626
rect 27466 13574 27478 13626
rect 27478 13574 27492 13626
rect 27516 13574 27530 13626
rect 27530 13574 27542 13626
rect 27542 13574 27572 13626
rect 27596 13574 27606 13626
rect 27606 13574 27652 13626
rect 27356 13572 27412 13574
rect 27436 13572 27492 13574
rect 27516 13572 27572 13574
rect 27596 13572 27652 13574
rect 28354 13676 28356 13696
rect 28356 13676 28408 13696
rect 28408 13676 28410 13696
rect 28354 13640 28410 13676
rect 22556 11450 22612 11452
rect 22636 11450 22692 11452
rect 22716 11450 22772 11452
rect 22796 11450 22852 11452
rect 22556 11398 22602 11450
rect 22602 11398 22612 11450
rect 22636 11398 22666 11450
rect 22666 11398 22678 11450
rect 22678 11398 22692 11450
rect 22716 11398 22730 11450
rect 22730 11398 22742 11450
rect 22742 11398 22772 11450
rect 22796 11398 22806 11450
rect 22806 11398 22852 11450
rect 22556 11396 22612 11398
rect 22636 11396 22692 11398
rect 22716 11396 22772 11398
rect 22796 11396 22852 11398
rect 22556 10362 22612 10364
rect 22636 10362 22692 10364
rect 22716 10362 22772 10364
rect 22796 10362 22852 10364
rect 22556 10310 22602 10362
rect 22602 10310 22612 10362
rect 22636 10310 22666 10362
rect 22666 10310 22678 10362
rect 22678 10310 22692 10362
rect 22716 10310 22730 10362
rect 22730 10310 22742 10362
rect 22742 10310 22772 10362
rect 22796 10310 22806 10362
rect 22806 10310 22852 10362
rect 22556 10308 22612 10310
rect 22636 10308 22692 10310
rect 22716 10308 22772 10310
rect 22796 10308 22852 10310
rect 24956 11994 25012 11996
rect 25036 11994 25092 11996
rect 25116 11994 25172 11996
rect 25196 11994 25252 11996
rect 24956 11942 25002 11994
rect 25002 11942 25012 11994
rect 25036 11942 25066 11994
rect 25066 11942 25078 11994
rect 25078 11942 25092 11994
rect 25116 11942 25130 11994
rect 25130 11942 25142 11994
rect 25142 11942 25172 11994
rect 25196 11942 25206 11994
rect 25206 11942 25252 11994
rect 24956 11940 25012 11942
rect 25036 11940 25092 11942
rect 25116 11940 25172 11942
rect 25196 11940 25252 11942
rect 27356 12538 27412 12540
rect 27436 12538 27492 12540
rect 27516 12538 27572 12540
rect 27596 12538 27652 12540
rect 27356 12486 27402 12538
rect 27402 12486 27412 12538
rect 27436 12486 27466 12538
rect 27466 12486 27478 12538
rect 27478 12486 27492 12538
rect 27516 12486 27530 12538
rect 27530 12486 27542 12538
rect 27542 12486 27572 12538
rect 27596 12486 27606 12538
rect 27606 12486 27652 12538
rect 27356 12484 27412 12486
rect 27436 12484 27492 12486
rect 27516 12484 27572 12486
rect 27596 12484 27652 12486
rect 24956 10906 25012 10908
rect 25036 10906 25092 10908
rect 25116 10906 25172 10908
rect 25196 10906 25252 10908
rect 24956 10854 25002 10906
rect 25002 10854 25012 10906
rect 25036 10854 25066 10906
rect 25066 10854 25078 10906
rect 25078 10854 25092 10906
rect 25116 10854 25130 10906
rect 25130 10854 25142 10906
rect 25142 10854 25172 10906
rect 25196 10854 25206 10906
rect 25206 10854 25252 10906
rect 24956 10852 25012 10854
rect 25036 10852 25092 10854
rect 25116 10852 25172 10854
rect 25196 10852 25252 10854
rect 22556 9274 22612 9276
rect 22636 9274 22692 9276
rect 22716 9274 22772 9276
rect 22796 9274 22852 9276
rect 22556 9222 22602 9274
rect 22602 9222 22612 9274
rect 22636 9222 22666 9274
rect 22666 9222 22678 9274
rect 22678 9222 22692 9274
rect 22716 9222 22730 9274
rect 22730 9222 22742 9274
rect 22742 9222 22772 9274
rect 22796 9222 22806 9274
rect 22806 9222 22852 9274
rect 22556 9220 22612 9222
rect 22636 9220 22692 9222
rect 22716 9220 22772 9222
rect 22796 9220 22852 9222
rect 20156 7642 20212 7644
rect 20236 7642 20292 7644
rect 20316 7642 20372 7644
rect 20396 7642 20452 7644
rect 20156 7590 20202 7642
rect 20202 7590 20212 7642
rect 20236 7590 20266 7642
rect 20266 7590 20278 7642
rect 20278 7590 20292 7642
rect 20316 7590 20330 7642
rect 20330 7590 20342 7642
rect 20342 7590 20372 7642
rect 20396 7590 20406 7642
rect 20406 7590 20452 7642
rect 20156 7588 20212 7590
rect 20236 7588 20292 7590
rect 20316 7588 20372 7590
rect 20396 7588 20452 7590
rect 22556 8186 22612 8188
rect 22636 8186 22692 8188
rect 22716 8186 22772 8188
rect 22796 8186 22852 8188
rect 22556 8134 22602 8186
rect 22602 8134 22612 8186
rect 22636 8134 22666 8186
rect 22666 8134 22678 8186
rect 22678 8134 22692 8186
rect 22716 8134 22730 8186
rect 22730 8134 22742 8186
rect 22742 8134 22772 8186
rect 22796 8134 22806 8186
rect 22806 8134 22852 8186
rect 22556 8132 22612 8134
rect 22636 8132 22692 8134
rect 22716 8132 22772 8134
rect 22796 8132 22852 8134
rect 20156 6554 20212 6556
rect 20236 6554 20292 6556
rect 20316 6554 20372 6556
rect 20396 6554 20452 6556
rect 20156 6502 20202 6554
rect 20202 6502 20212 6554
rect 20236 6502 20266 6554
rect 20266 6502 20278 6554
rect 20278 6502 20292 6554
rect 20316 6502 20330 6554
rect 20330 6502 20342 6554
rect 20342 6502 20372 6554
rect 20396 6502 20406 6554
rect 20406 6502 20452 6554
rect 20156 6500 20212 6502
rect 20236 6500 20292 6502
rect 20316 6500 20372 6502
rect 20396 6500 20452 6502
rect 22556 7098 22612 7100
rect 22636 7098 22692 7100
rect 22716 7098 22772 7100
rect 22796 7098 22852 7100
rect 22556 7046 22602 7098
rect 22602 7046 22612 7098
rect 22636 7046 22666 7098
rect 22666 7046 22678 7098
rect 22678 7046 22692 7098
rect 22716 7046 22730 7098
rect 22730 7046 22742 7098
rect 22742 7046 22772 7098
rect 22796 7046 22806 7098
rect 22806 7046 22852 7098
rect 22556 7044 22612 7046
rect 22636 7044 22692 7046
rect 22716 7044 22772 7046
rect 22796 7044 22852 7046
rect 20156 5466 20212 5468
rect 20236 5466 20292 5468
rect 20316 5466 20372 5468
rect 20396 5466 20452 5468
rect 20156 5414 20202 5466
rect 20202 5414 20212 5466
rect 20236 5414 20266 5466
rect 20266 5414 20278 5466
rect 20278 5414 20292 5466
rect 20316 5414 20330 5466
rect 20330 5414 20342 5466
rect 20342 5414 20372 5466
rect 20396 5414 20406 5466
rect 20406 5414 20452 5466
rect 20156 5412 20212 5414
rect 20236 5412 20292 5414
rect 20316 5412 20372 5414
rect 20396 5412 20452 5414
rect 20156 4378 20212 4380
rect 20236 4378 20292 4380
rect 20316 4378 20372 4380
rect 20396 4378 20452 4380
rect 20156 4326 20202 4378
rect 20202 4326 20212 4378
rect 20236 4326 20266 4378
rect 20266 4326 20278 4378
rect 20278 4326 20292 4378
rect 20316 4326 20330 4378
rect 20330 4326 20342 4378
rect 20342 4326 20372 4378
rect 20396 4326 20406 4378
rect 20406 4326 20452 4378
rect 20156 4324 20212 4326
rect 20236 4324 20292 4326
rect 20316 4324 20372 4326
rect 20396 4324 20452 4326
rect 22556 6010 22612 6012
rect 22636 6010 22692 6012
rect 22716 6010 22772 6012
rect 22796 6010 22852 6012
rect 22556 5958 22602 6010
rect 22602 5958 22612 6010
rect 22636 5958 22666 6010
rect 22666 5958 22678 6010
rect 22678 5958 22692 6010
rect 22716 5958 22730 6010
rect 22730 5958 22742 6010
rect 22742 5958 22772 6010
rect 22796 5958 22806 6010
rect 22806 5958 22852 6010
rect 22556 5956 22612 5958
rect 22636 5956 22692 5958
rect 22716 5956 22772 5958
rect 22796 5956 22852 5958
rect 22556 4922 22612 4924
rect 22636 4922 22692 4924
rect 22716 4922 22772 4924
rect 22796 4922 22852 4924
rect 22556 4870 22602 4922
rect 22602 4870 22612 4922
rect 22636 4870 22666 4922
rect 22666 4870 22678 4922
rect 22678 4870 22692 4922
rect 22716 4870 22730 4922
rect 22730 4870 22742 4922
rect 22742 4870 22772 4922
rect 22796 4870 22806 4922
rect 22806 4870 22852 4922
rect 22556 4868 22612 4870
rect 22636 4868 22692 4870
rect 22716 4868 22772 4870
rect 22796 4868 22852 4870
rect 24956 9818 25012 9820
rect 25036 9818 25092 9820
rect 25116 9818 25172 9820
rect 25196 9818 25252 9820
rect 24956 9766 25002 9818
rect 25002 9766 25012 9818
rect 25036 9766 25066 9818
rect 25066 9766 25078 9818
rect 25078 9766 25092 9818
rect 25116 9766 25130 9818
rect 25130 9766 25142 9818
rect 25142 9766 25172 9818
rect 25196 9766 25206 9818
rect 25206 9766 25252 9818
rect 24956 9764 25012 9766
rect 25036 9764 25092 9766
rect 25116 9764 25172 9766
rect 25196 9764 25252 9766
rect 27356 11450 27412 11452
rect 27436 11450 27492 11452
rect 27516 11450 27572 11452
rect 27596 11450 27652 11452
rect 27356 11398 27402 11450
rect 27402 11398 27412 11450
rect 27436 11398 27466 11450
rect 27466 11398 27478 11450
rect 27478 11398 27492 11450
rect 27516 11398 27530 11450
rect 27530 11398 27542 11450
rect 27542 11398 27572 11450
rect 27596 11398 27606 11450
rect 27606 11398 27652 11450
rect 27356 11396 27412 11398
rect 27436 11396 27492 11398
rect 27516 11396 27572 11398
rect 27596 11396 27652 11398
rect 24956 8730 25012 8732
rect 25036 8730 25092 8732
rect 25116 8730 25172 8732
rect 25196 8730 25252 8732
rect 24956 8678 25002 8730
rect 25002 8678 25012 8730
rect 25036 8678 25066 8730
rect 25066 8678 25078 8730
rect 25078 8678 25092 8730
rect 25116 8678 25130 8730
rect 25130 8678 25142 8730
rect 25142 8678 25172 8730
rect 25196 8678 25206 8730
rect 25206 8678 25252 8730
rect 24956 8676 25012 8678
rect 25036 8676 25092 8678
rect 25116 8676 25172 8678
rect 25196 8676 25252 8678
rect 24956 7642 25012 7644
rect 25036 7642 25092 7644
rect 25116 7642 25172 7644
rect 25196 7642 25252 7644
rect 24956 7590 25002 7642
rect 25002 7590 25012 7642
rect 25036 7590 25066 7642
rect 25066 7590 25078 7642
rect 25078 7590 25092 7642
rect 25116 7590 25130 7642
rect 25130 7590 25142 7642
rect 25142 7590 25172 7642
rect 25196 7590 25206 7642
rect 25206 7590 25252 7642
rect 24956 7588 25012 7590
rect 25036 7588 25092 7590
rect 25116 7588 25172 7590
rect 25196 7588 25252 7590
rect 27356 10362 27412 10364
rect 27436 10362 27492 10364
rect 27516 10362 27572 10364
rect 27596 10362 27652 10364
rect 27356 10310 27402 10362
rect 27402 10310 27412 10362
rect 27436 10310 27466 10362
rect 27466 10310 27478 10362
rect 27478 10310 27492 10362
rect 27516 10310 27530 10362
rect 27530 10310 27542 10362
rect 27542 10310 27572 10362
rect 27596 10310 27606 10362
rect 27606 10310 27652 10362
rect 27356 10308 27412 10310
rect 27436 10308 27492 10310
rect 27516 10308 27572 10310
rect 27596 10308 27652 10310
rect 27356 9274 27412 9276
rect 27436 9274 27492 9276
rect 27516 9274 27572 9276
rect 27596 9274 27652 9276
rect 27356 9222 27402 9274
rect 27402 9222 27412 9274
rect 27436 9222 27466 9274
rect 27466 9222 27478 9274
rect 27478 9222 27492 9274
rect 27516 9222 27530 9274
rect 27530 9222 27542 9274
rect 27542 9222 27572 9274
rect 27596 9222 27606 9274
rect 27606 9222 27652 9274
rect 27356 9220 27412 9222
rect 27436 9220 27492 9222
rect 27516 9220 27572 9222
rect 27596 9220 27652 9222
rect 28354 11192 28410 11248
rect 27356 8186 27412 8188
rect 27436 8186 27492 8188
rect 27516 8186 27572 8188
rect 27596 8186 27652 8188
rect 27356 8134 27402 8186
rect 27402 8134 27412 8186
rect 27436 8134 27466 8186
rect 27466 8134 27478 8186
rect 27478 8134 27492 8186
rect 27516 8134 27530 8186
rect 27530 8134 27542 8186
rect 27542 8134 27572 8186
rect 27596 8134 27606 8186
rect 27606 8134 27652 8186
rect 27356 8132 27412 8134
rect 27436 8132 27492 8134
rect 27516 8132 27572 8134
rect 27596 8132 27652 8134
rect 27356 7098 27412 7100
rect 27436 7098 27492 7100
rect 27516 7098 27572 7100
rect 27596 7098 27652 7100
rect 27356 7046 27402 7098
rect 27402 7046 27412 7098
rect 27436 7046 27466 7098
rect 27466 7046 27478 7098
rect 27478 7046 27492 7098
rect 27516 7046 27530 7098
rect 27530 7046 27542 7098
rect 27542 7046 27572 7098
rect 27596 7046 27606 7098
rect 27606 7046 27652 7098
rect 27356 7044 27412 7046
rect 27436 7044 27492 7046
rect 27516 7044 27572 7046
rect 27596 7044 27652 7046
rect 24956 6554 25012 6556
rect 25036 6554 25092 6556
rect 25116 6554 25172 6556
rect 25196 6554 25252 6556
rect 24956 6502 25002 6554
rect 25002 6502 25012 6554
rect 25036 6502 25066 6554
rect 25066 6502 25078 6554
rect 25078 6502 25092 6554
rect 25116 6502 25130 6554
rect 25130 6502 25142 6554
rect 25142 6502 25172 6554
rect 25196 6502 25206 6554
rect 25206 6502 25252 6554
rect 24956 6500 25012 6502
rect 25036 6500 25092 6502
rect 25116 6500 25172 6502
rect 25196 6500 25252 6502
rect 28354 8744 28410 8800
rect 27356 6010 27412 6012
rect 27436 6010 27492 6012
rect 27516 6010 27572 6012
rect 27596 6010 27652 6012
rect 27356 5958 27402 6010
rect 27402 5958 27412 6010
rect 27436 5958 27466 6010
rect 27466 5958 27478 6010
rect 27478 5958 27492 6010
rect 27516 5958 27530 6010
rect 27530 5958 27542 6010
rect 27542 5958 27572 6010
rect 27596 5958 27606 6010
rect 27606 5958 27652 6010
rect 27356 5956 27412 5958
rect 27436 5956 27492 5958
rect 27516 5956 27572 5958
rect 27596 5956 27652 5958
rect 24956 5466 25012 5468
rect 25036 5466 25092 5468
rect 25116 5466 25172 5468
rect 25196 5466 25252 5468
rect 24956 5414 25002 5466
rect 25002 5414 25012 5466
rect 25036 5414 25066 5466
rect 25066 5414 25078 5466
rect 25078 5414 25092 5466
rect 25116 5414 25130 5466
rect 25130 5414 25142 5466
rect 25142 5414 25172 5466
rect 25196 5414 25206 5466
rect 25206 5414 25252 5466
rect 24956 5412 25012 5414
rect 25036 5412 25092 5414
rect 25116 5412 25172 5414
rect 25196 5412 25252 5414
rect 27356 4922 27412 4924
rect 27436 4922 27492 4924
rect 27516 4922 27572 4924
rect 27596 4922 27652 4924
rect 27356 4870 27402 4922
rect 27402 4870 27412 4922
rect 27436 4870 27466 4922
rect 27466 4870 27478 4922
rect 27478 4870 27492 4922
rect 27516 4870 27530 4922
rect 27530 4870 27542 4922
rect 27542 4870 27572 4922
rect 27596 4870 27606 4922
rect 27606 4870 27652 4922
rect 27356 4868 27412 4870
rect 27436 4868 27492 4870
rect 27516 4868 27572 4870
rect 27596 4868 27652 4870
rect 22556 3834 22612 3836
rect 22636 3834 22692 3836
rect 22716 3834 22772 3836
rect 22796 3834 22852 3836
rect 22556 3782 22602 3834
rect 22602 3782 22612 3834
rect 22636 3782 22666 3834
rect 22666 3782 22678 3834
rect 22678 3782 22692 3834
rect 22716 3782 22730 3834
rect 22730 3782 22742 3834
rect 22742 3782 22772 3834
rect 22796 3782 22806 3834
rect 22806 3782 22852 3834
rect 22556 3780 22612 3782
rect 22636 3780 22692 3782
rect 22716 3780 22772 3782
rect 22796 3780 22852 3782
rect 20156 3290 20212 3292
rect 20236 3290 20292 3292
rect 20316 3290 20372 3292
rect 20396 3290 20452 3292
rect 20156 3238 20202 3290
rect 20202 3238 20212 3290
rect 20236 3238 20266 3290
rect 20266 3238 20278 3290
rect 20278 3238 20292 3290
rect 20316 3238 20330 3290
rect 20330 3238 20342 3290
rect 20342 3238 20372 3290
rect 20396 3238 20406 3290
rect 20406 3238 20452 3290
rect 20156 3236 20212 3238
rect 20236 3236 20292 3238
rect 20316 3236 20372 3238
rect 20396 3236 20452 3238
rect 24956 4378 25012 4380
rect 25036 4378 25092 4380
rect 25116 4378 25172 4380
rect 25196 4378 25252 4380
rect 24956 4326 25002 4378
rect 25002 4326 25012 4378
rect 25036 4326 25066 4378
rect 25066 4326 25078 4378
rect 25078 4326 25092 4378
rect 25116 4326 25130 4378
rect 25130 4326 25142 4378
rect 25142 4326 25172 4378
rect 25196 4326 25206 4378
rect 25206 4326 25252 4378
rect 24956 4324 25012 4326
rect 25036 4324 25092 4326
rect 25116 4324 25172 4326
rect 25196 4324 25252 4326
rect 24956 3290 25012 3292
rect 25036 3290 25092 3292
rect 25116 3290 25172 3292
rect 25196 3290 25252 3292
rect 24956 3238 25002 3290
rect 25002 3238 25012 3290
rect 25036 3238 25066 3290
rect 25066 3238 25078 3290
rect 25078 3238 25092 3290
rect 25116 3238 25130 3290
rect 25130 3238 25142 3290
rect 25142 3238 25172 3290
rect 25196 3238 25206 3290
rect 25206 3238 25252 3290
rect 24956 3236 25012 3238
rect 25036 3236 25092 3238
rect 25116 3236 25172 3238
rect 25196 3236 25252 3238
rect 28354 6296 28410 6352
rect 27356 3834 27412 3836
rect 27436 3834 27492 3836
rect 27516 3834 27572 3836
rect 27596 3834 27652 3836
rect 27356 3782 27402 3834
rect 27402 3782 27412 3834
rect 27436 3782 27466 3834
rect 27466 3782 27478 3834
rect 27478 3782 27492 3834
rect 27516 3782 27530 3834
rect 27530 3782 27542 3834
rect 27542 3782 27572 3834
rect 27596 3782 27606 3834
rect 27606 3782 27652 3834
rect 27356 3780 27412 3782
rect 27436 3780 27492 3782
rect 27516 3780 27572 3782
rect 27596 3780 27652 3782
rect 28354 3848 28410 3904
rect 22556 2746 22612 2748
rect 22636 2746 22692 2748
rect 22716 2746 22772 2748
rect 22796 2746 22852 2748
rect 22556 2694 22602 2746
rect 22602 2694 22612 2746
rect 22636 2694 22666 2746
rect 22666 2694 22678 2746
rect 22678 2694 22692 2746
rect 22716 2694 22730 2746
rect 22730 2694 22742 2746
rect 22742 2694 22772 2746
rect 22796 2694 22806 2746
rect 22806 2694 22852 2746
rect 22556 2692 22612 2694
rect 22636 2692 22692 2694
rect 22716 2692 22772 2694
rect 22796 2692 22852 2694
rect 27356 2746 27412 2748
rect 27436 2746 27492 2748
rect 27516 2746 27572 2748
rect 27596 2746 27652 2748
rect 27356 2694 27402 2746
rect 27402 2694 27412 2746
rect 27436 2694 27466 2746
rect 27466 2694 27478 2746
rect 27478 2694 27492 2746
rect 27516 2694 27530 2746
rect 27530 2694 27542 2746
rect 27542 2694 27572 2746
rect 27596 2694 27606 2746
rect 27606 2694 27652 2746
rect 27356 2692 27412 2694
rect 27436 2692 27492 2694
rect 27516 2692 27572 2694
rect 27596 2692 27652 2694
rect 5756 2202 5812 2204
rect 5836 2202 5892 2204
rect 5916 2202 5972 2204
rect 5996 2202 6052 2204
rect 5756 2150 5802 2202
rect 5802 2150 5812 2202
rect 5836 2150 5866 2202
rect 5866 2150 5878 2202
rect 5878 2150 5892 2202
rect 5916 2150 5930 2202
rect 5930 2150 5942 2202
rect 5942 2150 5972 2202
rect 5996 2150 6006 2202
rect 6006 2150 6052 2202
rect 5756 2148 5812 2150
rect 5836 2148 5892 2150
rect 5916 2148 5972 2150
rect 5996 2148 6052 2150
rect 10556 2202 10612 2204
rect 10636 2202 10692 2204
rect 10716 2202 10772 2204
rect 10796 2202 10852 2204
rect 10556 2150 10602 2202
rect 10602 2150 10612 2202
rect 10636 2150 10666 2202
rect 10666 2150 10678 2202
rect 10678 2150 10692 2202
rect 10716 2150 10730 2202
rect 10730 2150 10742 2202
rect 10742 2150 10772 2202
rect 10796 2150 10806 2202
rect 10806 2150 10852 2202
rect 10556 2148 10612 2150
rect 10636 2148 10692 2150
rect 10716 2148 10772 2150
rect 10796 2148 10852 2150
rect 15356 2202 15412 2204
rect 15436 2202 15492 2204
rect 15516 2202 15572 2204
rect 15596 2202 15652 2204
rect 15356 2150 15402 2202
rect 15402 2150 15412 2202
rect 15436 2150 15466 2202
rect 15466 2150 15478 2202
rect 15478 2150 15492 2202
rect 15516 2150 15530 2202
rect 15530 2150 15542 2202
rect 15542 2150 15572 2202
rect 15596 2150 15606 2202
rect 15606 2150 15652 2202
rect 15356 2148 15412 2150
rect 15436 2148 15492 2150
rect 15516 2148 15572 2150
rect 15596 2148 15652 2150
rect 20156 2202 20212 2204
rect 20236 2202 20292 2204
rect 20316 2202 20372 2204
rect 20396 2202 20452 2204
rect 20156 2150 20202 2202
rect 20202 2150 20212 2202
rect 20236 2150 20266 2202
rect 20266 2150 20278 2202
rect 20278 2150 20292 2202
rect 20316 2150 20330 2202
rect 20330 2150 20342 2202
rect 20342 2150 20372 2202
rect 20396 2150 20406 2202
rect 20406 2150 20452 2202
rect 20156 2148 20212 2150
rect 20236 2148 20292 2150
rect 20316 2148 20372 2150
rect 20396 2148 20452 2150
rect 24956 2202 25012 2204
rect 25036 2202 25092 2204
rect 25116 2202 25172 2204
rect 25196 2202 25252 2204
rect 24956 2150 25002 2202
rect 25002 2150 25012 2202
rect 25036 2150 25066 2202
rect 25066 2150 25078 2202
rect 25078 2150 25092 2202
rect 25116 2150 25130 2202
rect 25130 2150 25142 2202
rect 25142 2150 25172 2202
rect 25196 2150 25206 2202
rect 25206 2150 25252 2202
rect 24956 2148 25012 2150
rect 25036 2148 25092 2150
rect 25116 2148 25172 2150
rect 25196 2148 25252 2150
rect 28354 1400 28410 1456
<< metal3 >>
rect 28349 28386 28415 28389
rect 29200 28386 30000 28416
rect 28349 28384 30000 28386
rect 28349 28328 28354 28384
rect 28410 28328 30000 28384
rect 28349 28326 30000 28328
rect 28349 28323 28415 28326
rect 29200 28296 30000 28326
rect 3346 27776 3662 27777
rect 3346 27712 3352 27776
rect 3416 27712 3432 27776
rect 3496 27712 3512 27776
rect 3576 27712 3592 27776
rect 3656 27712 3662 27776
rect 3346 27711 3662 27712
rect 8146 27776 8462 27777
rect 8146 27712 8152 27776
rect 8216 27712 8232 27776
rect 8296 27712 8312 27776
rect 8376 27712 8392 27776
rect 8456 27712 8462 27776
rect 8146 27711 8462 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 17746 27776 18062 27777
rect 17746 27712 17752 27776
rect 17816 27712 17832 27776
rect 17896 27712 17912 27776
rect 17976 27712 17992 27776
rect 18056 27712 18062 27776
rect 17746 27711 18062 27712
rect 22546 27776 22862 27777
rect 22546 27712 22552 27776
rect 22616 27712 22632 27776
rect 22696 27712 22712 27776
rect 22776 27712 22792 27776
rect 22856 27712 22862 27776
rect 22546 27711 22862 27712
rect 27346 27776 27662 27777
rect 27346 27712 27352 27776
rect 27416 27712 27432 27776
rect 27496 27712 27512 27776
rect 27576 27712 27592 27776
rect 27656 27712 27662 27776
rect 27346 27711 27662 27712
rect 5746 27232 6062 27233
rect 0 27162 800 27192
rect 5746 27168 5752 27232
rect 5816 27168 5832 27232
rect 5896 27168 5912 27232
rect 5976 27168 5992 27232
rect 6056 27168 6062 27232
rect 5746 27167 6062 27168
rect 10546 27232 10862 27233
rect 10546 27168 10552 27232
rect 10616 27168 10632 27232
rect 10696 27168 10712 27232
rect 10776 27168 10792 27232
rect 10856 27168 10862 27232
rect 10546 27167 10862 27168
rect 15346 27232 15662 27233
rect 15346 27168 15352 27232
rect 15416 27168 15432 27232
rect 15496 27168 15512 27232
rect 15576 27168 15592 27232
rect 15656 27168 15662 27232
rect 15346 27167 15662 27168
rect 20146 27232 20462 27233
rect 20146 27168 20152 27232
rect 20216 27168 20232 27232
rect 20296 27168 20312 27232
rect 20376 27168 20392 27232
rect 20456 27168 20462 27232
rect 20146 27167 20462 27168
rect 24946 27232 25262 27233
rect 24946 27168 24952 27232
rect 25016 27168 25032 27232
rect 25096 27168 25112 27232
rect 25176 27168 25192 27232
rect 25256 27168 25262 27232
rect 24946 27167 25262 27168
rect 1577 27162 1643 27165
rect 0 27160 1643 27162
rect 0 27104 1582 27160
rect 1638 27104 1643 27160
rect 0 27102 1643 27104
rect 0 27072 800 27102
rect 1577 27099 1643 27102
rect 3346 26688 3662 26689
rect 3346 26624 3352 26688
rect 3416 26624 3432 26688
rect 3496 26624 3512 26688
rect 3576 26624 3592 26688
rect 3656 26624 3662 26688
rect 3346 26623 3662 26624
rect 8146 26688 8462 26689
rect 8146 26624 8152 26688
rect 8216 26624 8232 26688
rect 8296 26624 8312 26688
rect 8376 26624 8392 26688
rect 8456 26624 8462 26688
rect 8146 26623 8462 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 17746 26688 18062 26689
rect 17746 26624 17752 26688
rect 17816 26624 17832 26688
rect 17896 26624 17912 26688
rect 17976 26624 17992 26688
rect 18056 26624 18062 26688
rect 17746 26623 18062 26624
rect 22546 26688 22862 26689
rect 22546 26624 22552 26688
rect 22616 26624 22632 26688
rect 22696 26624 22712 26688
rect 22776 26624 22792 26688
rect 22856 26624 22862 26688
rect 22546 26623 22862 26624
rect 27346 26688 27662 26689
rect 27346 26624 27352 26688
rect 27416 26624 27432 26688
rect 27496 26624 27512 26688
rect 27576 26624 27592 26688
rect 27656 26624 27662 26688
rect 27346 26623 27662 26624
rect 5746 26144 6062 26145
rect 5746 26080 5752 26144
rect 5816 26080 5832 26144
rect 5896 26080 5912 26144
rect 5976 26080 5992 26144
rect 6056 26080 6062 26144
rect 5746 26079 6062 26080
rect 10546 26144 10862 26145
rect 10546 26080 10552 26144
rect 10616 26080 10632 26144
rect 10696 26080 10712 26144
rect 10776 26080 10792 26144
rect 10856 26080 10862 26144
rect 10546 26079 10862 26080
rect 15346 26144 15662 26145
rect 15346 26080 15352 26144
rect 15416 26080 15432 26144
rect 15496 26080 15512 26144
rect 15576 26080 15592 26144
rect 15656 26080 15662 26144
rect 15346 26079 15662 26080
rect 20146 26144 20462 26145
rect 20146 26080 20152 26144
rect 20216 26080 20232 26144
rect 20296 26080 20312 26144
rect 20376 26080 20392 26144
rect 20456 26080 20462 26144
rect 20146 26079 20462 26080
rect 24946 26144 25262 26145
rect 24946 26080 24952 26144
rect 25016 26080 25032 26144
rect 25096 26080 25112 26144
rect 25176 26080 25192 26144
rect 25256 26080 25262 26144
rect 24946 26079 25262 26080
rect 28349 25938 28415 25941
rect 29200 25938 30000 25968
rect 28349 25936 30000 25938
rect 28349 25880 28354 25936
rect 28410 25880 30000 25936
rect 28349 25878 30000 25880
rect 28349 25875 28415 25878
rect 29200 25848 30000 25878
rect 3346 25600 3662 25601
rect 3346 25536 3352 25600
rect 3416 25536 3432 25600
rect 3496 25536 3512 25600
rect 3576 25536 3592 25600
rect 3656 25536 3662 25600
rect 3346 25535 3662 25536
rect 8146 25600 8462 25601
rect 8146 25536 8152 25600
rect 8216 25536 8232 25600
rect 8296 25536 8312 25600
rect 8376 25536 8392 25600
rect 8456 25536 8462 25600
rect 8146 25535 8462 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 17746 25600 18062 25601
rect 17746 25536 17752 25600
rect 17816 25536 17832 25600
rect 17896 25536 17912 25600
rect 17976 25536 17992 25600
rect 18056 25536 18062 25600
rect 17746 25535 18062 25536
rect 22546 25600 22862 25601
rect 22546 25536 22552 25600
rect 22616 25536 22632 25600
rect 22696 25536 22712 25600
rect 22776 25536 22792 25600
rect 22856 25536 22862 25600
rect 22546 25535 22862 25536
rect 27346 25600 27662 25601
rect 27346 25536 27352 25600
rect 27416 25536 27432 25600
rect 27496 25536 27512 25600
rect 27576 25536 27592 25600
rect 27656 25536 27662 25600
rect 27346 25535 27662 25536
rect 5746 25056 6062 25057
rect 5746 24992 5752 25056
rect 5816 24992 5832 25056
rect 5896 24992 5912 25056
rect 5976 24992 5992 25056
rect 6056 24992 6062 25056
rect 5746 24991 6062 24992
rect 10546 25056 10862 25057
rect 10546 24992 10552 25056
rect 10616 24992 10632 25056
rect 10696 24992 10712 25056
rect 10776 24992 10792 25056
rect 10856 24992 10862 25056
rect 10546 24991 10862 24992
rect 15346 25056 15662 25057
rect 15346 24992 15352 25056
rect 15416 24992 15432 25056
rect 15496 24992 15512 25056
rect 15576 24992 15592 25056
rect 15656 24992 15662 25056
rect 15346 24991 15662 24992
rect 20146 25056 20462 25057
rect 20146 24992 20152 25056
rect 20216 24992 20232 25056
rect 20296 24992 20312 25056
rect 20376 24992 20392 25056
rect 20456 24992 20462 25056
rect 20146 24991 20462 24992
rect 24946 25056 25262 25057
rect 24946 24992 24952 25056
rect 25016 24992 25032 25056
rect 25096 24992 25112 25056
rect 25176 24992 25192 25056
rect 25256 24992 25262 25056
rect 24946 24991 25262 24992
rect 3346 24512 3662 24513
rect 3346 24448 3352 24512
rect 3416 24448 3432 24512
rect 3496 24448 3512 24512
rect 3576 24448 3592 24512
rect 3656 24448 3662 24512
rect 3346 24447 3662 24448
rect 8146 24512 8462 24513
rect 8146 24448 8152 24512
rect 8216 24448 8232 24512
rect 8296 24448 8312 24512
rect 8376 24448 8392 24512
rect 8456 24448 8462 24512
rect 8146 24447 8462 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 17746 24512 18062 24513
rect 17746 24448 17752 24512
rect 17816 24448 17832 24512
rect 17896 24448 17912 24512
rect 17976 24448 17992 24512
rect 18056 24448 18062 24512
rect 17746 24447 18062 24448
rect 22546 24512 22862 24513
rect 22546 24448 22552 24512
rect 22616 24448 22632 24512
rect 22696 24448 22712 24512
rect 22776 24448 22792 24512
rect 22856 24448 22862 24512
rect 22546 24447 22862 24448
rect 27346 24512 27662 24513
rect 27346 24448 27352 24512
rect 27416 24448 27432 24512
rect 27496 24448 27512 24512
rect 27576 24448 27592 24512
rect 27656 24448 27662 24512
rect 27346 24447 27662 24448
rect 5746 23968 6062 23969
rect 5746 23904 5752 23968
rect 5816 23904 5832 23968
rect 5896 23904 5912 23968
rect 5976 23904 5992 23968
rect 6056 23904 6062 23968
rect 5746 23903 6062 23904
rect 10546 23968 10862 23969
rect 10546 23904 10552 23968
rect 10616 23904 10632 23968
rect 10696 23904 10712 23968
rect 10776 23904 10792 23968
rect 10856 23904 10862 23968
rect 10546 23903 10862 23904
rect 15346 23968 15662 23969
rect 15346 23904 15352 23968
rect 15416 23904 15432 23968
rect 15496 23904 15512 23968
rect 15576 23904 15592 23968
rect 15656 23904 15662 23968
rect 15346 23903 15662 23904
rect 20146 23968 20462 23969
rect 20146 23904 20152 23968
rect 20216 23904 20232 23968
rect 20296 23904 20312 23968
rect 20376 23904 20392 23968
rect 20456 23904 20462 23968
rect 20146 23903 20462 23904
rect 24946 23968 25262 23969
rect 24946 23904 24952 23968
rect 25016 23904 25032 23968
rect 25096 23904 25112 23968
rect 25176 23904 25192 23968
rect 25256 23904 25262 23968
rect 24946 23903 25262 23904
rect 28349 23490 28415 23493
rect 29200 23490 30000 23520
rect 28349 23488 30000 23490
rect 28349 23432 28354 23488
rect 28410 23432 30000 23488
rect 28349 23430 30000 23432
rect 28349 23427 28415 23430
rect 3346 23424 3662 23425
rect 3346 23360 3352 23424
rect 3416 23360 3432 23424
rect 3496 23360 3512 23424
rect 3576 23360 3592 23424
rect 3656 23360 3662 23424
rect 3346 23359 3662 23360
rect 8146 23424 8462 23425
rect 8146 23360 8152 23424
rect 8216 23360 8232 23424
rect 8296 23360 8312 23424
rect 8376 23360 8392 23424
rect 8456 23360 8462 23424
rect 8146 23359 8462 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 17746 23424 18062 23425
rect 17746 23360 17752 23424
rect 17816 23360 17832 23424
rect 17896 23360 17912 23424
rect 17976 23360 17992 23424
rect 18056 23360 18062 23424
rect 17746 23359 18062 23360
rect 22546 23424 22862 23425
rect 22546 23360 22552 23424
rect 22616 23360 22632 23424
rect 22696 23360 22712 23424
rect 22776 23360 22792 23424
rect 22856 23360 22862 23424
rect 22546 23359 22862 23360
rect 27346 23424 27662 23425
rect 27346 23360 27352 23424
rect 27416 23360 27432 23424
rect 27496 23360 27512 23424
rect 27576 23360 27592 23424
rect 27656 23360 27662 23424
rect 29200 23400 30000 23430
rect 27346 23359 27662 23360
rect 5746 22880 6062 22881
rect 5746 22816 5752 22880
rect 5816 22816 5832 22880
rect 5896 22816 5912 22880
rect 5976 22816 5992 22880
rect 6056 22816 6062 22880
rect 5746 22815 6062 22816
rect 10546 22880 10862 22881
rect 10546 22816 10552 22880
rect 10616 22816 10632 22880
rect 10696 22816 10712 22880
rect 10776 22816 10792 22880
rect 10856 22816 10862 22880
rect 10546 22815 10862 22816
rect 15346 22880 15662 22881
rect 15346 22816 15352 22880
rect 15416 22816 15432 22880
rect 15496 22816 15512 22880
rect 15576 22816 15592 22880
rect 15656 22816 15662 22880
rect 15346 22815 15662 22816
rect 20146 22880 20462 22881
rect 20146 22816 20152 22880
rect 20216 22816 20232 22880
rect 20296 22816 20312 22880
rect 20376 22816 20392 22880
rect 20456 22816 20462 22880
rect 20146 22815 20462 22816
rect 24946 22880 25262 22881
rect 24946 22816 24952 22880
rect 25016 22816 25032 22880
rect 25096 22816 25112 22880
rect 25176 22816 25192 22880
rect 25256 22816 25262 22880
rect 24946 22815 25262 22816
rect 3346 22336 3662 22337
rect 0 22266 800 22296
rect 3346 22272 3352 22336
rect 3416 22272 3432 22336
rect 3496 22272 3512 22336
rect 3576 22272 3592 22336
rect 3656 22272 3662 22336
rect 3346 22271 3662 22272
rect 8146 22336 8462 22337
rect 8146 22272 8152 22336
rect 8216 22272 8232 22336
rect 8296 22272 8312 22336
rect 8376 22272 8392 22336
rect 8456 22272 8462 22336
rect 8146 22271 8462 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 17746 22336 18062 22337
rect 17746 22272 17752 22336
rect 17816 22272 17832 22336
rect 17896 22272 17912 22336
rect 17976 22272 17992 22336
rect 18056 22272 18062 22336
rect 17746 22271 18062 22272
rect 22546 22336 22862 22337
rect 22546 22272 22552 22336
rect 22616 22272 22632 22336
rect 22696 22272 22712 22336
rect 22776 22272 22792 22336
rect 22856 22272 22862 22336
rect 22546 22271 22862 22272
rect 27346 22336 27662 22337
rect 27346 22272 27352 22336
rect 27416 22272 27432 22336
rect 27496 22272 27512 22336
rect 27576 22272 27592 22336
rect 27656 22272 27662 22336
rect 27346 22271 27662 22272
rect 1577 22266 1643 22269
rect 0 22264 1643 22266
rect 0 22208 1582 22264
rect 1638 22208 1643 22264
rect 0 22206 1643 22208
rect 0 22176 800 22206
rect 1577 22203 1643 22206
rect 5746 21792 6062 21793
rect 5746 21728 5752 21792
rect 5816 21728 5832 21792
rect 5896 21728 5912 21792
rect 5976 21728 5992 21792
rect 6056 21728 6062 21792
rect 5746 21727 6062 21728
rect 10546 21792 10862 21793
rect 10546 21728 10552 21792
rect 10616 21728 10632 21792
rect 10696 21728 10712 21792
rect 10776 21728 10792 21792
rect 10856 21728 10862 21792
rect 10546 21727 10862 21728
rect 15346 21792 15662 21793
rect 15346 21728 15352 21792
rect 15416 21728 15432 21792
rect 15496 21728 15512 21792
rect 15576 21728 15592 21792
rect 15656 21728 15662 21792
rect 15346 21727 15662 21728
rect 20146 21792 20462 21793
rect 20146 21728 20152 21792
rect 20216 21728 20232 21792
rect 20296 21728 20312 21792
rect 20376 21728 20392 21792
rect 20456 21728 20462 21792
rect 20146 21727 20462 21728
rect 24946 21792 25262 21793
rect 24946 21728 24952 21792
rect 25016 21728 25032 21792
rect 25096 21728 25112 21792
rect 25176 21728 25192 21792
rect 25256 21728 25262 21792
rect 24946 21727 25262 21728
rect 3346 21248 3662 21249
rect 3346 21184 3352 21248
rect 3416 21184 3432 21248
rect 3496 21184 3512 21248
rect 3576 21184 3592 21248
rect 3656 21184 3662 21248
rect 3346 21183 3662 21184
rect 8146 21248 8462 21249
rect 8146 21184 8152 21248
rect 8216 21184 8232 21248
rect 8296 21184 8312 21248
rect 8376 21184 8392 21248
rect 8456 21184 8462 21248
rect 8146 21183 8462 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 17746 21248 18062 21249
rect 17746 21184 17752 21248
rect 17816 21184 17832 21248
rect 17896 21184 17912 21248
rect 17976 21184 17992 21248
rect 18056 21184 18062 21248
rect 17746 21183 18062 21184
rect 22546 21248 22862 21249
rect 22546 21184 22552 21248
rect 22616 21184 22632 21248
rect 22696 21184 22712 21248
rect 22776 21184 22792 21248
rect 22856 21184 22862 21248
rect 22546 21183 22862 21184
rect 27346 21248 27662 21249
rect 27346 21184 27352 21248
rect 27416 21184 27432 21248
rect 27496 21184 27512 21248
rect 27576 21184 27592 21248
rect 27656 21184 27662 21248
rect 27346 21183 27662 21184
rect 28349 21042 28415 21045
rect 29200 21042 30000 21072
rect 28349 21040 30000 21042
rect 28349 20984 28354 21040
rect 28410 20984 30000 21040
rect 28349 20982 30000 20984
rect 28349 20979 28415 20982
rect 29200 20952 30000 20982
rect 5746 20704 6062 20705
rect 5746 20640 5752 20704
rect 5816 20640 5832 20704
rect 5896 20640 5912 20704
rect 5976 20640 5992 20704
rect 6056 20640 6062 20704
rect 5746 20639 6062 20640
rect 10546 20704 10862 20705
rect 10546 20640 10552 20704
rect 10616 20640 10632 20704
rect 10696 20640 10712 20704
rect 10776 20640 10792 20704
rect 10856 20640 10862 20704
rect 10546 20639 10862 20640
rect 15346 20704 15662 20705
rect 15346 20640 15352 20704
rect 15416 20640 15432 20704
rect 15496 20640 15512 20704
rect 15576 20640 15592 20704
rect 15656 20640 15662 20704
rect 15346 20639 15662 20640
rect 20146 20704 20462 20705
rect 20146 20640 20152 20704
rect 20216 20640 20232 20704
rect 20296 20640 20312 20704
rect 20376 20640 20392 20704
rect 20456 20640 20462 20704
rect 20146 20639 20462 20640
rect 24946 20704 25262 20705
rect 24946 20640 24952 20704
rect 25016 20640 25032 20704
rect 25096 20640 25112 20704
rect 25176 20640 25192 20704
rect 25256 20640 25262 20704
rect 24946 20639 25262 20640
rect 3346 20160 3662 20161
rect 3346 20096 3352 20160
rect 3416 20096 3432 20160
rect 3496 20096 3512 20160
rect 3576 20096 3592 20160
rect 3656 20096 3662 20160
rect 3346 20095 3662 20096
rect 8146 20160 8462 20161
rect 8146 20096 8152 20160
rect 8216 20096 8232 20160
rect 8296 20096 8312 20160
rect 8376 20096 8392 20160
rect 8456 20096 8462 20160
rect 8146 20095 8462 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 17746 20160 18062 20161
rect 17746 20096 17752 20160
rect 17816 20096 17832 20160
rect 17896 20096 17912 20160
rect 17976 20096 17992 20160
rect 18056 20096 18062 20160
rect 17746 20095 18062 20096
rect 22546 20160 22862 20161
rect 22546 20096 22552 20160
rect 22616 20096 22632 20160
rect 22696 20096 22712 20160
rect 22776 20096 22792 20160
rect 22856 20096 22862 20160
rect 22546 20095 22862 20096
rect 27346 20160 27662 20161
rect 27346 20096 27352 20160
rect 27416 20096 27432 20160
rect 27496 20096 27512 20160
rect 27576 20096 27592 20160
rect 27656 20096 27662 20160
rect 27346 20095 27662 20096
rect 5746 19616 6062 19617
rect 5746 19552 5752 19616
rect 5816 19552 5832 19616
rect 5896 19552 5912 19616
rect 5976 19552 5992 19616
rect 6056 19552 6062 19616
rect 5746 19551 6062 19552
rect 10546 19616 10862 19617
rect 10546 19552 10552 19616
rect 10616 19552 10632 19616
rect 10696 19552 10712 19616
rect 10776 19552 10792 19616
rect 10856 19552 10862 19616
rect 10546 19551 10862 19552
rect 15346 19616 15662 19617
rect 15346 19552 15352 19616
rect 15416 19552 15432 19616
rect 15496 19552 15512 19616
rect 15576 19552 15592 19616
rect 15656 19552 15662 19616
rect 15346 19551 15662 19552
rect 20146 19616 20462 19617
rect 20146 19552 20152 19616
rect 20216 19552 20232 19616
rect 20296 19552 20312 19616
rect 20376 19552 20392 19616
rect 20456 19552 20462 19616
rect 20146 19551 20462 19552
rect 24946 19616 25262 19617
rect 24946 19552 24952 19616
rect 25016 19552 25032 19616
rect 25096 19552 25112 19616
rect 25176 19552 25192 19616
rect 25256 19552 25262 19616
rect 24946 19551 25262 19552
rect 3346 19072 3662 19073
rect 3346 19008 3352 19072
rect 3416 19008 3432 19072
rect 3496 19008 3512 19072
rect 3576 19008 3592 19072
rect 3656 19008 3662 19072
rect 3346 19007 3662 19008
rect 8146 19072 8462 19073
rect 8146 19008 8152 19072
rect 8216 19008 8232 19072
rect 8296 19008 8312 19072
rect 8376 19008 8392 19072
rect 8456 19008 8462 19072
rect 8146 19007 8462 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 17746 19072 18062 19073
rect 17746 19008 17752 19072
rect 17816 19008 17832 19072
rect 17896 19008 17912 19072
rect 17976 19008 17992 19072
rect 18056 19008 18062 19072
rect 17746 19007 18062 19008
rect 22546 19072 22862 19073
rect 22546 19008 22552 19072
rect 22616 19008 22632 19072
rect 22696 19008 22712 19072
rect 22776 19008 22792 19072
rect 22856 19008 22862 19072
rect 22546 19007 22862 19008
rect 27346 19072 27662 19073
rect 27346 19008 27352 19072
rect 27416 19008 27432 19072
rect 27496 19008 27512 19072
rect 27576 19008 27592 19072
rect 27656 19008 27662 19072
rect 27346 19007 27662 19008
rect 28349 18594 28415 18597
rect 29200 18594 30000 18624
rect 28349 18592 30000 18594
rect 28349 18536 28354 18592
rect 28410 18536 30000 18592
rect 28349 18534 30000 18536
rect 28349 18531 28415 18534
rect 5746 18528 6062 18529
rect 5746 18464 5752 18528
rect 5816 18464 5832 18528
rect 5896 18464 5912 18528
rect 5976 18464 5992 18528
rect 6056 18464 6062 18528
rect 5746 18463 6062 18464
rect 10546 18528 10862 18529
rect 10546 18464 10552 18528
rect 10616 18464 10632 18528
rect 10696 18464 10712 18528
rect 10776 18464 10792 18528
rect 10856 18464 10862 18528
rect 10546 18463 10862 18464
rect 15346 18528 15662 18529
rect 15346 18464 15352 18528
rect 15416 18464 15432 18528
rect 15496 18464 15512 18528
rect 15576 18464 15592 18528
rect 15656 18464 15662 18528
rect 15346 18463 15662 18464
rect 20146 18528 20462 18529
rect 20146 18464 20152 18528
rect 20216 18464 20232 18528
rect 20296 18464 20312 18528
rect 20376 18464 20392 18528
rect 20456 18464 20462 18528
rect 20146 18463 20462 18464
rect 24946 18528 25262 18529
rect 24946 18464 24952 18528
rect 25016 18464 25032 18528
rect 25096 18464 25112 18528
rect 25176 18464 25192 18528
rect 25256 18464 25262 18528
rect 29200 18504 30000 18534
rect 24946 18463 25262 18464
rect 3346 17984 3662 17985
rect 3346 17920 3352 17984
rect 3416 17920 3432 17984
rect 3496 17920 3512 17984
rect 3576 17920 3592 17984
rect 3656 17920 3662 17984
rect 3346 17919 3662 17920
rect 8146 17984 8462 17985
rect 8146 17920 8152 17984
rect 8216 17920 8232 17984
rect 8296 17920 8312 17984
rect 8376 17920 8392 17984
rect 8456 17920 8462 17984
rect 8146 17919 8462 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 17746 17984 18062 17985
rect 17746 17920 17752 17984
rect 17816 17920 17832 17984
rect 17896 17920 17912 17984
rect 17976 17920 17992 17984
rect 18056 17920 18062 17984
rect 17746 17919 18062 17920
rect 22546 17984 22862 17985
rect 22546 17920 22552 17984
rect 22616 17920 22632 17984
rect 22696 17920 22712 17984
rect 22776 17920 22792 17984
rect 22856 17920 22862 17984
rect 22546 17919 22862 17920
rect 27346 17984 27662 17985
rect 27346 17920 27352 17984
rect 27416 17920 27432 17984
rect 27496 17920 27512 17984
rect 27576 17920 27592 17984
rect 27656 17920 27662 17984
rect 27346 17919 27662 17920
rect 5746 17440 6062 17441
rect 0 17370 800 17400
rect 5746 17376 5752 17440
rect 5816 17376 5832 17440
rect 5896 17376 5912 17440
rect 5976 17376 5992 17440
rect 6056 17376 6062 17440
rect 5746 17375 6062 17376
rect 10546 17440 10862 17441
rect 10546 17376 10552 17440
rect 10616 17376 10632 17440
rect 10696 17376 10712 17440
rect 10776 17376 10792 17440
rect 10856 17376 10862 17440
rect 10546 17375 10862 17376
rect 15346 17440 15662 17441
rect 15346 17376 15352 17440
rect 15416 17376 15432 17440
rect 15496 17376 15512 17440
rect 15576 17376 15592 17440
rect 15656 17376 15662 17440
rect 15346 17375 15662 17376
rect 20146 17440 20462 17441
rect 20146 17376 20152 17440
rect 20216 17376 20232 17440
rect 20296 17376 20312 17440
rect 20376 17376 20392 17440
rect 20456 17376 20462 17440
rect 20146 17375 20462 17376
rect 24946 17440 25262 17441
rect 24946 17376 24952 17440
rect 25016 17376 25032 17440
rect 25096 17376 25112 17440
rect 25176 17376 25192 17440
rect 25256 17376 25262 17440
rect 24946 17375 25262 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 3346 16896 3662 16897
rect 3346 16832 3352 16896
rect 3416 16832 3432 16896
rect 3496 16832 3512 16896
rect 3576 16832 3592 16896
rect 3656 16832 3662 16896
rect 3346 16831 3662 16832
rect 8146 16896 8462 16897
rect 8146 16832 8152 16896
rect 8216 16832 8232 16896
rect 8296 16832 8312 16896
rect 8376 16832 8392 16896
rect 8456 16832 8462 16896
rect 8146 16831 8462 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 17746 16896 18062 16897
rect 17746 16832 17752 16896
rect 17816 16832 17832 16896
rect 17896 16832 17912 16896
rect 17976 16832 17992 16896
rect 18056 16832 18062 16896
rect 17746 16831 18062 16832
rect 22546 16896 22862 16897
rect 22546 16832 22552 16896
rect 22616 16832 22632 16896
rect 22696 16832 22712 16896
rect 22776 16832 22792 16896
rect 22856 16832 22862 16896
rect 22546 16831 22862 16832
rect 27346 16896 27662 16897
rect 27346 16832 27352 16896
rect 27416 16832 27432 16896
rect 27496 16832 27512 16896
rect 27576 16832 27592 16896
rect 27656 16832 27662 16896
rect 27346 16831 27662 16832
rect 5746 16352 6062 16353
rect 5746 16288 5752 16352
rect 5816 16288 5832 16352
rect 5896 16288 5912 16352
rect 5976 16288 5992 16352
rect 6056 16288 6062 16352
rect 5746 16287 6062 16288
rect 10546 16352 10862 16353
rect 10546 16288 10552 16352
rect 10616 16288 10632 16352
rect 10696 16288 10712 16352
rect 10776 16288 10792 16352
rect 10856 16288 10862 16352
rect 10546 16287 10862 16288
rect 15346 16352 15662 16353
rect 15346 16288 15352 16352
rect 15416 16288 15432 16352
rect 15496 16288 15512 16352
rect 15576 16288 15592 16352
rect 15656 16288 15662 16352
rect 15346 16287 15662 16288
rect 20146 16352 20462 16353
rect 20146 16288 20152 16352
rect 20216 16288 20232 16352
rect 20296 16288 20312 16352
rect 20376 16288 20392 16352
rect 20456 16288 20462 16352
rect 20146 16287 20462 16288
rect 24946 16352 25262 16353
rect 24946 16288 24952 16352
rect 25016 16288 25032 16352
rect 25096 16288 25112 16352
rect 25176 16288 25192 16352
rect 25256 16288 25262 16352
rect 24946 16287 25262 16288
rect 28349 16146 28415 16149
rect 29200 16146 30000 16176
rect 28349 16144 30000 16146
rect 28349 16088 28354 16144
rect 28410 16088 30000 16144
rect 28349 16086 30000 16088
rect 28349 16083 28415 16086
rect 29200 16056 30000 16086
rect 3346 15808 3662 15809
rect 3346 15744 3352 15808
rect 3416 15744 3432 15808
rect 3496 15744 3512 15808
rect 3576 15744 3592 15808
rect 3656 15744 3662 15808
rect 3346 15743 3662 15744
rect 8146 15808 8462 15809
rect 8146 15744 8152 15808
rect 8216 15744 8232 15808
rect 8296 15744 8312 15808
rect 8376 15744 8392 15808
rect 8456 15744 8462 15808
rect 8146 15743 8462 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 17746 15808 18062 15809
rect 17746 15744 17752 15808
rect 17816 15744 17832 15808
rect 17896 15744 17912 15808
rect 17976 15744 17992 15808
rect 18056 15744 18062 15808
rect 17746 15743 18062 15744
rect 22546 15808 22862 15809
rect 22546 15744 22552 15808
rect 22616 15744 22632 15808
rect 22696 15744 22712 15808
rect 22776 15744 22792 15808
rect 22856 15744 22862 15808
rect 22546 15743 22862 15744
rect 27346 15808 27662 15809
rect 27346 15744 27352 15808
rect 27416 15744 27432 15808
rect 27496 15744 27512 15808
rect 27576 15744 27592 15808
rect 27656 15744 27662 15808
rect 27346 15743 27662 15744
rect 5746 15264 6062 15265
rect 5746 15200 5752 15264
rect 5816 15200 5832 15264
rect 5896 15200 5912 15264
rect 5976 15200 5992 15264
rect 6056 15200 6062 15264
rect 5746 15199 6062 15200
rect 10546 15264 10862 15265
rect 10546 15200 10552 15264
rect 10616 15200 10632 15264
rect 10696 15200 10712 15264
rect 10776 15200 10792 15264
rect 10856 15200 10862 15264
rect 10546 15199 10862 15200
rect 15346 15264 15662 15265
rect 15346 15200 15352 15264
rect 15416 15200 15432 15264
rect 15496 15200 15512 15264
rect 15576 15200 15592 15264
rect 15656 15200 15662 15264
rect 15346 15199 15662 15200
rect 20146 15264 20462 15265
rect 20146 15200 20152 15264
rect 20216 15200 20232 15264
rect 20296 15200 20312 15264
rect 20376 15200 20392 15264
rect 20456 15200 20462 15264
rect 20146 15199 20462 15200
rect 24946 15264 25262 15265
rect 24946 15200 24952 15264
rect 25016 15200 25032 15264
rect 25096 15200 25112 15264
rect 25176 15200 25192 15264
rect 25256 15200 25262 15264
rect 24946 15199 25262 15200
rect 3346 14720 3662 14721
rect 3346 14656 3352 14720
rect 3416 14656 3432 14720
rect 3496 14656 3512 14720
rect 3576 14656 3592 14720
rect 3656 14656 3662 14720
rect 3346 14655 3662 14656
rect 8146 14720 8462 14721
rect 8146 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8312 14720
rect 8376 14656 8392 14720
rect 8456 14656 8462 14720
rect 8146 14655 8462 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 17746 14720 18062 14721
rect 17746 14656 17752 14720
rect 17816 14656 17832 14720
rect 17896 14656 17912 14720
rect 17976 14656 17992 14720
rect 18056 14656 18062 14720
rect 17746 14655 18062 14656
rect 22546 14720 22862 14721
rect 22546 14656 22552 14720
rect 22616 14656 22632 14720
rect 22696 14656 22712 14720
rect 22776 14656 22792 14720
rect 22856 14656 22862 14720
rect 22546 14655 22862 14656
rect 27346 14720 27662 14721
rect 27346 14656 27352 14720
rect 27416 14656 27432 14720
rect 27496 14656 27512 14720
rect 27576 14656 27592 14720
rect 27656 14656 27662 14720
rect 27346 14655 27662 14656
rect 5746 14176 6062 14177
rect 5746 14112 5752 14176
rect 5816 14112 5832 14176
rect 5896 14112 5912 14176
rect 5976 14112 5992 14176
rect 6056 14112 6062 14176
rect 5746 14111 6062 14112
rect 10546 14176 10862 14177
rect 10546 14112 10552 14176
rect 10616 14112 10632 14176
rect 10696 14112 10712 14176
rect 10776 14112 10792 14176
rect 10856 14112 10862 14176
rect 10546 14111 10862 14112
rect 15346 14176 15662 14177
rect 15346 14112 15352 14176
rect 15416 14112 15432 14176
rect 15496 14112 15512 14176
rect 15576 14112 15592 14176
rect 15656 14112 15662 14176
rect 15346 14111 15662 14112
rect 20146 14176 20462 14177
rect 20146 14112 20152 14176
rect 20216 14112 20232 14176
rect 20296 14112 20312 14176
rect 20376 14112 20392 14176
rect 20456 14112 20462 14176
rect 20146 14111 20462 14112
rect 24946 14176 25262 14177
rect 24946 14112 24952 14176
rect 25016 14112 25032 14176
rect 25096 14112 25112 14176
rect 25176 14112 25192 14176
rect 25256 14112 25262 14176
rect 24946 14111 25262 14112
rect 28349 13698 28415 13701
rect 29200 13698 30000 13728
rect 28349 13696 30000 13698
rect 28349 13640 28354 13696
rect 28410 13640 30000 13696
rect 28349 13638 30000 13640
rect 28349 13635 28415 13638
rect 3346 13632 3662 13633
rect 3346 13568 3352 13632
rect 3416 13568 3432 13632
rect 3496 13568 3512 13632
rect 3576 13568 3592 13632
rect 3656 13568 3662 13632
rect 3346 13567 3662 13568
rect 8146 13632 8462 13633
rect 8146 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8312 13632
rect 8376 13568 8392 13632
rect 8456 13568 8462 13632
rect 8146 13567 8462 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 17746 13632 18062 13633
rect 17746 13568 17752 13632
rect 17816 13568 17832 13632
rect 17896 13568 17912 13632
rect 17976 13568 17992 13632
rect 18056 13568 18062 13632
rect 17746 13567 18062 13568
rect 22546 13632 22862 13633
rect 22546 13568 22552 13632
rect 22616 13568 22632 13632
rect 22696 13568 22712 13632
rect 22776 13568 22792 13632
rect 22856 13568 22862 13632
rect 22546 13567 22862 13568
rect 27346 13632 27662 13633
rect 27346 13568 27352 13632
rect 27416 13568 27432 13632
rect 27496 13568 27512 13632
rect 27576 13568 27592 13632
rect 27656 13568 27662 13632
rect 29200 13608 30000 13638
rect 27346 13567 27662 13568
rect 5746 13088 6062 13089
rect 5746 13024 5752 13088
rect 5816 13024 5832 13088
rect 5896 13024 5912 13088
rect 5976 13024 5992 13088
rect 6056 13024 6062 13088
rect 5746 13023 6062 13024
rect 10546 13088 10862 13089
rect 10546 13024 10552 13088
rect 10616 13024 10632 13088
rect 10696 13024 10712 13088
rect 10776 13024 10792 13088
rect 10856 13024 10862 13088
rect 10546 13023 10862 13024
rect 15346 13088 15662 13089
rect 15346 13024 15352 13088
rect 15416 13024 15432 13088
rect 15496 13024 15512 13088
rect 15576 13024 15592 13088
rect 15656 13024 15662 13088
rect 15346 13023 15662 13024
rect 20146 13088 20462 13089
rect 20146 13024 20152 13088
rect 20216 13024 20232 13088
rect 20296 13024 20312 13088
rect 20376 13024 20392 13088
rect 20456 13024 20462 13088
rect 20146 13023 20462 13024
rect 24946 13088 25262 13089
rect 24946 13024 24952 13088
rect 25016 13024 25032 13088
rect 25096 13024 25112 13088
rect 25176 13024 25192 13088
rect 25256 13024 25262 13088
rect 24946 13023 25262 13024
rect 3346 12544 3662 12545
rect 0 12474 800 12504
rect 3346 12480 3352 12544
rect 3416 12480 3432 12544
rect 3496 12480 3512 12544
rect 3576 12480 3592 12544
rect 3656 12480 3662 12544
rect 3346 12479 3662 12480
rect 8146 12544 8462 12545
rect 8146 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8312 12544
rect 8376 12480 8392 12544
rect 8456 12480 8462 12544
rect 8146 12479 8462 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 17746 12544 18062 12545
rect 17746 12480 17752 12544
rect 17816 12480 17832 12544
rect 17896 12480 17912 12544
rect 17976 12480 17992 12544
rect 18056 12480 18062 12544
rect 17746 12479 18062 12480
rect 22546 12544 22862 12545
rect 22546 12480 22552 12544
rect 22616 12480 22632 12544
rect 22696 12480 22712 12544
rect 22776 12480 22792 12544
rect 22856 12480 22862 12544
rect 22546 12479 22862 12480
rect 27346 12544 27662 12545
rect 27346 12480 27352 12544
rect 27416 12480 27432 12544
rect 27496 12480 27512 12544
rect 27576 12480 27592 12544
rect 27656 12480 27662 12544
rect 27346 12479 27662 12480
rect 1485 12474 1551 12477
rect 0 12472 1551 12474
rect 0 12416 1490 12472
rect 1546 12416 1551 12472
rect 0 12414 1551 12416
rect 0 12384 800 12414
rect 1485 12411 1551 12414
rect 5746 12000 6062 12001
rect 5746 11936 5752 12000
rect 5816 11936 5832 12000
rect 5896 11936 5912 12000
rect 5976 11936 5992 12000
rect 6056 11936 6062 12000
rect 5746 11935 6062 11936
rect 10546 12000 10862 12001
rect 10546 11936 10552 12000
rect 10616 11936 10632 12000
rect 10696 11936 10712 12000
rect 10776 11936 10792 12000
rect 10856 11936 10862 12000
rect 10546 11935 10862 11936
rect 15346 12000 15662 12001
rect 15346 11936 15352 12000
rect 15416 11936 15432 12000
rect 15496 11936 15512 12000
rect 15576 11936 15592 12000
rect 15656 11936 15662 12000
rect 15346 11935 15662 11936
rect 20146 12000 20462 12001
rect 20146 11936 20152 12000
rect 20216 11936 20232 12000
rect 20296 11936 20312 12000
rect 20376 11936 20392 12000
rect 20456 11936 20462 12000
rect 20146 11935 20462 11936
rect 24946 12000 25262 12001
rect 24946 11936 24952 12000
rect 25016 11936 25032 12000
rect 25096 11936 25112 12000
rect 25176 11936 25192 12000
rect 25256 11936 25262 12000
rect 24946 11935 25262 11936
rect 3346 11456 3662 11457
rect 3346 11392 3352 11456
rect 3416 11392 3432 11456
rect 3496 11392 3512 11456
rect 3576 11392 3592 11456
rect 3656 11392 3662 11456
rect 3346 11391 3662 11392
rect 8146 11456 8462 11457
rect 8146 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8312 11456
rect 8376 11392 8392 11456
rect 8456 11392 8462 11456
rect 8146 11391 8462 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 17746 11456 18062 11457
rect 17746 11392 17752 11456
rect 17816 11392 17832 11456
rect 17896 11392 17912 11456
rect 17976 11392 17992 11456
rect 18056 11392 18062 11456
rect 17746 11391 18062 11392
rect 22546 11456 22862 11457
rect 22546 11392 22552 11456
rect 22616 11392 22632 11456
rect 22696 11392 22712 11456
rect 22776 11392 22792 11456
rect 22856 11392 22862 11456
rect 22546 11391 22862 11392
rect 27346 11456 27662 11457
rect 27346 11392 27352 11456
rect 27416 11392 27432 11456
rect 27496 11392 27512 11456
rect 27576 11392 27592 11456
rect 27656 11392 27662 11456
rect 27346 11391 27662 11392
rect 28349 11250 28415 11253
rect 29200 11250 30000 11280
rect 28349 11248 30000 11250
rect 28349 11192 28354 11248
rect 28410 11192 30000 11248
rect 28349 11190 30000 11192
rect 28349 11187 28415 11190
rect 29200 11160 30000 11190
rect 5746 10912 6062 10913
rect 5746 10848 5752 10912
rect 5816 10848 5832 10912
rect 5896 10848 5912 10912
rect 5976 10848 5992 10912
rect 6056 10848 6062 10912
rect 5746 10847 6062 10848
rect 10546 10912 10862 10913
rect 10546 10848 10552 10912
rect 10616 10848 10632 10912
rect 10696 10848 10712 10912
rect 10776 10848 10792 10912
rect 10856 10848 10862 10912
rect 10546 10847 10862 10848
rect 15346 10912 15662 10913
rect 15346 10848 15352 10912
rect 15416 10848 15432 10912
rect 15496 10848 15512 10912
rect 15576 10848 15592 10912
rect 15656 10848 15662 10912
rect 15346 10847 15662 10848
rect 20146 10912 20462 10913
rect 20146 10848 20152 10912
rect 20216 10848 20232 10912
rect 20296 10848 20312 10912
rect 20376 10848 20392 10912
rect 20456 10848 20462 10912
rect 20146 10847 20462 10848
rect 24946 10912 25262 10913
rect 24946 10848 24952 10912
rect 25016 10848 25032 10912
rect 25096 10848 25112 10912
rect 25176 10848 25192 10912
rect 25256 10848 25262 10912
rect 24946 10847 25262 10848
rect 3346 10368 3662 10369
rect 3346 10304 3352 10368
rect 3416 10304 3432 10368
rect 3496 10304 3512 10368
rect 3576 10304 3592 10368
rect 3656 10304 3662 10368
rect 3346 10303 3662 10304
rect 8146 10368 8462 10369
rect 8146 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8312 10368
rect 8376 10304 8392 10368
rect 8456 10304 8462 10368
rect 8146 10303 8462 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 17746 10368 18062 10369
rect 17746 10304 17752 10368
rect 17816 10304 17832 10368
rect 17896 10304 17912 10368
rect 17976 10304 17992 10368
rect 18056 10304 18062 10368
rect 17746 10303 18062 10304
rect 22546 10368 22862 10369
rect 22546 10304 22552 10368
rect 22616 10304 22632 10368
rect 22696 10304 22712 10368
rect 22776 10304 22792 10368
rect 22856 10304 22862 10368
rect 22546 10303 22862 10304
rect 27346 10368 27662 10369
rect 27346 10304 27352 10368
rect 27416 10304 27432 10368
rect 27496 10304 27512 10368
rect 27576 10304 27592 10368
rect 27656 10304 27662 10368
rect 27346 10303 27662 10304
rect 5746 9824 6062 9825
rect 5746 9760 5752 9824
rect 5816 9760 5832 9824
rect 5896 9760 5912 9824
rect 5976 9760 5992 9824
rect 6056 9760 6062 9824
rect 5746 9759 6062 9760
rect 10546 9824 10862 9825
rect 10546 9760 10552 9824
rect 10616 9760 10632 9824
rect 10696 9760 10712 9824
rect 10776 9760 10792 9824
rect 10856 9760 10862 9824
rect 10546 9759 10862 9760
rect 15346 9824 15662 9825
rect 15346 9760 15352 9824
rect 15416 9760 15432 9824
rect 15496 9760 15512 9824
rect 15576 9760 15592 9824
rect 15656 9760 15662 9824
rect 15346 9759 15662 9760
rect 20146 9824 20462 9825
rect 20146 9760 20152 9824
rect 20216 9760 20232 9824
rect 20296 9760 20312 9824
rect 20376 9760 20392 9824
rect 20456 9760 20462 9824
rect 20146 9759 20462 9760
rect 24946 9824 25262 9825
rect 24946 9760 24952 9824
rect 25016 9760 25032 9824
rect 25096 9760 25112 9824
rect 25176 9760 25192 9824
rect 25256 9760 25262 9824
rect 24946 9759 25262 9760
rect 3346 9280 3662 9281
rect 3346 9216 3352 9280
rect 3416 9216 3432 9280
rect 3496 9216 3512 9280
rect 3576 9216 3592 9280
rect 3656 9216 3662 9280
rect 3346 9215 3662 9216
rect 8146 9280 8462 9281
rect 8146 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8312 9280
rect 8376 9216 8392 9280
rect 8456 9216 8462 9280
rect 8146 9215 8462 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 17746 9280 18062 9281
rect 17746 9216 17752 9280
rect 17816 9216 17832 9280
rect 17896 9216 17912 9280
rect 17976 9216 17992 9280
rect 18056 9216 18062 9280
rect 17746 9215 18062 9216
rect 22546 9280 22862 9281
rect 22546 9216 22552 9280
rect 22616 9216 22632 9280
rect 22696 9216 22712 9280
rect 22776 9216 22792 9280
rect 22856 9216 22862 9280
rect 22546 9215 22862 9216
rect 27346 9280 27662 9281
rect 27346 9216 27352 9280
rect 27416 9216 27432 9280
rect 27496 9216 27512 9280
rect 27576 9216 27592 9280
rect 27656 9216 27662 9280
rect 27346 9215 27662 9216
rect 28349 8802 28415 8805
rect 29200 8802 30000 8832
rect 28349 8800 30000 8802
rect 28349 8744 28354 8800
rect 28410 8744 30000 8800
rect 28349 8742 30000 8744
rect 28349 8739 28415 8742
rect 5746 8736 6062 8737
rect 5746 8672 5752 8736
rect 5816 8672 5832 8736
rect 5896 8672 5912 8736
rect 5976 8672 5992 8736
rect 6056 8672 6062 8736
rect 5746 8671 6062 8672
rect 10546 8736 10862 8737
rect 10546 8672 10552 8736
rect 10616 8672 10632 8736
rect 10696 8672 10712 8736
rect 10776 8672 10792 8736
rect 10856 8672 10862 8736
rect 10546 8671 10862 8672
rect 15346 8736 15662 8737
rect 15346 8672 15352 8736
rect 15416 8672 15432 8736
rect 15496 8672 15512 8736
rect 15576 8672 15592 8736
rect 15656 8672 15662 8736
rect 15346 8671 15662 8672
rect 20146 8736 20462 8737
rect 20146 8672 20152 8736
rect 20216 8672 20232 8736
rect 20296 8672 20312 8736
rect 20376 8672 20392 8736
rect 20456 8672 20462 8736
rect 20146 8671 20462 8672
rect 24946 8736 25262 8737
rect 24946 8672 24952 8736
rect 25016 8672 25032 8736
rect 25096 8672 25112 8736
rect 25176 8672 25192 8736
rect 25256 8672 25262 8736
rect 29200 8712 30000 8742
rect 24946 8671 25262 8672
rect 3346 8192 3662 8193
rect 3346 8128 3352 8192
rect 3416 8128 3432 8192
rect 3496 8128 3512 8192
rect 3576 8128 3592 8192
rect 3656 8128 3662 8192
rect 3346 8127 3662 8128
rect 8146 8192 8462 8193
rect 8146 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8312 8192
rect 8376 8128 8392 8192
rect 8456 8128 8462 8192
rect 8146 8127 8462 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 17746 8192 18062 8193
rect 17746 8128 17752 8192
rect 17816 8128 17832 8192
rect 17896 8128 17912 8192
rect 17976 8128 17992 8192
rect 18056 8128 18062 8192
rect 17746 8127 18062 8128
rect 22546 8192 22862 8193
rect 22546 8128 22552 8192
rect 22616 8128 22632 8192
rect 22696 8128 22712 8192
rect 22776 8128 22792 8192
rect 22856 8128 22862 8192
rect 22546 8127 22862 8128
rect 27346 8192 27662 8193
rect 27346 8128 27352 8192
rect 27416 8128 27432 8192
rect 27496 8128 27512 8192
rect 27576 8128 27592 8192
rect 27656 8128 27662 8192
rect 27346 8127 27662 8128
rect 5746 7648 6062 7649
rect 0 7578 800 7608
rect 5746 7584 5752 7648
rect 5816 7584 5832 7648
rect 5896 7584 5912 7648
rect 5976 7584 5992 7648
rect 6056 7584 6062 7648
rect 5746 7583 6062 7584
rect 10546 7648 10862 7649
rect 10546 7584 10552 7648
rect 10616 7584 10632 7648
rect 10696 7584 10712 7648
rect 10776 7584 10792 7648
rect 10856 7584 10862 7648
rect 10546 7583 10862 7584
rect 15346 7648 15662 7649
rect 15346 7584 15352 7648
rect 15416 7584 15432 7648
rect 15496 7584 15512 7648
rect 15576 7584 15592 7648
rect 15656 7584 15662 7648
rect 15346 7583 15662 7584
rect 20146 7648 20462 7649
rect 20146 7584 20152 7648
rect 20216 7584 20232 7648
rect 20296 7584 20312 7648
rect 20376 7584 20392 7648
rect 20456 7584 20462 7648
rect 20146 7583 20462 7584
rect 24946 7648 25262 7649
rect 24946 7584 24952 7648
rect 25016 7584 25032 7648
rect 25096 7584 25112 7648
rect 25176 7584 25192 7648
rect 25256 7584 25262 7648
rect 24946 7583 25262 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 3346 7104 3662 7105
rect 3346 7040 3352 7104
rect 3416 7040 3432 7104
rect 3496 7040 3512 7104
rect 3576 7040 3592 7104
rect 3656 7040 3662 7104
rect 3346 7039 3662 7040
rect 8146 7104 8462 7105
rect 8146 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8312 7104
rect 8376 7040 8392 7104
rect 8456 7040 8462 7104
rect 8146 7039 8462 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 17746 7104 18062 7105
rect 17746 7040 17752 7104
rect 17816 7040 17832 7104
rect 17896 7040 17912 7104
rect 17976 7040 17992 7104
rect 18056 7040 18062 7104
rect 17746 7039 18062 7040
rect 22546 7104 22862 7105
rect 22546 7040 22552 7104
rect 22616 7040 22632 7104
rect 22696 7040 22712 7104
rect 22776 7040 22792 7104
rect 22856 7040 22862 7104
rect 22546 7039 22862 7040
rect 27346 7104 27662 7105
rect 27346 7040 27352 7104
rect 27416 7040 27432 7104
rect 27496 7040 27512 7104
rect 27576 7040 27592 7104
rect 27656 7040 27662 7104
rect 27346 7039 27662 7040
rect 5746 6560 6062 6561
rect 5746 6496 5752 6560
rect 5816 6496 5832 6560
rect 5896 6496 5912 6560
rect 5976 6496 5992 6560
rect 6056 6496 6062 6560
rect 5746 6495 6062 6496
rect 10546 6560 10862 6561
rect 10546 6496 10552 6560
rect 10616 6496 10632 6560
rect 10696 6496 10712 6560
rect 10776 6496 10792 6560
rect 10856 6496 10862 6560
rect 10546 6495 10862 6496
rect 15346 6560 15662 6561
rect 15346 6496 15352 6560
rect 15416 6496 15432 6560
rect 15496 6496 15512 6560
rect 15576 6496 15592 6560
rect 15656 6496 15662 6560
rect 15346 6495 15662 6496
rect 20146 6560 20462 6561
rect 20146 6496 20152 6560
rect 20216 6496 20232 6560
rect 20296 6496 20312 6560
rect 20376 6496 20392 6560
rect 20456 6496 20462 6560
rect 20146 6495 20462 6496
rect 24946 6560 25262 6561
rect 24946 6496 24952 6560
rect 25016 6496 25032 6560
rect 25096 6496 25112 6560
rect 25176 6496 25192 6560
rect 25256 6496 25262 6560
rect 24946 6495 25262 6496
rect 28349 6354 28415 6357
rect 29200 6354 30000 6384
rect 28349 6352 30000 6354
rect 28349 6296 28354 6352
rect 28410 6296 30000 6352
rect 28349 6294 30000 6296
rect 28349 6291 28415 6294
rect 29200 6264 30000 6294
rect 3346 6016 3662 6017
rect 3346 5952 3352 6016
rect 3416 5952 3432 6016
rect 3496 5952 3512 6016
rect 3576 5952 3592 6016
rect 3656 5952 3662 6016
rect 3346 5951 3662 5952
rect 8146 6016 8462 6017
rect 8146 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8312 6016
rect 8376 5952 8392 6016
rect 8456 5952 8462 6016
rect 8146 5951 8462 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 17746 6016 18062 6017
rect 17746 5952 17752 6016
rect 17816 5952 17832 6016
rect 17896 5952 17912 6016
rect 17976 5952 17992 6016
rect 18056 5952 18062 6016
rect 17746 5951 18062 5952
rect 22546 6016 22862 6017
rect 22546 5952 22552 6016
rect 22616 5952 22632 6016
rect 22696 5952 22712 6016
rect 22776 5952 22792 6016
rect 22856 5952 22862 6016
rect 22546 5951 22862 5952
rect 27346 6016 27662 6017
rect 27346 5952 27352 6016
rect 27416 5952 27432 6016
rect 27496 5952 27512 6016
rect 27576 5952 27592 6016
rect 27656 5952 27662 6016
rect 27346 5951 27662 5952
rect 5746 5472 6062 5473
rect 5746 5408 5752 5472
rect 5816 5408 5832 5472
rect 5896 5408 5912 5472
rect 5976 5408 5992 5472
rect 6056 5408 6062 5472
rect 5746 5407 6062 5408
rect 10546 5472 10862 5473
rect 10546 5408 10552 5472
rect 10616 5408 10632 5472
rect 10696 5408 10712 5472
rect 10776 5408 10792 5472
rect 10856 5408 10862 5472
rect 10546 5407 10862 5408
rect 15346 5472 15662 5473
rect 15346 5408 15352 5472
rect 15416 5408 15432 5472
rect 15496 5408 15512 5472
rect 15576 5408 15592 5472
rect 15656 5408 15662 5472
rect 15346 5407 15662 5408
rect 20146 5472 20462 5473
rect 20146 5408 20152 5472
rect 20216 5408 20232 5472
rect 20296 5408 20312 5472
rect 20376 5408 20392 5472
rect 20456 5408 20462 5472
rect 20146 5407 20462 5408
rect 24946 5472 25262 5473
rect 24946 5408 24952 5472
rect 25016 5408 25032 5472
rect 25096 5408 25112 5472
rect 25176 5408 25192 5472
rect 25256 5408 25262 5472
rect 24946 5407 25262 5408
rect 3346 4928 3662 4929
rect 3346 4864 3352 4928
rect 3416 4864 3432 4928
rect 3496 4864 3512 4928
rect 3576 4864 3592 4928
rect 3656 4864 3662 4928
rect 3346 4863 3662 4864
rect 8146 4928 8462 4929
rect 8146 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8312 4928
rect 8376 4864 8392 4928
rect 8456 4864 8462 4928
rect 8146 4863 8462 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 17746 4928 18062 4929
rect 17746 4864 17752 4928
rect 17816 4864 17832 4928
rect 17896 4864 17912 4928
rect 17976 4864 17992 4928
rect 18056 4864 18062 4928
rect 17746 4863 18062 4864
rect 22546 4928 22862 4929
rect 22546 4864 22552 4928
rect 22616 4864 22632 4928
rect 22696 4864 22712 4928
rect 22776 4864 22792 4928
rect 22856 4864 22862 4928
rect 22546 4863 22862 4864
rect 27346 4928 27662 4929
rect 27346 4864 27352 4928
rect 27416 4864 27432 4928
rect 27496 4864 27512 4928
rect 27576 4864 27592 4928
rect 27656 4864 27662 4928
rect 27346 4863 27662 4864
rect 5746 4384 6062 4385
rect 5746 4320 5752 4384
rect 5816 4320 5832 4384
rect 5896 4320 5912 4384
rect 5976 4320 5992 4384
rect 6056 4320 6062 4384
rect 5746 4319 6062 4320
rect 10546 4384 10862 4385
rect 10546 4320 10552 4384
rect 10616 4320 10632 4384
rect 10696 4320 10712 4384
rect 10776 4320 10792 4384
rect 10856 4320 10862 4384
rect 10546 4319 10862 4320
rect 15346 4384 15662 4385
rect 15346 4320 15352 4384
rect 15416 4320 15432 4384
rect 15496 4320 15512 4384
rect 15576 4320 15592 4384
rect 15656 4320 15662 4384
rect 15346 4319 15662 4320
rect 20146 4384 20462 4385
rect 20146 4320 20152 4384
rect 20216 4320 20232 4384
rect 20296 4320 20312 4384
rect 20376 4320 20392 4384
rect 20456 4320 20462 4384
rect 20146 4319 20462 4320
rect 24946 4384 25262 4385
rect 24946 4320 24952 4384
rect 25016 4320 25032 4384
rect 25096 4320 25112 4384
rect 25176 4320 25192 4384
rect 25256 4320 25262 4384
rect 24946 4319 25262 4320
rect 28349 3906 28415 3909
rect 29200 3906 30000 3936
rect 28349 3904 30000 3906
rect 28349 3848 28354 3904
rect 28410 3848 30000 3904
rect 28349 3846 30000 3848
rect 28349 3843 28415 3846
rect 3346 3840 3662 3841
rect 3346 3776 3352 3840
rect 3416 3776 3432 3840
rect 3496 3776 3512 3840
rect 3576 3776 3592 3840
rect 3656 3776 3662 3840
rect 3346 3775 3662 3776
rect 8146 3840 8462 3841
rect 8146 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8312 3840
rect 8376 3776 8392 3840
rect 8456 3776 8462 3840
rect 8146 3775 8462 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 17746 3840 18062 3841
rect 17746 3776 17752 3840
rect 17816 3776 17832 3840
rect 17896 3776 17912 3840
rect 17976 3776 17992 3840
rect 18056 3776 18062 3840
rect 17746 3775 18062 3776
rect 22546 3840 22862 3841
rect 22546 3776 22552 3840
rect 22616 3776 22632 3840
rect 22696 3776 22712 3840
rect 22776 3776 22792 3840
rect 22856 3776 22862 3840
rect 22546 3775 22862 3776
rect 27346 3840 27662 3841
rect 27346 3776 27352 3840
rect 27416 3776 27432 3840
rect 27496 3776 27512 3840
rect 27576 3776 27592 3840
rect 27656 3776 27662 3840
rect 29200 3816 30000 3846
rect 27346 3775 27662 3776
rect 5746 3296 6062 3297
rect 5746 3232 5752 3296
rect 5816 3232 5832 3296
rect 5896 3232 5912 3296
rect 5976 3232 5992 3296
rect 6056 3232 6062 3296
rect 5746 3231 6062 3232
rect 10546 3296 10862 3297
rect 10546 3232 10552 3296
rect 10616 3232 10632 3296
rect 10696 3232 10712 3296
rect 10776 3232 10792 3296
rect 10856 3232 10862 3296
rect 10546 3231 10862 3232
rect 15346 3296 15662 3297
rect 15346 3232 15352 3296
rect 15416 3232 15432 3296
rect 15496 3232 15512 3296
rect 15576 3232 15592 3296
rect 15656 3232 15662 3296
rect 15346 3231 15662 3232
rect 20146 3296 20462 3297
rect 20146 3232 20152 3296
rect 20216 3232 20232 3296
rect 20296 3232 20312 3296
rect 20376 3232 20392 3296
rect 20456 3232 20462 3296
rect 20146 3231 20462 3232
rect 24946 3296 25262 3297
rect 24946 3232 24952 3296
rect 25016 3232 25032 3296
rect 25096 3232 25112 3296
rect 25176 3232 25192 3296
rect 25256 3232 25262 3296
rect 24946 3231 25262 3232
rect 3346 2752 3662 2753
rect 0 2682 800 2712
rect 3346 2688 3352 2752
rect 3416 2688 3432 2752
rect 3496 2688 3512 2752
rect 3576 2688 3592 2752
rect 3656 2688 3662 2752
rect 3346 2687 3662 2688
rect 8146 2752 8462 2753
rect 8146 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8312 2752
rect 8376 2688 8392 2752
rect 8456 2688 8462 2752
rect 8146 2687 8462 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 17746 2752 18062 2753
rect 17746 2688 17752 2752
rect 17816 2688 17832 2752
rect 17896 2688 17912 2752
rect 17976 2688 17992 2752
rect 18056 2688 18062 2752
rect 17746 2687 18062 2688
rect 22546 2752 22862 2753
rect 22546 2688 22552 2752
rect 22616 2688 22632 2752
rect 22696 2688 22712 2752
rect 22776 2688 22792 2752
rect 22856 2688 22862 2752
rect 22546 2687 22862 2688
rect 27346 2752 27662 2753
rect 27346 2688 27352 2752
rect 27416 2688 27432 2752
rect 27496 2688 27512 2752
rect 27576 2688 27592 2752
rect 27656 2688 27662 2752
rect 27346 2687 27662 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 0 2592 800 2622
rect 1577 2619 1643 2622
rect 5746 2208 6062 2209
rect 5746 2144 5752 2208
rect 5816 2144 5832 2208
rect 5896 2144 5912 2208
rect 5976 2144 5992 2208
rect 6056 2144 6062 2208
rect 5746 2143 6062 2144
rect 10546 2208 10862 2209
rect 10546 2144 10552 2208
rect 10616 2144 10632 2208
rect 10696 2144 10712 2208
rect 10776 2144 10792 2208
rect 10856 2144 10862 2208
rect 10546 2143 10862 2144
rect 15346 2208 15662 2209
rect 15346 2144 15352 2208
rect 15416 2144 15432 2208
rect 15496 2144 15512 2208
rect 15576 2144 15592 2208
rect 15656 2144 15662 2208
rect 15346 2143 15662 2144
rect 20146 2208 20462 2209
rect 20146 2144 20152 2208
rect 20216 2144 20232 2208
rect 20296 2144 20312 2208
rect 20376 2144 20392 2208
rect 20456 2144 20462 2208
rect 20146 2143 20462 2144
rect 24946 2208 25262 2209
rect 24946 2144 24952 2208
rect 25016 2144 25032 2208
rect 25096 2144 25112 2208
rect 25176 2144 25192 2208
rect 25256 2144 25262 2208
rect 24946 2143 25262 2144
rect 28349 1458 28415 1461
rect 29200 1458 30000 1488
rect 28349 1456 30000 1458
rect 28349 1400 28354 1456
rect 28410 1400 30000 1456
rect 28349 1398 30000 1400
rect 28349 1395 28415 1398
rect 29200 1368 30000 1398
<< via3 >>
rect 3352 27772 3416 27776
rect 3352 27716 3356 27772
rect 3356 27716 3412 27772
rect 3412 27716 3416 27772
rect 3352 27712 3416 27716
rect 3432 27772 3496 27776
rect 3432 27716 3436 27772
rect 3436 27716 3492 27772
rect 3492 27716 3496 27772
rect 3432 27712 3496 27716
rect 3512 27772 3576 27776
rect 3512 27716 3516 27772
rect 3516 27716 3572 27772
rect 3572 27716 3576 27772
rect 3512 27712 3576 27716
rect 3592 27772 3656 27776
rect 3592 27716 3596 27772
rect 3596 27716 3652 27772
rect 3652 27716 3656 27772
rect 3592 27712 3656 27716
rect 8152 27772 8216 27776
rect 8152 27716 8156 27772
rect 8156 27716 8212 27772
rect 8212 27716 8216 27772
rect 8152 27712 8216 27716
rect 8232 27772 8296 27776
rect 8232 27716 8236 27772
rect 8236 27716 8292 27772
rect 8292 27716 8296 27772
rect 8232 27712 8296 27716
rect 8312 27772 8376 27776
rect 8312 27716 8316 27772
rect 8316 27716 8372 27772
rect 8372 27716 8376 27772
rect 8312 27712 8376 27716
rect 8392 27772 8456 27776
rect 8392 27716 8396 27772
rect 8396 27716 8452 27772
rect 8452 27716 8456 27772
rect 8392 27712 8456 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 17752 27772 17816 27776
rect 17752 27716 17756 27772
rect 17756 27716 17812 27772
rect 17812 27716 17816 27772
rect 17752 27712 17816 27716
rect 17832 27772 17896 27776
rect 17832 27716 17836 27772
rect 17836 27716 17892 27772
rect 17892 27716 17896 27772
rect 17832 27712 17896 27716
rect 17912 27772 17976 27776
rect 17912 27716 17916 27772
rect 17916 27716 17972 27772
rect 17972 27716 17976 27772
rect 17912 27712 17976 27716
rect 17992 27772 18056 27776
rect 17992 27716 17996 27772
rect 17996 27716 18052 27772
rect 18052 27716 18056 27772
rect 17992 27712 18056 27716
rect 22552 27772 22616 27776
rect 22552 27716 22556 27772
rect 22556 27716 22612 27772
rect 22612 27716 22616 27772
rect 22552 27712 22616 27716
rect 22632 27772 22696 27776
rect 22632 27716 22636 27772
rect 22636 27716 22692 27772
rect 22692 27716 22696 27772
rect 22632 27712 22696 27716
rect 22712 27772 22776 27776
rect 22712 27716 22716 27772
rect 22716 27716 22772 27772
rect 22772 27716 22776 27772
rect 22712 27712 22776 27716
rect 22792 27772 22856 27776
rect 22792 27716 22796 27772
rect 22796 27716 22852 27772
rect 22852 27716 22856 27772
rect 22792 27712 22856 27716
rect 27352 27772 27416 27776
rect 27352 27716 27356 27772
rect 27356 27716 27412 27772
rect 27412 27716 27416 27772
rect 27352 27712 27416 27716
rect 27432 27772 27496 27776
rect 27432 27716 27436 27772
rect 27436 27716 27492 27772
rect 27492 27716 27496 27772
rect 27432 27712 27496 27716
rect 27512 27772 27576 27776
rect 27512 27716 27516 27772
rect 27516 27716 27572 27772
rect 27572 27716 27576 27772
rect 27512 27712 27576 27716
rect 27592 27772 27656 27776
rect 27592 27716 27596 27772
rect 27596 27716 27652 27772
rect 27652 27716 27656 27772
rect 27592 27712 27656 27716
rect 5752 27228 5816 27232
rect 5752 27172 5756 27228
rect 5756 27172 5812 27228
rect 5812 27172 5816 27228
rect 5752 27168 5816 27172
rect 5832 27228 5896 27232
rect 5832 27172 5836 27228
rect 5836 27172 5892 27228
rect 5892 27172 5896 27228
rect 5832 27168 5896 27172
rect 5912 27228 5976 27232
rect 5912 27172 5916 27228
rect 5916 27172 5972 27228
rect 5972 27172 5976 27228
rect 5912 27168 5976 27172
rect 5992 27228 6056 27232
rect 5992 27172 5996 27228
rect 5996 27172 6052 27228
rect 6052 27172 6056 27228
rect 5992 27168 6056 27172
rect 10552 27228 10616 27232
rect 10552 27172 10556 27228
rect 10556 27172 10612 27228
rect 10612 27172 10616 27228
rect 10552 27168 10616 27172
rect 10632 27228 10696 27232
rect 10632 27172 10636 27228
rect 10636 27172 10692 27228
rect 10692 27172 10696 27228
rect 10632 27168 10696 27172
rect 10712 27228 10776 27232
rect 10712 27172 10716 27228
rect 10716 27172 10772 27228
rect 10772 27172 10776 27228
rect 10712 27168 10776 27172
rect 10792 27228 10856 27232
rect 10792 27172 10796 27228
rect 10796 27172 10852 27228
rect 10852 27172 10856 27228
rect 10792 27168 10856 27172
rect 15352 27228 15416 27232
rect 15352 27172 15356 27228
rect 15356 27172 15412 27228
rect 15412 27172 15416 27228
rect 15352 27168 15416 27172
rect 15432 27228 15496 27232
rect 15432 27172 15436 27228
rect 15436 27172 15492 27228
rect 15492 27172 15496 27228
rect 15432 27168 15496 27172
rect 15512 27228 15576 27232
rect 15512 27172 15516 27228
rect 15516 27172 15572 27228
rect 15572 27172 15576 27228
rect 15512 27168 15576 27172
rect 15592 27228 15656 27232
rect 15592 27172 15596 27228
rect 15596 27172 15652 27228
rect 15652 27172 15656 27228
rect 15592 27168 15656 27172
rect 20152 27228 20216 27232
rect 20152 27172 20156 27228
rect 20156 27172 20212 27228
rect 20212 27172 20216 27228
rect 20152 27168 20216 27172
rect 20232 27228 20296 27232
rect 20232 27172 20236 27228
rect 20236 27172 20292 27228
rect 20292 27172 20296 27228
rect 20232 27168 20296 27172
rect 20312 27228 20376 27232
rect 20312 27172 20316 27228
rect 20316 27172 20372 27228
rect 20372 27172 20376 27228
rect 20312 27168 20376 27172
rect 20392 27228 20456 27232
rect 20392 27172 20396 27228
rect 20396 27172 20452 27228
rect 20452 27172 20456 27228
rect 20392 27168 20456 27172
rect 24952 27228 25016 27232
rect 24952 27172 24956 27228
rect 24956 27172 25012 27228
rect 25012 27172 25016 27228
rect 24952 27168 25016 27172
rect 25032 27228 25096 27232
rect 25032 27172 25036 27228
rect 25036 27172 25092 27228
rect 25092 27172 25096 27228
rect 25032 27168 25096 27172
rect 25112 27228 25176 27232
rect 25112 27172 25116 27228
rect 25116 27172 25172 27228
rect 25172 27172 25176 27228
rect 25112 27168 25176 27172
rect 25192 27228 25256 27232
rect 25192 27172 25196 27228
rect 25196 27172 25252 27228
rect 25252 27172 25256 27228
rect 25192 27168 25256 27172
rect 3352 26684 3416 26688
rect 3352 26628 3356 26684
rect 3356 26628 3412 26684
rect 3412 26628 3416 26684
rect 3352 26624 3416 26628
rect 3432 26684 3496 26688
rect 3432 26628 3436 26684
rect 3436 26628 3492 26684
rect 3492 26628 3496 26684
rect 3432 26624 3496 26628
rect 3512 26684 3576 26688
rect 3512 26628 3516 26684
rect 3516 26628 3572 26684
rect 3572 26628 3576 26684
rect 3512 26624 3576 26628
rect 3592 26684 3656 26688
rect 3592 26628 3596 26684
rect 3596 26628 3652 26684
rect 3652 26628 3656 26684
rect 3592 26624 3656 26628
rect 8152 26684 8216 26688
rect 8152 26628 8156 26684
rect 8156 26628 8212 26684
rect 8212 26628 8216 26684
rect 8152 26624 8216 26628
rect 8232 26684 8296 26688
rect 8232 26628 8236 26684
rect 8236 26628 8292 26684
rect 8292 26628 8296 26684
rect 8232 26624 8296 26628
rect 8312 26684 8376 26688
rect 8312 26628 8316 26684
rect 8316 26628 8372 26684
rect 8372 26628 8376 26684
rect 8312 26624 8376 26628
rect 8392 26684 8456 26688
rect 8392 26628 8396 26684
rect 8396 26628 8452 26684
rect 8452 26628 8456 26684
rect 8392 26624 8456 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 17752 26684 17816 26688
rect 17752 26628 17756 26684
rect 17756 26628 17812 26684
rect 17812 26628 17816 26684
rect 17752 26624 17816 26628
rect 17832 26684 17896 26688
rect 17832 26628 17836 26684
rect 17836 26628 17892 26684
rect 17892 26628 17896 26684
rect 17832 26624 17896 26628
rect 17912 26684 17976 26688
rect 17912 26628 17916 26684
rect 17916 26628 17972 26684
rect 17972 26628 17976 26684
rect 17912 26624 17976 26628
rect 17992 26684 18056 26688
rect 17992 26628 17996 26684
rect 17996 26628 18052 26684
rect 18052 26628 18056 26684
rect 17992 26624 18056 26628
rect 22552 26684 22616 26688
rect 22552 26628 22556 26684
rect 22556 26628 22612 26684
rect 22612 26628 22616 26684
rect 22552 26624 22616 26628
rect 22632 26684 22696 26688
rect 22632 26628 22636 26684
rect 22636 26628 22692 26684
rect 22692 26628 22696 26684
rect 22632 26624 22696 26628
rect 22712 26684 22776 26688
rect 22712 26628 22716 26684
rect 22716 26628 22772 26684
rect 22772 26628 22776 26684
rect 22712 26624 22776 26628
rect 22792 26684 22856 26688
rect 22792 26628 22796 26684
rect 22796 26628 22852 26684
rect 22852 26628 22856 26684
rect 22792 26624 22856 26628
rect 27352 26684 27416 26688
rect 27352 26628 27356 26684
rect 27356 26628 27412 26684
rect 27412 26628 27416 26684
rect 27352 26624 27416 26628
rect 27432 26684 27496 26688
rect 27432 26628 27436 26684
rect 27436 26628 27492 26684
rect 27492 26628 27496 26684
rect 27432 26624 27496 26628
rect 27512 26684 27576 26688
rect 27512 26628 27516 26684
rect 27516 26628 27572 26684
rect 27572 26628 27576 26684
rect 27512 26624 27576 26628
rect 27592 26684 27656 26688
rect 27592 26628 27596 26684
rect 27596 26628 27652 26684
rect 27652 26628 27656 26684
rect 27592 26624 27656 26628
rect 5752 26140 5816 26144
rect 5752 26084 5756 26140
rect 5756 26084 5812 26140
rect 5812 26084 5816 26140
rect 5752 26080 5816 26084
rect 5832 26140 5896 26144
rect 5832 26084 5836 26140
rect 5836 26084 5892 26140
rect 5892 26084 5896 26140
rect 5832 26080 5896 26084
rect 5912 26140 5976 26144
rect 5912 26084 5916 26140
rect 5916 26084 5972 26140
rect 5972 26084 5976 26140
rect 5912 26080 5976 26084
rect 5992 26140 6056 26144
rect 5992 26084 5996 26140
rect 5996 26084 6052 26140
rect 6052 26084 6056 26140
rect 5992 26080 6056 26084
rect 10552 26140 10616 26144
rect 10552 26084 10556 26140
rect 10556 26084 10612 26140
rect 10612 26084 10616 26140
rect 10552 26080 10616 26084
rect 10632 26140 10696 26144
rect 10632 26084 10636 26140
rect 10636 26084 10692 26140
rect 10692 26084 10696 26140
rect 10632 26080 10696 26084
rect 10712 26140 10776 26144
rect 10712 26084 10716 26140
rect 10716 26084 10772 26140
rect 10772 26084 10776 26140
rect 10712 26080 10776 26084
rect 10792 26140 10856 26144
rect 10792 26084 10796 26140
rect 10796 26084 10852 26140
rect 10852 26084 10856 26140
rect 10792 26080 10856 26084
rect 15352 26140 15416 26144
rect 15352 26084 15356 26140
rect 15356 26084 15412 26140
rect 15412 26084 15416 26140
rect 15352 26080 15416 26084
rect 15432 26140 15496 26144
rect 15432 26084 15436 26140
rect 15436 26084 15492 26140
rect 15492 26084 15496 26140
rect 15432 26080 15496 26084
rect 15512 26140 15576 26144
rect 15512 26084 15516 26140
rect 15516 26084 15572 26140
rect 15572 26084 15576 26140
rect 15512 26080 15576 26084
rect 15592 26140 15656 26144
rect 15592 26084 15596 26140
rect 15596 26084 15652 26140
rect 15652 26084 15656 26140
rect 15592 26080 15656 26084
rect 20152 26140 20216 26144
rect 20152 26084 20156 26140
rect 20156 26084 20212 26140
rect 20212 26084 20216 26140
rect 20152 26080 20216 26084
rect 20232 26140 20296 26144
rect 20232 26084 20236 26140
rect 20236 26084 20292 26140
rect 20292 26084 20296 26140
rect 20232 26080 20296 26084
rect 20312 26140 20376 26144
rect 20312 26084 20316 26140
rect 20316 26084 20372 26140
rect 20372 26084 20376 26140
rect 20312 26080 20376 26084
rect 20392 26140 20456 26144
rect 20392 26084 20396 26140
rect 20396 26084 20452 26140
rect 20452 26084 20456 26140
rect 20392 26080 20456 26084
rect 24952 26140 25016 26144
rect 24952 26084 24956 26140
rect 24956 26084 25012 26140
rect 25012 26084 25016 26140
rect 24952 26080 25016 26084
rect 25032 26140 25096 26144
rect 25032 26084 25036 26140
rect 25036 26084 25092 26140
rect 25092 26084 25096 26140
rect 25032 26080 25096 26084
rect 25112 26140 25176 26144
rect 25112 26084 25116 26140
rect 25116 26084 25172 26140
rect 25172 26084 25176 26140
rect 25112 26080 25176 26084
rect 25192 26140 25256 26144
rect 25192 26084 25196 26140
rect 25196 26084 25252 26140
rect 25252 26084 25256 26140
rect 25192 26080 25256 26084
rect 3352 25596 3416 25600
rect 3352 25540 3356 25596
rect 3356 25540 3412 25596
rect 3412 25540 3416 25596
rect 3352 25536 3416 25540
rect 3432 25596 3496 25600
rect 3432 25540 3436 25596
rect 3436 25540 3492 25596
rect 3492 25540 3496 25596
rect 3432 25536 3496 25540
rect 3512 25596 3576 25600
rect 3512 25540 3516 25596
rect 3516 25540 3572 25596
rect 3572 25540 3576 25596
rect 3512 25536 3576 25540
rect 3592 25596 3656 25600
rect 3592 25540 3596 25596
rect 3596 25540 3652 25596
rect 3652 25540 3656 25596
rect 3592 25536 3656 25540
rect 8152 25596 8216 25600
rect 8152 25540 8156 25596
rect 8156 25540 8212 25596
rect 8212 25540 8216 25596
rect 8152 25536 8216 25540
rect 8232 25596 8296 25600
rect 8232 25540 8236 25596
rect 8236 25540 8292 25596
rect 8292 25540 8296 25596
rect 8232 25536 8296 25540
rect 8312 25596 8376 25600
rect 8312 25540 8316 25596
rect 8316 25540 8372 25596
rect 8372 25540 8376 25596
rect 8312 25536 8376 25540
rect 8392 25596 8456 25600
rect 8392 25540 8396 25596
rect 8396 25540 8452 25596
rect 8452 25540 8456 25596
rect 8392 25536 8456 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 17752 25596 17816 25600
rect 17752 25540 17756 25596
rect 17756 25540 17812 25596
rect 17812 25540 17816 25596
rect 17752 25536 17816 25540
rect 17832 25596 17896 25600
rect 17832 25540 17836 25596
rect 17836 25540 17892 25596
rect 17892 25540 17896 25596
rect 17832 25536 17896 25540
rect 17912 25596 17976 25600
rect 17912 25540 17916 25596
rect 17916 25540 17972 25596
rect 17972 25540 17976 25596
rect 17912 25536 17976 25540
rect 17992 25596 18056 25600
rect 17992 25540 17996 25596
rect 17996 25540 18052 25596
rect 18052 25540 18056 25596
rect 17992 25536 18056 25540
rect 22552 25596 22616 25600
rect 22552 25540 22556 25596
rect 22556 25540 22612 25596
rect 22612 25540 22616 25596
rect 22552 25536 22616 25540
rect 22632 25596 22696 25600
rect 22632 25540 22636 25596
rect 22636 25540 22692 25596
rect 22692 25540 22696 25596
rect 22632 25536 22696 25540
rect 22712 25596 22776 25600
rect 22712 25540 22716 25596
rect 22716 25540 22772 25596
rect 22772 25540 22776 25596
rect 22712 25536 22776 25540
rect 22792 25596 22856 25600
rect 22792 25540 22796 25596
rect 22796 25540 22852 25596
rect 22852 25540 22856 25596
rect 22792 25536 22856 25540
rect 27352 25596 27416 25600
rect 27352 25540 27356 25596
rect 27356 25540 27412 25596
rect 27412 25540 27416 25596
rect 27352 25536 27416 25540
rect 27432 25596 27496 25600
rect 27432 25540 27436 25596
rect 27436 25540 27492 25596
rect 27492 25540 27496 25596
rect 27432 25536 27496 25540
rect 27512 25596 27576 25600
rect 27512 25540 27516 25596
rect 27516 25540 27572 25596
rect 27572 25540 27576 25596
rect 27512 25536 27576 25540
rect 27592 25596 27656 25600
rect 27592 25540 27596 25596
rect 27596 25540 27652 25596
rect 27652 25540 27656 25596
rect 27592 25536 27656 25540
rect 5752 25052 5816 25056
rect 5752 24996 5756 25052
rect 5756 24996 5812 25052
rect 5812 24996 5816 25052
rect 5752 24992 5816 24996
rect 5832 25052 5896 25056
rect 5832 24996 5836 25052
rect 5836 24996 5892 25052
rect 5892 24996 5896 25052
rect 5832 24992 5896 24996
rect 5912 25052 5976 25056
rect 5912 24996 5916 25052
rect 5916 24996 5972 25052
rect 5972 24996 5976 25052
rect 5912 24992 5976 24996
rect 5992 25052 6056 25056
rect 5992 24996 5996 25052
rect 5996 24996 6052 25052
rect 6052 24996 6056 25052
rect 5992 24992 6056 24996
rect 10552 25052 10616 25056
rect 10552 24996 10556 25052
rect 10556 24996 10612 25052
rect 10612 24996 10616 25052
rect 10552 24992 10616 24996
rect 10632 25052 10696 25056
rect 10632 24996 10636 25052
rect 10636 24996 10692 25052
rect 10692 24996 10696 25052
rect 10632 24992 10696 24996
rect 10712 25052 10776 25056
rect 10712 24996 10716 25052
rect 10716 24996 10772 25052
rect 10772 24996 10776 25052
rect 10712 24992 10776 24996
rect 10792 25052 10856 25056
rect 10792 24996 10796 25052
rect 10796 24996 10852 25052
rect 10852 24996 10856 25052
rect 10792 24992 10856 24996
rect 15352 25052 15416 25056
rect 15352 24996 15356 25052
rect 15356 24996 15412 25052
rect 15412 24996 15416 25052
rect 15352 24992 15416 24996
rect 15432 25052 15496 25056
rect 15432 24996 15436 25052
rect 15436 24996 15492 25052
rect 15492 24996 15496 25052
rect 15432 24992 15496 24996
rect 15512 25052 15576 25056
rect 15512 24996 15516 25052
rect 15516 24996 15572 25052
rect 15572 24996 15576 25052
rect 15512 24992 15576 24996
rect 15592 25052 15656 25056
rect 15592 24996 15596 25052
rect 15596 24996 15652 25052
rect 15652 24996 15656 25052
rect 15592 24992 15656 24996
rect 20152 25052 20216 25056
rect 20152 24996 20156 25052
rect 20156 24996 20212 25052
rect 20212 24996 20216 25052
rect 20152 24992 20216 24996
rect 20232 25052 20296 25056
rect 20232 24996 20236 25052
rect 20236 24996 20292 25052
rect 20292 24996 20296 25052
rect 20232 24992 20296 24996
rect 20312 25052 20376 25056
rect 20312 24996 20316 25052
rect 20316 24996 20372 25052
rect 20372 24996 20376 25052
rect 20312 24992 20376 24996
rect 20392 25052 20456 25056
rect 20392 24996 20396 25052
rect 20396 24996 20452 25052
rect 20452 24996 20456 25052
rect 20392 24992 20456 24996
rect 24952 25052 25016 25056
rect 24952 24996 24956 25052
rect 24956 24996 25012 25052
rect 25012 24996 25016 25052
rect 24952 24992 25016 24996
rect 25032 25052 25096 25056
rect 25032 24996 25036 25052
rect 25036 24996 25092 25052
rect 25092 24996 25096 25052
rect 25032 24992 25096 24996
rect 25112 25052 25176 25056
rect 25112 24996 25116 25052
rect 25116 24996 25172 25052
rect 25172 24996 25176 25052
rect 25112 24992 25176 24996
rect 25192 25052 25256 25056
rect 25192 24996 25196 25052
rect 25196 24996 25252 25052
rect 25252 24996 25256 25052
rect 25192 24992 25256 24996
rect 3352 24508 3416 24512
rect 3352 24452 3356 24508
rect 3356 24452 3412 24508
rect 3412 24452 3416 24508
rect 3352 24448 3416 24452
rect 3432 24508 3496 24512
rect 3432 24452 3436 24508
rect 3436 24452 3492 24508
rect 3492 24452 3496 24508
rect 3432 24448 3496 24452
rect 3512 24508 3576 24512
rect 3512 24452 3516 24508
rect 3516 24452 3572 24508
rect 3572 24452 3576 24508
rect 3512 24448 3576 24452
rect 3592 24508 3656 24512
rect 3592 24452 3596 24508
rect 3596 24452 3652 24508
rect 3652 24452 3656 24508
rect 3592 24448 3656 24452
rect 8152 24508 8216 24512
rect 8152 24452 8156 24508
rect 8156 24452 8212 24508
rect 8212 24452 8216 24508
rect 8152 24448 8216 24452
rect 8232 24508 8296 24512
rect 8232 24452 8236 24508
rect 8236 24452 8292 24508
rect 8292 24452 8296 24508
rect 8232 24448 8296 24452
rect 8312 24508 8376 24512
rect 8312 24452 8316 24508
rect 8316 24452 8372 24508
rect 8372 24452 8376 24508
rect 8312 24448 8376 24452
rect 8392 24508 8456 24512
rect 8392 24452 8396 24508
rect 8396 24452 8452 24508
rect 8452 24452 8456 24508
rect 8392 24448 8456 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 17752 24508 17816 24512
rect 17752 24452 17756 24508
rect 17756 24452 17812 24508
rect 17812 24452 17816 24508
rect 17752 24448 17816 24452
rect 17832 24508 17896 24512
rect 17832 24452 17836 24508
rect 17836 24452 17892 24508
rect 17892 24452 17896 24508
rect 17832 24448 17896 24452
rect 17912 24508 17976 24512
rect 17912 24452 17916 24508
rect 17916 24452 17972 24508
rect 17972 24452 17976 24508
rect 17912 24448 17976 24452
rect 17992 24508 18056 24512
rect 17992 24452 17996 24508
rect 17996 24452 18052 24508
rect 18052 24452 18056 24508
rect 17992 24448 18056 24452
rect 22552 24508 22616 24512
rect 22552 24452 22556 24508
rect 22556 24452 22612 24508
rect 22612 24452 22616 24508
rect 22552 24448 22616 24452
rect 22632 24508 22696 24512
rect 22632 24452 22636 24508
rect 22636 24452 22692 24508
rect 22692 24452 22696 24508
rect 22632 24448 22696 24452
rect 22712 24508 22776 24512
rect 22712 24452 22716 24508
rect 22716 24452 22772 24508
rect 22772 24452 22776 24508
rect 22712 24448 22776 24452
rect 22792 24508 22856 24512
rect 22792 24452 22796 24508
rect 22796 24452 22852 24508
rect 22852 24452 22856 24508
rect 22792 24448 22856 24452
rect 27352 24508 27416 24512
rect 27352 24452 27356 24508
rect 27356 24452 27412 24508
rect 27412 24452 27416 24508
rect 27352 24448 27416 24452
rect 27432 24508 27496 24512
rect 27432 24452 27436 24508
rect 27436 24452 27492 24508
rect 27492 24452 27496 24508
rect 27432 24448 27496 24452
rect 27512 24508 27576 24512
rect 27512 24452 27516 24508
rect 27516 24452 27572 24508
rect 27572 24452 27576 24508
rect 27512 24448 27576 24452
rect 27592 24508 27656 24512
rect 27592 24452 27596 24508
rect 27596 24452 27652 24508
rect 27652 24452 27656 24508
rect 27592 24448 27656 24452
rect 5752 23964 5816 23968
rect 5752 23908 5756 23964
rect 5756 23908 5812 23964
rect 5812 23908 5816 23964
rect 5752 23904 5816 23908
rect 5832 23964 5896 23968
rect 5832 23908 5836 23964
rect 5836 23908 5892 23964
rect 5892 23908 5896 23964
rect 5832 23904 5896 23908
rect 5912 23964 5976 23968
rect 5912 23908 5916 23964
rect 5916 23908 5972 23964
rect 5972 23908 5976 23964
rect 5912 23904 5976 23908
rect 5992 23964 6056 23968
rect 5992 23908 5996 23964
rect 5996 23908 6052 23964
rect 6052 23908 6056 23964
rect 5992 23904 6056 23908
rect 10552 23964 10616 23968
rect 10552 23908 10556 23964
rect 10556 23908 10612 23964
rect 10612 23908 10616 23964
rect 10552 23904 10616 23908
rect 10632 23964 10696 23968
rect 10632 23908 10636 23964
rect 10636 23908 10692 23964
rect 10692 23908 10696 23964
rect 10632 23904 10696 23908
rect 10712 23964 10776 23968
rect 10712 23908 10716 23964
rect 10716 23908 10772 23964
rect 10772 23908 10776 23964
rect 10712 23904 10776 23908
rect 10792 23964 10856 23968
rect 10792 23908 10796 23964
rect 10796 23908 10852 23964
rect 10852 23908 10856 23964
rect 10792 23904 10856 23908
rect 15352 23964 15416 23968
rect 15352 23908 15356 23964
rect 15356 23908 15412 23964
rect 15412 23908 15416 23964
rect 15352 23904 15416 23908
rect 15432 23964 15496 23968
rect 15432 23908 15436 23964
rect 15436 23908 15492 23964
rect 15492 23908 15496 23964
rect 15432 23904 15496 23908
rect 15512 23964 15576 23968
rect 15512 23908 15516 23964
rect 15516 23908 15572 23964
rect 15572 23908 15576 23964
rect 15512 23904 15576 23908
rect 15592 23964 15656 23968
rect 15592 23908 15596 23964
rect 15596 23908 15652 23964
rect 15652 23908 15656 23964
rect 15592 23904 15656 23908
rect 20152 23964 20216 23968
rect 20152 23908 20156 23964
rect 20156 23908 20212 23964
rect 20212 23908 20216 23964
rect 20152 23904 20216 23908
rect 20232 23964 20296 23968
rect 20232 23908 20236 23964
rect 20236 23908 20292 23964
rect 20292 23908 20296 23964
rect 20232 23904 20296 23908
rect 20312 23964 20376 23968
rect 20312 23908 20316 23964
rect 20316 23908 20372 23964
rect 20372 23908 20376 23964
rect 20312 23904 20376 23908
rect 20392 23964 20456 23968
rect 20392 23908 20396 23964
rect 20396 23908 20452 23964
rect 20452 23908 20456 23964
rect 20392 23904 20456 23908
rect 24952 23964 25016 23968
rect 24952 23908 24956 23964
rect 24956 23908 25012 23964
rect 25012 23908 25016 23964
rect 24952 23904 25016 23908
rect 25032 23964 25096 23968
rect 25032 23908 25036 23964
rect 25036 23908 25092 23964
rect 25092 23908 25096 23964
rect 25032 23904 25096 23908
rect 25112 23964 25176 23968
rect 25112 23908 25116 23964
rect 25116 23908 25172 23964
rect 25172 23908 25176 23964
rect 25112 23904 25176 23908
rect 25192 23964 25256 23968
rect 25192 23908 25196 23964
rect 25196 23908 25252 23964
rect 25252 23908 25256 23964
rect 25192 23904 25256 23908
rect 3352 23420 3416 23424
rect 3352 23364 3356 23420
rect 3356 23364 3412 23420
rect 3412 23364 3416 23420
rect 3352 23360 3416 23364
rect 3432 23420 3496 23424
rect 3432 23364 3436 23420
rect 3436 23364 3492 23420
rect 3492 23364 3496 23420
rect 3432 23360 3496 23364
rect 3512 23420 3576 23424
rect 3512 23364 3516 23420
rect 3516 23364 3572 23420
rect 3572 23364 3576 23420
rect 3512 23360 3576 23364
rect 3592 23420 3656 23424
rect 3592 23364 3596 23420
rect 3596 23364 3652 23420
rect 3652 23364 3656 23420
rect 3592 23360 3656 23364
rect 8152 23420 8216 23424
rect 8152 23364 8156 23420
rect 8156 23364 8212 23420
rect 8212 23364 8216 23420
rect 8152 23360 8216 23364
rect 8232 23420 8296 23424
rect 8232 23364 8236 23420
rect 8236 23364 8292 23420
rect 8292 23364 8296 23420
rect 8232 23360 8296 23364
rect 8312 23420 8376 23424
rect 8312 23364 8316 23420
rect 8316 23364 8372 23420
rect 8372 23364 8376 23420
rect 8312 23360 8376 23364
rect 8392 23420 8456 23424
rect 8392 23364 8396 23420
rect 8396 23364 8452 23420
rect 8452 23364 8456 23420
rect 8392 23360 8456 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 17752 23420 17816 23424
rect 17752 23364 17756 23420
rect 17756 23364 17812 23420
rect 17812 23364 17816 23420
rect 17752 23360 17816 23364
rect 17832 23420 17896 23424
rect 17832 23364 17836 23420
rect 17836 23364 17892 23420
rect 17892 23364 17896 23420
rect 17832 23360 17896 23364
rect 17912 23420 17976 23424
rect 17912 23364 17916 23420
rect 17916 23364 17972 23420
rect 17972 23364 17976 23420
rect 17912 23360 17976 23364
rect 17992 23420 18056 23424
rect 17992 23364 17996 23420
rect 17996 23364 18052 23420
rect 18052 23364 18056 23420
rect 17992 23360 18056 23364
rect 22552 23420 22616 23424
rect 22552 23364 22556 23420
rect 22556 23364 22612 23420
rect 22612 23364 22616 23420
rect 22552 23360 22616 23364
rect 22632 23420 22696 23424
rect 22632 23364 22636 23420
rect 22636 23364 22692 23420
rect 22692 23364 22696 23420
rect 22632 23360 22696 23364
rect 22712 23420 22776 23424
rect 22712 23364 22716 23420
rect 22716 23364 22772 23420
rect 22772 23364 22776 23420
rect 22712 23360 22776 23364
rect 22792 23420 22856 23424
rect 22792 23364 22796 23420
rect 22796 23364 22852 23420
rect 22852 23364 22856 23420
rect 22792 23360 22856 23364
rect 27352 23420 27416 23424
rect 27352 23364 27356 23420
rect 27356 23364 27412 23420
rect 27412 23364 27416 23420
rect 27352 23360 27416 23364
rect 27432 23420 27496 23424
rect 27432 23364 27436 23420
rect 27436 23364 27492 23420
rect 27492 23364 27496 23420
rect 27432 23360 27496 23364
rect 27512 23420 27576 23424
rect 27512 23364 27516 23420
rect 27516 23364 27572 23420
rect 27572 23364 27576 23420
rect 27512 23360 27576 23364
rect 27592 23420 27656 23424
rect 27592 23364 27596 23420
rect 27596 23364 27652 23420
rect 27652 23364 27656 23420
rect 27592 23360 27656 23364
rect 5752 22876 5816 22880
rect 5752 22820 5756 22876
rect 5756 22820 5812 22876
rect 5812 22820 5816 22876
rect 5752 22816 5816 22820
rect 5832 22876 5896 22880
rect 5832 22820 5836 22876
rect 5836 22820 5892 22876
rect 5892 22820 5896 22876
rect 5832 22816 5896 22820
rect 5912 22876 5976 22880
rect 5912 22820 5916 22876
rect 5916 22820 5972 22876
rect 5972 22820 5976 22876
rect 5912 22816 5976 22820
rect 5992 22876 6056 22880
rect 5992 22820 5996 22876
rect 5996 22820 6052 22876
rect 6052 22820 6056 22876
rect 5992 22816 6056 22820
rect 10552 22876 10616 22880
rect 10552 22820 10556 22876
rect 10556 22820 10612 22876
rect 10612 22820 10616 22876
rect 10552 22816 10616 22820
rect 10632 22876 10696 22880
rect 10632 22820 10636 22876
rect 10636 22820 10692 22876
rect 10692 22820 10696 22876
rect 10632 22816 10696 22820
rect 10712 22876 10776 22880
rect 10712 22820 10716 22876
rect 10716 22820 10772 22876
rect 10772 22820 10776 22876
rect 10712 22816 10776 22820
rect 10792 22876 10856 22880
rect 10792 22820 10796 22876
rect 10796 22820 10852 22876
rect 10852 22820 10856 22876
rect 10792 22816 10856 22820
rect 15352 22876 15416 22880
rect 15352 22820 15356 22876
rect 15356 22820 15412 22876
rect 15412 22820 15416 22876
rect 15352 22816 15416 22820
rect 15432 22876 15496 22880
rect 15432 22820 15436 22876
rect 15436 22820 15492 22876
rect 15492 22820 15496 22876
rect 15432 22816 15496 22820
rect 15512 22876 15576 22880
rect 15512 22820 15516 22876
rect 15516 22820 15572 22876
rect 15572 22820 15576 22876
rect 15512 22816 15576 22820
rect 15592 22876 15656 22880
rect 15592 22820 15596 22876
rect 15596 22820 15652 22876
rect 15652 22820 15656 22876
rect 15592 22816 15656 22820
rect 20152 22876 20216 22880
rect 20152 22820 20156 22876
rect 20156 22820 20212 22876
rect 20212 22820 20216 22876
rect 20152 22816 20216 22820
rect 20232 22876 20296 22880
rect 20232 22820 20236 22876
rect 20236 22820 20292 22876
rect 20292 22820 20296 22876
rect 20232 22816 20296 22820
rect 20312 22876 20376 22880
rect 20312 22820 20316 22876
rect 20316 22820 20372 22876
rect 20372 22820 20376 22876
rect 20312 22816 20376 22820
rect 20392 22876 20456 22880
rect 20392 22820 20396 22876
rect 20396 22820 20452 22876
rect 20452 22820 20456 22876
rect 20392 22816 20456 22820
rect 24952 22876 25016 22880
rect 24952 22820 24956 22876
rect 24956 22820 25012 22876
rect 25012 22820 25016 22876
rect 24952 22816 25016 22820
rect 25032 22876 25096 22880
rect 25032 22820 25036 22876
rect 25036 22820 25092 22876
rect 25092 22820 25096 22876
rect 25032 22816 25096 22820
rect 25112 22876 25176 22880
rect 25112 22820 25116 22876
rect 25116 22820 25172 22876
rect 25172 22820 25176 22876
rect 25112 22816 25176 22820
rect 25192 22876 25256 22880
rect 25192 22820 25196 22876
rect 25196 22820 25252 22876
rect 25252 22820 25256 22876
rect 25192 22816 25256 22820
rect 3352 22332 3416 22336
rect 3352 22276 3356 22332
rect 3356 22276 3412 22332
rect 3412 22276 3416 22332
rect 3352 22272 3416 22276
rect 3432 22332 3496 22336
rect 3432 22276 3436 22332
rect 3436 22276 3492 22332
rect 3492 22276 3496 22332
rect 3432 22272 3496 22276
rect 3512 22332 3576 22336
rect 3512 22276 3516 22332
rect 3516 22276 3572 22332
rect 3572 22276 3576 22332
rect 3512 22272 3576 22276
rect 3592 22332 3656 22336
rect 3592 22276 3596 22332
rect 3596 22276 3652 22332
rect 3652 22276 3656 22332
rect 3592 22272 3656 22276
rect 8152 22332 8216 22336
rect 8152 22276 8156 22332
rect 8156 22276 8212 22332
rect 8212 22276 8216 22332
rect 8152 22272 8216 22276
rect 8232 22332 8296 22336
rect 8232 22276 8236 22332
rect 8236 22276 8292 22332
rect 8292 22276 8296 22332
rect 8232 22272 8296 22276
rect 8312 22332 8376 22336
rect 8312 22276 8316 22332
rect 8316 22276 8372 22332
rect 8372 22276 8376 22332
rect 8312 22272 8376 22276
rect 8392 22332 8456 22336
rect 8392 22276 8396 22332
rect 8396 22276 8452 22332
rect 8452 22276 8456 22332
rect 8392 22272 8456 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 17752 22332 17816 22336
rect 17752 22276 17756 22332
rect 17756 22276 17812 22332
rect 17812 22276 17816 22332
rect 17752 22272 17816 22276
rect 17832 22332 17896 22336
rect 17832 22276 17836 22332
rect 17836 22276 17892 22332
rect 17892 22276 17896 22332
rect 17832 22272 17896 22276
rect 17912 22332 17976 22336
rect 17912 22276 17916 22332
rect 17916 22276 17972 22332
rect 17972 22276 17976 22332
rect 17912 22272 17976 22276
rect 17992 22332 18056 22336
rect 17992 22276 17996 22332
rect 17996 22276 18052 22332
rect 18052 22276 18056 22332
rect 17992 22272 18056 22276
rect 22552 22332 22616 22336
rect 22552 22276 22556 22332
rect 22556 22276 22612 22332
rect 22612 22276 22616 22332
rect 22552 22272 22616 22276
rect 22632 22332 22696 22336
rect 22632 22276 22636 22332
rect 22636 22276 22692 22332
rect 22692 22276 22696 22332
rect 22632 22272 22696 22276
rect 22712 22332 22776 22336
rect 22712 22276 22716 22332
rect 22716 22276 22772 22332
rect 22772 22276 22776 22332
rect 22712 22272 22776 22276
rect 22792 22332 22856 22336
rect 22792 22276 22796 22332
rect 22796 22276 22852 22332
rect 22852 22276 22856 22332
rect 22792 22272 22856 22276
rect 27352 22332 27416 22336
rect 27352 22276 27356 22332
rect 27356 22276 27412 22332
rect 27412 22276 27416 22332
rect 27352 22272 27416 22276
rect 27432 22332 27496 22336
rect 27432 22276 27436 22332
rect 27436 22276 27492 22332
rect 27492 22276 27496 22332
rect 27432 22272 27496 22276
rect 27512 22332 27576 22336
rect 27512 22276 27516 22332
rect 27516 22276 27572 22332
rect 27572 22276 27576 22332
rect 27512 22272 27576 22276
rect 27592 22332 27656 22336
rect 27592 22276 27596 22332
rect 27596 22276 27652 22332
rect 27652 22276 27656 22332
rect 27592 22272 27656 22276
rect 5752 21788 5816 21792
rect 5752 21732 5756 21788
rect 5756 21732 5812 21788
rect 5812 21732 5816 21788
rect 5752 21728 5816 21732
rect 5832 21788 5896 21792
rect 5832 21732 5836 21788
rect 5836 21732 5892 21788
rect 5892 21732 5896 21788
rect 5832 21728 5896 21732
rect 5912 21788 5976 21792
rect 5912 21732 5916 21788
rect 5916 21732 5972 21788
rect 5972 21732 5976 21788
rect 5912 21728 5976 21732
rect 5992 21788 6056 21792
rect 5992 21732 5996 21788
rect 5996 21732 6052 21788
rect 6052 21732 6056 21788
rect 5992 21728 6056 21732
rect 10552 21788 10616 21792
rect 10552 21732 10556 21788
rect 10556 21732 10612 21788
rect 10612 21732 10616 21788
rect 10552 21728 10616 21732
rect 10632 21788 10696 21792
rect 10632 21732 10636 21788
rect 10636 21732 10692 21788
rect 10692 21732 10696 21788
rect 10632 21728 10696 21732
rect 10712 21788 10776 21792
rect 10712 21732 10716 21788
rect 10716 21732 10772 21788
rect 10772 21732 10776 21788
rect 10712 21728 10776 21732
rect 10792 21788 10856 21792
rect 10792 21732 10796 21788
rect 10796 21732 10852 21788
rect 10852 21732 10856 21788
rect 10792 21728 10856 21732
rect 15352 21788 15416 21792
rect 15352 21732 15356 21788
rect 15356 21732 15412 21788
rect 15412 21732 15416 21788
rect 15352 21728 15416 21732
rect 15432 21788 15496 21792
rect 15432 21732 15436 21788
rect 15436 21732 15492 21788
rect 15492 21732 15496 21788
rect 15432 21728 15496 21732
rect 15512 21788 15576 21792
rect 15512 21732 15516 21788
rect 15516 21732 15572 21788
rect 15572 21732 15576 21788
rect 15512 21728 15576 21732
rect 15592 21788 15656 21792
rect 15592 21732 15596 21788
rect 15596 21732 15652 21788
rect 15652 21732 15656 21788
rect 15592 21728 15656 21732
rect 20152 21788 20216 21792
rect 20152 21732 20156 21788
rect 20156 21732 20212 21788
rect 20212 21732 20216 21788
rect 20152 21728 20216 21732
rect 20232 21788 20296 21792
rect 20232 21732 20236 21788
rect 20236 21732 20292 21788
rect 20292 21732 20296 21788
rect 20232 21728 20296 21732
rect 20312 21788 20376 21792
rect 20312 21732 20316 21788
rect 20316 21732 20372 21788
rect 20372 21732 20376 21788
rect 20312 21728 20376 21732
rect 20392 21788 20456 21792
rect 20392 21732 20396 21788
rect 20396 21732 20452 21788
rect 20452 21732 20456 21788
rect 20392 21728 20456 21732
rect 24952 21788 25016 21792
rect 24952 21732 24956 21788
rect 24956 21732 25012 21788
rect 25012 21732 25016 21788
rect 24952 21728 25016 21732
rect 25032 21788 25096 21792
rect 25032 21732 25036 21788
rect 25036 21732 25092 21788
rect 25092 21732 25096 21788
rect 25032 21728 25096 21732
rect 25112 21788 25176 21792
rect 25112 21732 25116 21788
rect 25116 21732 25172 21788
rect 25172 21732 25176 21788
rect 25112 21728 25176 21732
rect 25192 21788 25256 21792
rect 25192 21732 25196 21788
rect 25196 21732 25252 21788
rect 25252 21732 25256 21788
rect 25192 21728 25256 21732
rect 3352 21244 3416 21248
rect 3352 21188 3356 21244
rect 3356 21188 3412 21244
rect 3412 21188 3416 21244
rect 3352 21184 3416 21188
rect 3432 21244 3496 21248
rect 3432 21188 3436 21244
rect 3436 21188 3492 21244
rect 3492 21188 3496 21244
rect 3432 21184 3496 21188
rect 3512 21244 3576 21248
rect 3512 21188 3516 21244
rect 3516 21188 3572 21244
rect 3572 21188 3576 21244
rect 3512 21184 3576 21188
rect 3592 21244 3656 21248
rect 3592 21188 3596 21244
rect 3596 21188 3652 21244
rect 3652 21188 3656 21244
rect 3592 21184 3656 21188
rect 8152 21244 8216 21248
rect 8152 21188 8156 21244
rect 8156 21188 8212 21244
rect 8212 21188 8216 21244
rect 8152 21184 8216 21188
rect 8232 21244 8296 21248
rect 8232 21188 8236 21244
rect 8236 21188 8292 21244
rect 8292 21188 8296 21244
rect 8232 21184 8296 21188
rect 8312 21244 8376 21248
rect 8312 21188 8316 21244
rect 8316 21188 8372 21244
rect 8372 21188 8376 21244
rect 8312 21184 8376 21188
rect 8392 21244 8456 21248
rect 8392 21188 8396 21244
rect 8396 21188 8452 21244
rect 8452 21188 8456 21244
rect 8392 21184 8456 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 17752 21244 17816 21248
rect 17752 21188 17756 21244
rect 17756 21188 17812 21244
rect 17812 21188 17816 21244
rect 17752 21184 17816 21188
rect 17832 21244 17896 21248
rect 17832 21188 17836 21244
rect 17836 21188 17892 21244
rect 17892 21188 17896 21244
rect 17832 21184 17896 21188
rect 17912 21244 17976 21248
rect 17912 21188 17916 21244
rect 17916 21188 17972 21244
rect 17972 21188 17976 21244
rect 17912 21184 17976 21188
rect 17992 21244 18056 21248
rect 17992 21188 17996 21244
rect 17996 21188 18052 21244
rect 18052 21188 18056 21244
rect 17992 21184 18056 21188
rect 22552 21244 22616 21248
rect 22552 21188 22556 21244
rect 22556 21188 22612 21244
rect 22612 21188 22616 21244
rect 22552 21184 22616 21188
rect 22632 21244 22696 21248
rect 22632 21188 22636 21244
rect 22636 21188 22692 21244
rect 22692 21188 22696 21244
rect 22632 21184 22696 21188
rect 22712 21244 22776 21248
rect 22712 21188 22716 21244
rect 22716 21188 22772 21244
rect 22772 21188 22776 21244
rect 22712 21184 22776 21188
rect 22792 21244 22856 21248
rect 22792 21188 22796 21244
rect 22796 21188 22852 21244
rect 22852 21188 22856 21244
rect 22792 21184 22856 21188
rect 27352 21244 27416 21248
rect 27352 21188 27356 21244
rect 27356 21188 27412 21244
rect 27412 21188 27416 21244
rect 27352 21184 27416 21188
rect 27432 21244 27496 21248
rect 27432 21188 27436 21244
rect 27436 21188 27492 21244
rect 27492 21188 27496 21244
rect 27432 21184 27496 21188
rect 27512 21244 27576 21248
rect 27512 21188 27516 21244
rect 27516 21188 27572 21244
rect 27572 21188 27576 21244
rect 27512 21184 27576 21188
rect 27592 21244 27656 21248
rect 27592 21188 27596 21244
rect 27596 21188 27652 21244
rect 27652 21188 27656 21244
rect 27592 21184 27656 21188
rect 5752 20700 5816 20704
rect 5752 20644 5756 20700
rect 5756 20644 5812 20700
rect 5812 20644 5816 20700
rect 5752 20640 5816 20644
rect 5832 20700 5896 20704
rect 5832 20644 5836 20700
rect 5836 20644 5892 20700
rect 5892 20644 5896 20700
rect 5832 20640 5896 20644
rect 5912 20700 5976 20704
rect 5912 20644 5916 20700
rect 5916 20644 5972 20700
rect 5972 20644 5976 20700
rect 5912 20640 5976 20644
rect 5992 20700 6056 20704
rect 5992 20644 5996 20700
rect 5996 20644 6052 20700
rect 6052 20644 6056 20700
rect 5992 20640 6056 20644
rect 10552 20700 10616 20704
rect 10552 20644 10556 20700
rect 10556 20644 10612 20700
rect 10612 20644 10616 20700
rect 10552 20640 10616 20644
rect 10632 20700 10696 20704
rect 10632 20644 10636 20700
rect 10636 20644 10692 20700
rect 10692 20644 10696 20700
rect 10632 20640 10696 20644
rect 10712 20700 10776 20704
rect 10712 20644 10716 20700
rect 10716 20644 10772 20700
rect 10772 20644 10776 20700
rect 10712 20640 10776 20644
rect 10792 20700 10856 20704
rect 10792 20644 10796 20700
rect 10796 20644 10852 20700
rect 10852 20644 10856 20700
rect 10792 20640 10856 20644
rect 15352 20700 15416 20704
rect 15352 20644 15356 20700
rect 15356 20644 15412 20700
rect 15412 20644 15416 20700
rect 15352 20640 15416 20644
rect 15432 20700 15496 20704
rect 15432 20644 15436 20700
rect 15436 20644 15492 20700
rect 15492 20644 15496 20700
rect 15432 20640 15496 20644
rect 15512 20700 15576 20704
rect 15512 20644 15516 20700
rect 15516 20644 15572 20700
rect 15572 20644 15576 20700
rect 15512 20640 15576 20644
rect 15592 20700 15656 20704
rect 15592 20644 15596 20700
rect 15596 20644 15652 20700
rect 15652 20644 15656 20700
rect 15592 20640 15656 20644
rect 20152 20700 20216 20704
rect 20152 20644 20156 20700
rect 20156 20644 20212 20700
rect 20212 20644 20216 20700
rect 20152 20640 20216 20644
rect 20232 20700 20296 20704
rect 20232 20644 20236 20700
rect 20236 20644 20292 20700
rect 20292 20644 20296 20700
rect 20232 20640 20296 20644
rect 20312 20700 20376 20704
rect 20312 20644 20316 20700
rect 20316 20644 20372 20700
rect 20372 20644 20376 20700
rect 20312 20640 20376 20644
rect 20392 20700 20456 20704
rect 20392 20644 20396 20700
rect 20396 20644 20452 20700
rect 20452 20644 20456 20700
rect 20392 20640 20456 20644
rect 24952 20700 25016 20704
rect 24952 20644 24956 20700
rect 24956 20644 25012 20700
rect 25012 20644 25016 20700
rect 24952 20640 25016 20644
rect 25032 20700 25096 20704
rect 25032 20644 25036 20700
rect 25036 20644 25092 20700
rect 25092 20644 25096 20700
rect 25032 20640 25096 20644
rect 25112 20700 25176 20704
rect 25112 20644 25116 20700
rect 25116 20644 25172 20700
rect 25172 20644 25176 20700
rect 25112 20640 25176 20644
rect 25192 20700 25256 20704
rect 25192 20644 25196 20700
rect 25196 20644 25252 20700
rect 25252 20644 25256 20700
rect 25192 20640 25256 20644
rect 3352 20156 3416 20160
rect 3352 20100 3356 20156
rect 3356 20100 3412 20156
rect 3412 20100 3416 20156
rect 3352 20096 3416 20100
rect 3432 20156 3496 20160
rect 3432 20100 3436 20156
rect 3436 20100 3492 20156
rect 3492 20100 3496 20156
rect 3432 20096 3496 20100
rect 3512 20156 3576 20160
rect 3512 20100 3516 20156
rect 3516 20100 3572 20156
rect 3572 20100 3576 20156
rect 3512 20096 3576 20100
rect 3592 20156 3656 20160
rect 3592 20100 3596 20156
rect 3596 20100 3652 20156
rect 3652 20100 3656 20156
rect 3592 20096 3656 20100
rect 8152 20156 8216 20160
rect 8152 20100 8156 20156
rect 8156 20100 8212 20156
rect 8212 20100 8216 20156
rect 8152 20096 8216 20100
rect 8232 20156 8296 20160
rect 8232 20100 8236 20156
rect 8236 20100 8292 20156
rect 8292 20100 8296 20156
rect 8232 20096 8296 20100
rect 8312 20156 8376 20160
rect 8312 20100 8316 20156
rect 8316 20100 8372 20156
rect 8372 20100 8376 20156
rect 8312 20096 8376 20100
rect 8392 20156 8456 20160
rect 8392 20100 8396 20156
rect 8396 20100 8452 20156
rect 8452 20100 8456 20156
rect 8392 20096 8456 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 17752 20156 17816 20160
rect 17752 20100 17756 20156
rect 17756 20100 17812 20156
rect 17812 20100 17816 20156
rect 17752 20096 17816 20100
rect 17832 20156 17896 20160
rect 17832 20100 17836 20156
rect 17836 20100 17892 20156
rect 17892 20100 17896 20156
rect 17832 20096 17896 20100
rect 17912 20156 17976 20160
rect 17912 20100 17916 20156
rect 17916 20100 17972 20156
rect 17972 20100 17976 20156
rect 17912 20096 17976 20100
rect 17992 20156 18056 20160
rect 17992 20100 17996 20156
rect 17996 20100 18052 20156
rect 18052 20100 18056 20156
rect 17992 20096 18056 20100
rect 22552 20156 22616 20160
rect 22552 20100 22556 20156
rect 22556 20100 22612 20156
rect 22612 20100 22616 20156
rect 22552 20096 22616 20100
rect 22632 20156 22696 20160
rect 22632 20100 22636 20156
rect 22636 20100 22692 20156
rect 22692 20100 22696 20156
rect 22632 20096 22696 20100
rect 22712 20156 22776 20160
rect 22712 20100 22716 20156
rect 22716 20100 22772 20156
rect 22772 20100 22776 20156
rect 22712 20096 22776 20100
rect 22792 20156 22856 20160
rect 22792 20100 22796 20156
rect 22796 20100 22852 20156
rect 22852 20100 22856 20156
rect 22792 20096 22856 20100
rect 27352 20156 27416 20160
rect 27352 20100 27356 20156
rect 27356 20100 27412 20156
rect 27412 20100 27416 20156
rect 27352 20096 27416 20100
rect 27432 20156 27496 20160
rect 27432 20100 27436 20156
rect 27436 20100 27492 20156
rect 27492 20100 27496 20156
rect 27432 20096 27496 20100
rect 27512 20156 27576 20160
rect 27512 20100 27516 20156
rect 27516 20100 27572 20156
rect 27572 20100 27576 20156
rect 27512 20096 27576 20100
rect 27592 20156 27656 20160
rect 27592 20100 27596 20156
rect 27596 20100 27652 20156
rect 27652 20100 27656 20156
rect 27592 20096 27656 20100
rect 5752 19612 5816 19616
rect 5752 19556 5756 19612
rect 5756 19556 5812 19612
rect 5812 19556 5816 19612
rect 5752 19552 5816 19556
rect 5832 19612 5896 19616
rect 5832 19556 5836 19612
rect 5836 19556 5892 19612
rect 5892 19556 5896 19612
rect 5832 19552 5896 19556
rect 5912 19612 5976 19616
rect 5912 19556 5916 19612
rect 5916 19556 5972 19612
rect 5972 19556 5976 19612
rect 5912 19552 5976 19556
rect 5992 19612 6056 19616
rect 5992 19556 5996 19612
rect 5996 19556 6052 19612
rect 6052 19556 6056 19612
rect 5992 19552 6056 19556
rect 10552 19612 10616 19616
rect 10552 19556 10556 19612
rect 10556 19556 10612 19612
rect 10612 19556 10616 19612
rect 10552 19552 10616 19556
rect 10632 19612 10696 19616
rect 10632 19556 10636 19612
rect 10636 19556 10692 19612
rect 10692 19556 10696 19612
rect 10632 19552 10696 19556
rect 10712 19612 10776 19616
rect 10712 19556 10716 19612
rect 10716 19556 10772 19612
rect 10772 19556 10776 19612
rect 10712 19552 10776 19556
rect 10792 19612 10856 19616
rect 10792 19556 10796 19612
rect 10796 19556 10852 19612
rect 10852 19556 10856 19612
rect 10792 19552 10856 19556
rect 15352 19612 15416 19616
rect 15352 19556 15356 19612
rect 15356 19556 15412 19612
rect 15412 19556 15416 19612
rect 15352 19552 15416 19556
rect 15432 19612 15496 19616
rect 15432 19556 15436 19612
rect 15436 19556 15492 19612
rect 15492 19556 15496 19612
rect 15432 19552 15496 19556
rect 15512 19612 15576 19616
rect 15512 19556 15516 19612
rect 15516 19556 15572 19612
rect 15572 19556 15576 19612
rect 15512 19552 15576 19556
rect 15592 19612 15656 19616
rect 15592 19556 15596 19612
rect 15596 19556 15652 19612
rect 15652 19556 15656 19612
rect 15592 19552 15656 19556
rect 20152 19612 20216 19616
rect 20152 19556 20156 19612
rect 20156 19556 20212 19612
rect 20212 19556 20216 19612
rect 20152 19552 20216 19556
rect 20232 19612 20296 19616
rect 20232 19556 20236 19612
rect 20236 19556 20292 19612
rect 20292 19556 20296 19612
rect 20232 19552 20296 19556
rect 20312 19612 20376 19616
rect 20312 19556 20316 19612
rect 20316 19556 20372 19612
rect 20372 19556 20376 19612
rect 20312 19552 20376 19556
rect 20392 19612 20456 19616
rect 20392 19556 20396 19612
rect 20396 19556 20452 19612
rect 20452 19556 20456 19612
rect 20392 19552 20456 19556
rect 24952 19612 25016 19616
rect 24952 19556 24956 19612
rect 24956 19556 25012 19612
rect 25012 19556 25016 19612
rect 24952 19552 25016 19556
rect 25032 19612 25096 19616
rect 25032 19556 25036 19612
rect 25036 19556 25092 19612
rect 25092 19556 25096 19612
rect 25032 19552 25096 19556
rect 25112 19612 25176 19616
rect 25112 19556 25116 19612
rect 25116 19556 25172 19612
rect 25172 19556 25176 19612
rect 25112 19552 25176 19556
rect 25192 19612 25256 19616
rect 25192 19556 25196 19612
rect 25196 19556 25252 19612
rect 25252 19556 25256 19612
rect 25192 19552 25256 19556
rect 3352 19068 3416 19072
rect 3352 19012 3356 19068
rect 3356 19012 3412 19068
rect 3412 19012 3416 19068
rect 3352 19008 3416 19012
rect 3432 19068 3496 19072
rect 3432 19012 3436 19068
rect 3436 19012 3492 19068
rect 3492 19012 3496 19068
rect 3432 19008 3496 19012
rect 3512 19068 3576 19072
rect 3512 19012 3516 19068
rect 3516 19012 3572 19068
rect 3572 19012 3576 19068
rect 3512 19008 3576 19012
rect 3592 19068 3656 19072
rect 3592 19012 3596 19068
rect 3596 19012 3652 19068
rect 3652 19012 3656 19068
rect 3592 19008 3656 19012
rect 8152 19068 8216 19072
rect 8152 19012 8156 19068
rect 8156 19012 8212 19068
rect 8212 19012 8216 19068
rect 8152 19008 8216 19012
rect 8232 19068 8296 19072
rect 8232 19012 8236 19068
rect 8236 19012 8292 19068
rect 8292 19012 8296 19068
rect 8232 19008 8296 19012
rect 8312 19068 8376 19072
rect 8312 19012 8316 19068
rect 8316 19012 8372 19068
rect 8372 19012 8376 19068
rect 8312 19008 8376 19012
rect 8392 19068 8456 19072
rect 8392 19012 8396 19068
rect 8396 19012 8452 19068
rect 8452 19012 8456 19068
rect 8392 19008 8456 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 17752 19068 17816 19072
rect 17752 19012 17756 19068
rect 17756 19012 17812 19068
rect 17812 19012 17816 19068
rect 17752 19008 17816 19012
rect 17832 19068 17896 19072
rect 17832 19012 17836 19068
rect 17836 19012 17892 19068
rect 17892 19012 17896 19068
rect 17832 19008 17896 19012
rect 17912 19068 17976 19072
rect 17912 19012 17916 19068
rect 17916 19012 17972 19068
rect 17972 19012 17976 19068
rect 17912 19008 17976 19012
rect 17992 19068 18056 19072
rect 17992 19012 17996 19068
rect 17996 19012 18052 19068
rect 18052 19012 18056 19068
rect 17992 19008 18056 19012
rect 22552 19068 22616 19072
rect 22552 19012 22556 19068
rect 22556 19012 22612 19068
rect 22612 19012 22616 19068
rect 22552 19008 22616 19012
rect 22632 19068 22696 19072
rect 22632 19012 22636 19068
rect 22636 19012 22692 19068
rect 22692 19012 22696 19068
rect 22632 19008 22696 19012
rect 22712 19068 22776 19072
rect 22712 19012 22716 19068
rect 22716 19012 22772 19068
rect 22772 19012 22776 19068
rect 22712 19008 22776 19012
rect 22792 19068 22856 19072
rect 22792 19012 22796 19068
rect 22796 19012 22852 19068
rect 22852 19012 22856 19068
rect 22792 19008 22856 19012
rect 27352 19068 27416 19072
rect 27352 19012 27356 19068
rect 27356 19012 27412 19068
rect 27412 19012 27416 19068
rect 27352 19008 27416 19012
rect 27432 19068 27496 19072
rect 27432 19012 27436 19068
rect 27436 19012 27492 19068
rect 27492 19012 27496 19068
rect 27432 19008 27496 19012
rect 27512 19068 27576 19072
rect 27512 19012 27516 19068
rect 27516 19012 27572 19068
rect 27572 19012 27576 19068
rect 27512 19008 27576 19012
rect 27592 19068 27656 19072
rect 27592 19012 27596 19068
rect 27596 19012 27652 19068
rect 27652 19012 27656 19068
rect 27592 19008 27656 19012
rect 5752 18524 5816 18528
rect 5752 18468 5756 18524
rect 5756 18468 5812 18524
rect 5812 18468 5816 18524
rect 5752 18464 5816 18468
rect 5832 18524 5896 18528
rect 5832 18468 5836 18524
rect 5836 18468 5892 18524
rect 5892 18468 5896 18524
rect 5832 18464 5896 18468
rect 5912 18524 5976 18528
rect 5912 18468 5916 18524
rect 5916 18468 5972 18524
rect 5972 18468 5976 18524
rect 5912 18464 5976 18468
rect 5992 18524 6056 18528
rect 5992 18468 5996 18524
rect 5996 18468 6052 18524
rect 6052 18468 6056 18524
rect 5992 18464 6056 18468
rect 10552 18524 10616 18528
rect 10552 18468 10556 18524
rect 10556 18468 10612 18524
rect 10612 18468 10616 18524
rect 10552 18464 10616 18468
rect 10632 18524 10696 18528
rect 10632 18468 10636 18524
rect 10636 18468 10692 18524
rect 10692 18468 10696 18524
rect 10632 18464 10696 18468
rect 10712 18524 10776 18528
rect 10712 18468 10716 18524
rect 10716 18468 10772 18524
rect 10772 18468 10776 18524
rect 10712 18464 10776 18468
rect 10792 18524 10856 18528
rect 10792 18468 10796 18524
rect 10796 18468 10852 18524
rect 10852 18468 10856 18524
rect 10792 18464 10856 18468
rect 15352 18524 15416 18528
rect 15352 18468 15356 18524
rect 15356 18468 15412 18524
rect 15412 18468 15416 18524
rect 15352 18464 15416 18468
rect 15432 18524 15496 18528
rect 15432 18468 15436 18524
rect 15436 18468 15492 18524
rect 15492 18468 15496 18524
rect 15432 18464 15496 18468
rect 15512 18524 15576 18528
rect 15512 18468 15516 18524
rect 15516 18468 15572 18524
rect 15572 18468 15576 18524
rect 15512 18464 15576 18468
rect 15592 18524 15656 18528
rect 15592 18468 15596 18524
rect 15596 18468 15652 18524
rect 15652 18468 15656 18524
rect 15592 18464 15656 18468
rect 20152 18524 20216 18528
rect 20152 18468 20156 18524
rect 20156 18468 20212 18524
rect 20212 18468 20216 18524
rect 20152 18464 20216 18468
rect 20232 18524 20296 18528
rect 20232 18468 20236 18524
rect 20236 18468 20292 18524
rect 20292 18468 20296 18524
rect 20232 18464 20296 18468
rect 20312 18524 20376 18528
rect 20312 18468 20316 18524
rect 20316 18468 20372 18524
rect 20372 18468 20376 18524
rect 20312 18464 20376 18468
rect 20392 18524 20456 18528
rect 20392 18468 20396 18524
rect 20396 18468 20452 18524
rect 20452 18468 20456 18524
rect 20392 18464 20456 18468
rect 24952 18524 25016 18528
rect 24952 18468 24956 18524
rect 24956 18468 25012 18524
rect 25012 18468 25016 18524
rect 24952 18464 25016 18468
rect 25032 18524 25096 18528
rect 25032 18468 25036 18524
rect 25036 18468 25092 18524
rect 25092 18468 25096 18524
rect 25032 18464 25096 18468
rect 25112 18524 25176 18528
rect 25112 18468 25116 18524
rect 25116 18468 25172 18524
rect 25172 18468 25176 18524
rect 25112 18464 25176 18468
rect 25192 18524 25256 18528
rect 25192 18468 25196 18524
rect 25196 18468 25252 18524
rect 25252 18468 25256 18524
rect 25192 18464 25256 18468
rect 3352 17980 3416 17984
rect 3352 17924 3356 17980
rect 3356 17924 3412 17980
rect 3412 17924 3416 17980
rect 3352 17920 3416 17924
rect 3432 17980 3496 17984
rect 3432 17924 3436 17980
rect 3436 17924 3492 17980
rect 3492 17924 3496 17980
rect 3432 17920 3496 17924
rect 3512 17980 3576 17984
rect 3512 17924 3516 17980
rect 3516 17924 3572 17980
rect 3572 17924 3576 17980
rect 3512 17920 3576 17924
rect 3592 17980 3656 17984
rect 3592 17924 3596 17980
rect 3596 17924 3652 17980
rect 3652 17924 3656 17980
rect 3592 17920 3656 17924
rect 8152 17980 8216 17984
rect 8152 17924 8156 17980
rect 8156 17924 8212 17980
rect 8212 17924 8216 17980
rect 8152 17920 8216 17924
rect 8232 17980 8296 17984
rect 8232 17924 8236 17980
rect 8236 17924 8292 17980
rect 8292 17924 8296 17980
rect 8232 17920 8296 17924
rect 8312 17980 8376 17984
rect 8312 17924 8316 17980
rect 8316 17924 8372 17980
rect 8372 17924 8376 17980
rect 8312 17920 8376 17924
rect 8392 17980 8456 17984
rect 8392 17924 8396 17980
rect 8396 17924 8452 17980
rect 8452 17924 8456 17980
rect 8392 17920 8456 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 17752 17980 17816 17984
rect 17752 17924 17756 17980
rect 17756 17924 17812 17980
rect 17812 17924 17816 17980
rect 17752 17920 17816 17924
rect 17832 17980 17896 17984
rect 17832 17924 17836 17980
rect 17836 17924 17892 17980
rect 17892 17924 17896 17980
rect 17832 17920 17896 17924
rect 17912 17980 17976 17984
rect 17912 17924 17916 17980
rect 17916 17924 17972 17980
rect 17972 17924 17976 17980
rect 17912 17920 17976 17924
rect 17992 17980 18056 17984
rect 17992 17924 17996 17980
rect 17996 17924 18052 17980
rect 18052 17924 18056 17980
rect 17992 17920 18056 17924
rect 22552 17980 22616 17984
rect 22552 17924 22556 17980
rect 22556 17924 22612 17980
rect 22612 17924 22616 17980
rect 22552 17920 22616 17924
rect 22632 17980 22696 17984
rect 22632 17924 22636 17980
rect 22636 17924 22692 17980
rect 22692 17924 22696 17980
rect 22632 17920 22696 17924
rect 22712 17980 22776 17984
rect 22712 17924 22716 17980
rect 22716 17924 22772 17980
rect 22772 17924 22776 17980
rect 22712 17920 22776 17924
rect 22792 17980 22856 17984
rect 22792 17924 22796 17980
rect 22796 17924 22852 17980
rect 22852 17924 22856 17980
rect 22792 17920 22856 17924
rect 27352 17980 27416 17984
rect 27352 17924 27356 17980
rect 27356 17924 27412 17980
rect 27412 17924 27416 17980
rect 27352 17920 27416 17924
rect 27432 17980 27496 17984
rect 27432 17924 27436 17980
rect 27436 17924 27492 17980
rect 27492 17924 27496 17980
rect 27432 17920 27496 17924
rect 27512 17980 27576 17984
rect 27512 17924 27516 17980
rect 27516 17924 27572 17980
rect 27572 17924 27576 17980
rect 27512 17920 27576 17924
rect 27592 17980 27656 17984
rect 27592 17924 27596 17980
rect 27596 17924 27652 17980
rect 27652 17924 27656 17980
rect 27592 17920 27656 17924
rect 5752 17436 5816 17440
rect 5752 17380 5756 17436
rect 5756 17380 5812 17436
rect 5812 17380 5816 17436
rect 5752 17376 5816 17380
rect 5832 17436 5896 17440
rect 5832 17380 5836 17436
rect 5836 17380 5892 17436
rect 5892 17380 5896 17436
rect 5832 17376 5896 17380
rect 5912 17436 5976 17440
rect 5912 17380 5916 17436
rect 5916 17380 5972 17436
rect 5972 17380 5976 17436
rect 5912 17376 5976 17380
rect 5992 17436 6056 17440
rect 5992 17380 5996 17436
rect 5996 17380 6052 17436
rect 6052 17380 6056 17436
rect 5992 17376 6056 17380
rect 10552 17436 10616 17440
rect 10552 17380 10556 17436
rect 10556 17380 10612 17436
rect 10612 17380 10616 17436
rect 10552 17376 10616 17380
rect 10632 17436 10696 17440
rect 10632 17380 10636 17436
rect 10636 17380 10692 17436
rect 10692 17380 10696 17436
rect 10632 17376 10696 17380
rect 10712 17436 10776 17440
rect 10712 17380 10716 17436
rect 10716 17380 10772 17436
rect 10772 17380 10776 17436
rect 10712 17376 10776 17380
rect 10792 17436 10856 17440
rect 10792 17380 10796 17436
rect 10796 17380 10852 17436
rect 10852 17380 10856 17436
rect 10792 17376 10856 17380
rect 15352 17436 15416 17440
rect 15352 17380 15356 17436
rect 15356 17380 15412 17436
rect 15412 17380 15416 17436
rect 15352 17376 15416 17380
rect 15432 17436 15496 17440
rect 15432 17380 15436 17436
rect 15436 17380 15492 17436
rect 15492 17380 15496 17436
rect 15432 17376 15496 17380
rect 15512 17436 15576 17440
rect 15512 17380 15516 17436
rect 15516 17380 15572 17436
rect 15572 17380 15576 17436
rect 15512 17376 15576 17380
rect 15592 17436 15656 17440
rect 15592 17380 15596 17436
rect 15596 17380 15652 17436
rect 15652 17380 15656 17436
rect 15592 17376 15656 17380
rect 20152 17436 20216 17440
rect 20152 17380 20156 17436
rect 20156 17380 20212 17436
rect 20212 17380 20216 17436
rect 20152 17376 20216 17380
rect 20232 17436 20296 17440
rect 20232 17380 20236 17436
rect 20236 17380 20292 17436
rect 20292 17380 20296 17436
rect 20232 17376 20296 17380
rect 20312 17436 20376 17440
rect 20312 17380 20316 17436
rect 20316 17380 20372 17436
rect 20372 17380 20376 17436
rect 20312 17376 20376 17380
rect 20392 17436 20456 17440
rect 20392 17380 20396 17436
rect 20396 17380 20452 17436
rect 20452 17380 20456 17436
rect 20392 17376 20456 17380
rect 24952 17436 25016 17440
rect 24952 17380 24956 17436
rect 24956 17380 25012 17436
rect 25012 17380 25016 17436
rect 24952 17376 25016 17380
rect 25032 17436 25096 17440
rect 25032 17380 25036 17436
rect 25036 17380 25092 17436
rect 25092 17380 25096 17436
rect 25032 17376 25096 17380
rect 25112 17436 25176 17440
rect 25112 17380 25116 17436
rect 25116 17380 25172 17436
rect 25172 17380 25176 17436
rect 25112 17376 25176 17380
rect 25192 17436 25256 17440
rect 25192 17380 25196 17436
rect 25196 17380 25252 17436
rect 25252 17380 25256 17436
rect 25192 17376 25256 17380
rect 3352 16892 3416 16896
rect 3352 16836 3356 16892
rect 3356 16836 3412 16892
rect 3412 16836 3416 16892
rect 3352 16832 3416 16836
rect 3432 16892 3496 16896
rect 3432 16836 3436 16892
rect 3436 16836 3492 16892
rect 3492 16836 3496 16892
rect 3432 16832 3496 16836
rect 3512 16892 3576 16896
rect 3512 16836 3516 16892
rect 3516 16836 3572 16892
rect 3572 16836 3576 16892
rect 3512 16832 3576 16836
rect 3592 16892 3656 16896
rect 3592 16836 3596 16892
rect 3596 16836 3652 16892
rect 3652 16836 3656 16892
rect 3592 16832 3656 16836
rect 8152 16892 8216 16896
rect 8152 16836 8156 16892
rect 8156 16836 8212 16892
rect 8212 16836 8216 16892
rect 8152 16832 8216 16836
rect 8232 16892 8296 16896
rect 8232 16836 8236 16892
rect 8236 16836 8292 16892
rect 8292 16836 8296 16892
rect 8232 16832 8296 16836
rect 8312 16892 8376 16896
rect 8312 16836 8316 16892
rect 8316 16836 8372 16892
rect 8372 16836 8376 16892
rect 8312 16832 8376 16836
rect 8392 16892 8456 16896
rect 8392 16836 8396 16892
rect 8396 16836 8452 16892
rect 8452 16836 8456 16892
rect 8392 16832 8456 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 17752 16892 17816 16896
rect 17752 16836 17756 16892
rect 17756 16836 17812 16892
rect 17812 16836 17816 16892
rect 17752 16832 17816 16836
rect 17832 16892 17896 16896
rect 17832 16836 17836 16892
rect 17836 16836 17892 16892
rect 17892 16836 17896 16892
rect 17832 16832 17896 16836
rect 17912 16892 17976 16896
rect 17912 16836 17916 16892
rect 17916 16836 17972 16892
rect 17972 16836 17976 16892
rect 17912 16832 17976 16836
rect 17992 16892 18056 16896
rect 17992 16836 17996 16892
rect 17996 16836 18052 16892
rect 18052 16836 18056 16892
rect 17992 16832 18056 16836
rect 22552 16892 22616 16896
rect 22552 16836 22556 16892
rect 22556 16836 22612 16892
rect 22612 16836 22616 16892
rect 22552 16832 22616 16836
rect 22632 16892 22696 16896
rect 22632 16836 22636 16892
rect 22636 16836 22692 16892
rect 22692 16836 22696 16892
rect 22632 16832 22696 16836
rect 22712 16892 22776 16896
rect 22712 16836 22716 16892
rect 22716 16836 22772 16892
rect 22772 16836 22776 16892
rect 22712 16832 22776 16836
rect 22792 16892 22856 16896
rect 22792 16836 22796 16892
rect 22796 16836 22852 16892
rect 22852 16836 22856 16892
rect 22792 16832 22856 16836
rect 27352 16892 27416 16896
rect 27352 16836 27356 16892
rect 27356 16836 27412 16892
rect 27412 16836 27416 16892
rect 27352 16832 27416 16836
rect 27432 16892 27496 16896
rect 27432 16836 27436 16892
rect 27436 16836 27492 16892
rect 27492 16836 27496 16892
rect 27432 16832 27496 16836
rect 27512 16892 27576 16896
rect 27512 16836 27516 16892
rect 27516 16836 27572 16892
rect 27572 16836 27576 16892
rect 27512 16832 27576 16836
rect 27592 16892 27656 16896
rect 27592 16836 27596 16892
rect 27596 16836 27652 16892
rect 27652 16836 27656 16892
rect 27592 16832 27656 16836
rect 5752 16348 5816 16352
rect 5752 16292 5756 16348
rect 5756 16292 5812 16348
rect 5812 16292 5816 16348
rect 5752 16288 5816 16292
rect 5832 16348 5896 16352
rect 5832 16292 5836 16348
rect 5836 16292 5892 16348
rect 5892 16292 5896 16348
rect 5832 16288 5896 16292
rect 5912 16348 5976 16352
rect 5912 16292 5916 16348
rect 5916 16292 5972 16348
rect 5972 16292 5976 16348
rect 5912 16288 5976 16292
rect 5992 16348 6056 16352
rect 5992 16292 5996 16348
rect 5996 16292 6052 16348
rect 6052 16292 6056 16348
rect 5992 16288 6056 16292
rect 10552 16348 10616 16352
rect 10552 16292 10556 16348
rect 10556 16292 10612 16348
rect 10612 16292 10616 16348
rect 10552 16288 10616 16292
rect 10632 16348 10696 16352
rect 10632 16292 10636 16348
rect 10636 16292 10692 16348
rect 10692 16292 10696 16348
rect 10632 16288 10696 16292
rect 10712 16348 10776 16352
rect 10712 16292 10716 16348
rect 10716 16292 10772 16348
rect 10772 16292 10776 16348
rect 10712 16288 10776 16292
rect 10792 16348 10856 16352
rect 10792 16292 10796 16348
rect 10796 16292 10852 16348
rect 10852 16292 10856 16348
rect 10792 16288 10856 16292
rect 15352 16348 15416 16352
rect 15352 16292 15356 16348
rect 15356 16292 15412 16348
rect 15412 16292 15416 16348
rect 15352 16288 15416 16292
rect 15432 16348 15496 16352
rect 15432 16292 15436 16348
rect 15436 16292 15492 16348
rect 15492 16292 15496 16348
rect 15432 16288 15496 16292
rect 15512 16348 15576 16352
rect 15512 16292 15516 16348
rect 15516 16292 15572 16348
rect 15572 16292 15576 16348
rect 15512 16288 15576 16292
rect 15592 16348 15656 16352
rect 15592 16292 15596 16348
rect 15596 16292 15652 16348
rect 15652 16292 15656 16348
rect 15592 16288 15656 16292
rect 20152 16348 20216 16352
rect 20152 16292 20156 16348
rect 20156 16292 20212 16348
rect 20212 16292 20216 16348
rect 20152 16288 20216 16292
rect 20232 16348 20296 16352
rect 20232 16292 20236 16348
rect 20236 16292 20292 16348
rect 20292 16292 20296 16348
rect 20232 16288 20296 16292
rect 20312 16348 20376 16352
rect 20312 16292 20316 16348
rect 20316 16292 20372 16348
rect 20372 16292 20376 16348
rect 20312 16288 20376 16292
rect 20392 16348 20456 16352
rect 20392 16292 20396 16348
rect 20396 16292 20452 16348
rect 20452 16292 20456 16348
rect 20392 16288 20456 16292
rect 24952 16348 25016 16352
rect 24952 16292 24956 16348
rect 24956 16292 25012 16348
rect 25012 16292 25016 16348
rect 24952 16288 25016 16292
rect 25032 16348 25096 16352
rect 25032 16292 25036 16348
rect 25036 16292 25092 16348
rect 25092 16292 25096 16348
rect 25032 16288 25096 16292
rect 25112 16348 25176 16352
rect 25112 16292 25116 16348
rect 25116 16292 25172 16348
rect 25172 16292 25176 16348
rect 25112 16288 25176 16292
rect 25192 16348 25256 16352
rect 25192 16292 25196 16348
rect 25196 16292 25252 16348
rect 25252 16292 25256 16348
rect 25192 16288 25256 16292
rect 3352 15804 3416 15808
rect 3352 15748 3356 15804
rect 3356 15748 3412 15804
rect 3412 15748 3416 15804
rect 3352 15744 3416 15748
rect 3432 15804 3496 15808
rect 3432 15748 3436 15804
rect 3436 15748 3492 15804
rect 3492 15748 3496 15804
rect 3432 15744 3496 15748
rect 3512 15804 3576 15808
rect 3512 15748 3516 15804
rect 3516 15748 3572 15804
rect 3572 15748 3576 15804
rect 3512 15744 3576 15748
rect 3592 15804 3656 15808
rect 3592 15748 3596 15804
rect 3596 15748 3652 15804
rect 3652 15748 3656 15804
rect 3592 15744 3656 15748
rect 8152 15804 8216 15808
rect 8152 15748 8156 15804
rect 8156 15748 8212 15804
rect 8212 15748 8216 15804
rect 8152 15744 8216 15748
rect 8232 15804 8296 15808
rect 8232 15748 8236 15804
rect 8236 15748 8292 15804
rect 8292 15748 8296 15804
rect 8232 15744 8296 15748
rect 8312 15804 8376 15808
rect 8312 15748 8316 15804
rect 8316 15748 8372 15804
rect 8372 15748 8376 15804
rect 8312 15744 8376 15748
rect 8392 15804 8456 15808
rect 8392 15748 8396 15804
rect 8396 15748 8452 15804
rect 8452 15748 8456 15804
rect 8392 15744 8456 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 17752 15804 17816 15808
rect 17752 15748 17756 15804
rect 17756 15748 17812 15804
rect 17812 15748 17816 15804
rect 17752 15744 17816 15748
rect 17832 15804 17896 15808
rect 17832 15748 17836 15804
rect 17836 15748 17892 15804
rect 17892 15748 17896 15804
rect 17832 15744 17896 15748
rect 17912 15804 17976 15808
rect 17912 15748 17916 15804
rect 17916 15748 17972 15804
rect 17972 15748 17976 15804
rect 17912 15744 17976 15748
rect 17992 15804 18056 15808
rect 17992 15748 17996 15804
rect 17996 15748 18052 15804
rect 18052 15748 18056 15804
rect 17992 15744 18056 15748
rect 22552 15804 22616 15808
rect 22552 15748 22556 15804
rect 22556 15748 22612 15804
rect 22612 15748 22616 15804
rect 22552 15744 22616 15748
rect 22632 15804 22696 15808
rect 22632 15748 22636 15804
rect 22636 15748 22692 15804
rect 22692 15748 22696 15804
rect 22632 15744 22696 15748
rect 22712 15804 22776 15808
rect 22712 15748 22716 15804
rect 22716 15748 22772 15804
rect 22772 15748 22776 15804
rect 22712 15744 22776 15748
rect 22792 15804 22856 15808
rect 22792 15748 22796 15804
rect 22796 15748 22852 15804
rect 22852 15748 22856 15804
rect 22792 15744 22856 15748
rect 27352 15804 27416 15808
rect 27352 15748 27356 15804
rect 27356 15748 27412 15804
rect 27412 15748 27416 15804
rect 27352 15744 27416 15748
rect 27432 15804 27496 15808
rect 27432 15748 27436 15804
rect 27436 15748 27492 15804
rect 27492 15748 27496 15804
rect 27432 15744 27496 15748
rect 27512 15804 27576 15808
rect 27512 15748 27516 15804
rect 27516 15748 27572 15804
rect 27572 15748 27576 15804
rect 27512 15744 27576 15748
rect 27592 15804 27656 15808
rect 27592 15748 27596 15804
rect 27596 15748 27652 15804
rect 27652 15748 27656 15804
rect 27592 15744 27656 15748
rect 5752 15260 5816 15264
rect 5752 15204 5756 15260
rect 5756 15204 5812 15260
rect 5812 15204 5816 15260
rect 5752 15200 5816 15204
rect 5832 15260 5896 15264
rect 5832 15204 5836 15260
rect 5836 15204 5892 15260
rect 5892 15204 5896 15260
rect 5832 15200 5896 15204
rect 5912 15260 5976 15264
rect 5912 15204 5916 15260
rect 5916 15204 5972 15260
rect 5972 15204 5976 15260
rect 5912 15200 5976 15204
rect 5992 15260 6056 15264
rect 5992 15204 5996 15260
rect 5996 15204 6052 15260
rect 6052 15204 6056 15260
rect 5992 15200 6056 15204
rect 10552 15260 10616 15264
rect 10552 15204 10556 15260
rect 10556 15204 10612 15260
rect 10612 15204 10616 15260
rect 10552 15200 10616 15204
rect 10632 15260 10696 15264
rect 10632 15204 10636 15260
rect 10636 15204 10692 15260
rect 10692 15204 10696 15260
rect 10632 15200 10696 15204
rect 10712 15260 10776 15264
rect 10712 15204 10716 15260
rect 10716 15204 10772 15260
rect 10772 15204 10776 15260
rect 10712 15200 10776 15204
rect 10792 15260 10856 15264
rect 10792 15204 10796 15260
rect 10796 15204 10852 15260
rect 10852 15204 10856 15260
rect 10792 15200 10856 15204
rect 15352 15260 15416 15264
rect 15352 15204 15356 15260
rect 15356 15204 15412 15260
rect 15412 15204 15416 15260
rect 15352 15200 15416 15204
rect 15432 15260 15496 15264
rect 15432 15204 15436 15260
rect 15436 15204 15492 15260
rect 15492 15204 15496 15260
rect 15432 15200 15496 15204
rect 15512 15260 15576 15264
rect 15512 15204 15516 15260
rect 15516 15204 15572 15260
rect 15572 15204 15576 15260
rect 15512 15200 15576 15204
rect 15592 15260 15656 15264
rect 15592 15204 15596 15260
rect 15596 15204 15652 15260
rect 15652 15204 15656 15260
rect 15592 15200 15656 15204
rect 20152 15260 20216 15264
rect 20152 15204 20156 15260
rect 20156 15204 20212 15260
rect 20212 15204 20216 15260
rect 20152 15200 20216 15204
rect 20232 15260 20296 15264
rect 20232 15204 20236 15260
rect 20236 15204 20292 15260
rect 20292 15204 20296 15260
rect 20232 15200 20296 15204
rect 20312 15260 20376 15264
rect 20312 15204 20316 15260
rect 20316 15204 20372 15260
rect 20372 15204 20376 15260
rect 20312 15200 20376 15204
rect 20392 15260 20456 15264
rect 20392 15204 20396 15260
rect 20396 15204 20452 15260
rect 20452 15204 20456 15260
rect 20392 15200 20456 15204
rect 24952 15260 25016 15264
rect 24952 15204 24956 15260
rect 24956 15204 25012 15260
rect 25012 15204 25016 15260
rect 24952 15200 25016 15204
rect 25032 15260 25096 15264
rect 25032 15204 25036 15260
rect 25036 15204 25092 15260
rect 25092 15204 25096 15260
rect 25032 15200 25096 15204
rect 25112 15260 25176 15264
rect 25112 15204 25116 15260
rect 25116 15204 25172 15260
rect 25172 15204 25176 15260
rect 25112 15200 25176 15204
rect 25192 15260 25256 15264
rect 25192 15204 25196 15260
rect 25196 15204 25252 15260
rect 25252 15204 25256 15260
rect 25192 15200 25256 15204
rect 3352 14716 3416 14720
rect 3352 14660 3356 14716
rect 3356 14660 3412 14716
rect 3412 14660 3416 14716
rect 3352 14656 3416 14660
rect 3432 14716 3496 14720
rect 3432 14660 3436 14716
rect 3436 14660 3492 14716
rect 3492 14660 3496 14716
rect 3432 14656 3496 14660
rect 3512 14716 3576 14720
rect 3512 14660 3516 14716
rect 3516 14660 3572 14716
rect 3572 14660 3576 14716
rect 3512 14656 3576 14660
rect 3592 14716 3656 14720
rect 3592 14660 3596 14716
rect 3596 14660 3652 14716
rect 3652 14660 3656 14716
rect 3592 14656 3656 14660
rect 8152 14716 8216 14720
rect 8152 14660 8156 14716
rect 8156 14660 8212 14716
rect 8212 14660 8216 14716
rect 8152 14656 8216 14660
rect 8232 14716 8296 14720
rect 8232 14660 8236 14716
rect 8236 14660 8292 14716
rect 8292 14660 8296 14716
rect 8232 14656 8296 14660
rect 8312 14716 8376 14720
rect 8312 14660 8316 14716
rect 8316 14660 8372 14716
rect 8372 14660 8376 14716
rect 8312 14656 8376 14660
rect 8392 14716 8456 14720
rect 8392 14660 8396 14716
rect 8396 14660 8452 14716
rect 8452 14660 8456 14716
rect 8392 14656 8456 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 17752 14716 17816 14720
rect 17752 14660 17756 14716
rect 17756 14660 17812 14716
rect 17812 14660 17816 14716
rect 17752 14656 17816 14660
rect 17832 14716 17896 14720
rect 17832 14660 17836 14716
rect 17836 14660 17892 14716
rect 17892 14660 17896 14716
rect 17832 14656 17896 14660
rect 17912 14716 17976 14720
rect 17912 14660 17916 14716
rect 17916 14660 17972 14716
rect 17972 14660 17976 14716
rect 17912 14656 17976 14660
rect 17992 14716 18056 14720
rect 17992 14660 17996 14716
rect 17996 14660 18052 14716
rect 18052 14660 18056 14716
rect 17992 14656 18056 14660
rect 22552 14716 22616 14720
rect 22552 14660 22556 14716
rect 22556 14660 22612 14716
rect 22612 14660 22616 14716
rect 22552 14656 22616 14660
rect 22632 14716 22696 14720
rect 22632 14660 22636 14716
rect 22636 14660 22692 14716
rect 22692 14660 22696 14716
rect 22632 14656 22696 14660
rect 22712 14716 22776 14720
rect 22712 14660 22716 14716
rect 22716 14660 22772 14716
rect 22772 14660 22776 14716
rect 22712 14656 22776 14660
rect 22792 14716 22856 14720
rect 22792 14660 22796 14716
rect 22796 14660 22852 14716
rect 22852 14660 22856 14716
rect 22792 14656 22856 14660
rect 27352 14716 27416 14720
rect 27352 14660 27356 14716
rect 27356 14660 27412 14716
rect 27412 14660 27416 14716
rect 27352 14656 27416 14660
rect 27432 14716 27496 14720
rect 27432 14660 27436 14716
rect 27436 14660 27492 14716
rect 27492 14660 27496 14716
rect 27432 14656 27496 14660
rect 27512 14716 27576 14720
rect 27512 14660 27516 14716
rect 27516 14660 27572 14716
rect 27572 14660 27576 14716
rect 27512 14656 27576 14660
rect 27592 14716 27656 14720
rect 27592 14660 27596 14716
rect 27596 14660 27652 14716
rect 27652 14660 27656 14716
rect 27592 14656 27656 14660
rect 5752 14172 5816 14176
rect 5752 14116 5756 14172
rect 5756 14116 5812 14172
rect 5812 14116 5816 14172
rect 5752 14112 5816 14116
rect 5832 14172 5896 14176
rect 5832 14116 5836 14172
rect 5836 14116 5892 14172
rect 5892 14116 5896 14172
rect 5832 14112 5896 14116
rect 5912 14172 5976 14176
rect 5912 14116 5916 14172
rect 5916 14116 5972 14172
rect 5972 14116 5976 14172
rect 5912 14112 5976 14116
rect 5992 14172 6056 14176
rect 5992 14116 5996 14172
rect 5996 14116 6052 14172
rect 6052 14116 6056 14172
rect 5992 14112 6056 14116
rect 10552 14172 10616 14176
rect 10552 14116 10556 14172
rect 10556 14116 10612 14172
rect 10612 14116 10616 14172
rect 10552 14112 10616 14116
rect 10632 14172 10696 14176
rect 10632 14116 10636 14172
rect 10636 14116 10692 14172
rect 10692 14116 10696 14172
rect 10632 14112 10696 14116
rect 10712 14172 10776 14176
rect 10712 14116 10716 14172
rect 10716 14116 10772 14172
rect 10772 14116 10776 14172
rect 10712 14112 10776 14116
rect 10792 14172 10856 14176
rect 10792 14116 10796 14172
rect 10796 14116 10852 14172
rect 10852 14116 10856 14172
rect 10792 14112 10856 14116
rect 15352 14172 15416 14176
rect 15352 14116 15356 14172
rect 15356 14116 15412 14172
rect 15412 14116 15416 14172
rect 15352 14112 15416 14116
rect 15432 14172 15496 14176
rect 15432 14116 15436 14172
rect 15436 14116 15492 14172
rect 15492 14116 15496 14172
rect 15432 14112 15496 14116
rect 15512 14172 15576 14176
rect 15512 14116 15516 14172
rect 15516 14116 15572 14172
rect 15572 14116 15576 14172
rect 15512 14112 15576 14116
rect 15592 14172 15656 14176
rect 15592 14116 15596 14172
rect 15596 14116 15652 14172
rect 15652 14116 15656 14172
rect 15592 14112 15656 14116
rect 20152 14172 20216 14176
rect 20152 14116 20156 14172
rect 20156 14116 20212 14172
rect 20212 14116 20216 14172
rect 20152 14112 20216 14116
rect 20232 14172 20296 14176
rect 20232 14116 20236 14172
rect 20236 14116 20292 14172
rect 20292 14116 20296 14172
rect 20232 14112 20296 14116
rect 20312 14172 20376 14176
rect 20312 14116 20316 14172
rect 20316 14116 20372 14172
rect 20372 14116 20376 14172
rect 20312 14112 20376 14116
rect 20392 14172 20456 14176
rect 20392 14116 20396 14172
rect 20396 14116 20452 14172
rect 20452 14116 20456 14172
rect 20392 14112 20456 14116
rect 24952 14172 25016 14176
rect 24952 14116 24956 14172
rect 24956 14116 25012 14172
rect 25012 14116 25016 14172
rect 24952 14112 25016 14116
rect 25032 14172 25096 14176
rect 25032 14116 25036 14172
rect 25036 14116 25092 14172
rect 25092 14116 25096 14172
rect 25032 14112 25096 14116
rect 25112 14172 25176 14176
rect 25112 14116 25116 14172
rect 25116 14116 25172 14172
rect 25172 14116 25176 14172
rect 25112 14112 25176 14116
rect 25192 14172 25256 14176
rect 25192 14116 25196 14172
rect 25196 14116 25252 14172
rect 25252 14116 25256 14172
rect 25192 14112 25256 14116
rect 3352 13628 3416 13632
rect 3352 13572 3356 13628
rect 3356 13572 3412 13628
rect 3412 13572 3416 13628
rect 3352 13568 3416 13572
rect 3432 13628 3496 13632
rect 3432 13572 3436 13628
rect 3436 13572 3492 13628
rect 3492 13572 3496 13628
rect 3432 13568 3496 13572
rect 3512 13628 3576 13632
rect 3512 13572 3516 13628
rect 3516 13572 3572 13628
rect 3572 13572 3576 13628
rect 3512 13568 3576 13572
rect 3592 13628 3656 13632
rect 3592 13572 3596 13628
rect 3596 13572 3652 13628
rect 3652 13572 3656 13628
rect 3592 13568 3656 13572
rect 8152 13628 8216 13632
rect 8152 13572 8156 13628
rect 8156 13572 8212 13628
rect 8212 13572 8216 13628
rect 8152 13568 8216 13572
rect 8232 13628 8296 13632
rect 8232 13572 8236 13628
rect 8236 13572 8292 13628
rect 8292 13572 8296 13628
rect 8232 13568 8296 13572
rect 8312 13628 8376 13632
rect 8312 13572 8316 13628
rect 8316 13572 8372 13628
rect 8372 13572 8376 13628
rect 8312 13568 8376 13572
rect 8392 13628 8456 13632
rect 8392 13572 8396 13628
rect 8396 13572 8452 13628
rect 8452 13572 8456 13628
rect 8392 13568 8456 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 17752 13628 17816 13632
rect 17752 13572 17756 13628
rect 17756 13572 17812 13628
rect 17812 13572 17816 13628
rect 17752 13568 17816 13572
rect 17832 13628 17896 13632
rect 17832 13572 17836 13628
rect 17836 13572 17892 13628
rect 17892 13572 17896 13628
rect 17832 13568 17896 13572
rect 17912 13628 17976 13632
rect 17912 13572 17916 13628
rect 17916 13572 17972 13628
rect 17972 13572 17976 13628
rect 17912 13568 17976 13572
rect 17992 13628 18056 13632
rect 17992 13572 17996 13628
rect 17996 13572 18052 13628
rect 18052 13572 18056 13628
rect 17992 13568 18056 13572
rect 22552 13628 22616 13632
rect 22552 13572 22556 13628
rect 22556 13572 22612 13628
rect 22612 13572 22616 13628
rect 22552 13568 22616 13572
rect 22632 13628 22696 13632
rect 22632 13572 22636 13628
rect 22636 13572 22692 13628
rect 22692 13572 22696 13628
rect 22632 13568 22696 13572
rect 22712 13628 22776 13632
rect 22712 13572 22716 13628
rect 22716 13572 22772 13628
rect 22772 13572 22776 13628
rect 22712 13568 22776 13572
rect 22792 13628 22856 13632
rect 22792 13572 22796 13628
rect 22796 13572 22852 13628
rect 22852 13572 22856 13628
rect 22792 13568 22856 13572
rect 27352 13628 27416 13632
rect 27352 13572 27356 13628
rect 27356 13572 27412 13628
rect 27412 13572 27416 13628
rect 27352 13568 27416 13572
rect 27432 13628 27496 13632
rect 27432 13572 27436 13628
rect 27436 13572 27492 13628
rect 27492 13572 27496 13628
rect 27432 13568 27496 13572
rect 27512 13628 27576 13632
rect 27512 13572 27516 13628
rect 27516 13572 27572 13628
rect 27572 13572 27576 13628
rect 27512 13568 27576 13572
rect 27592 13628 27656 13632
rect 27592 13572 27596 13628
rect 27596 13572 27652 13628
rect 27652 13572 27656 13628
rect 27592 13568 27656 13572
rect 5752 13084 5816 13088
rect 5752 13028 5756 13084
rect 5756 13028 5812 13084
rect 5812 13028 5816 13084
rect 5752 13024 5816 13028
rect 5832 13084 5896 13088
rect 5832 13028 5836 13084
rect 5836 13028 5892 13084
rect 5892 13028 5896 13084
rect 5832 13024 5896 13028
rect 5912 13084 5976 13088
rect 5912 13028 5916 13084
rect 5916 13028 5972 13084
rect 5972 13028 5976 13084
rect 5912 13024 5976 13028
rect 5992 13084 6056 13088
rect 5992 13028 5996 13084
rect 5996 13028 6052 13084
rect 6052 13028 6056 13084
rect 5992 13024 6056 13028
rect 10552 13084 10616 13088
rect 10552 13028 10556 13084
rect 10556 13028 10612 13084
rect 10612 13028 10616 13084
rect 10552 13024 10616 13028
rect 10632 13084 10696 13088
rect 10632 13028 10636 13084
rect 10636 13028 10692 13084
rect 10692 13028 10696 13084
rect 10632 13024 10696 13028
rect 10712 13084 10776 13088
rect 10712 13028 10716 13084
rect 10716 13028 10772 13084
rect 10772 13028 10776 13084
rect 10712 13024 10776 13028
rect 10792 13084 10856 13088
rect 10792 13028 10796 13084
rect 10796 13028 10852 13084
rect 10852 13028 10856 13084
rect 10792 13024 10856 13028
rect 15352 13084 15416 13088
rect 15352 13028 15356 13084
rect 15356 13028 15412 13084
rect 15412 13028 15416 13084
rect 15352 13024 15416 13028
rect 15432 13084 15496 13088
rect 15432 13028 15436 13084
rect 15436 13028 15492 13084
rect 15492 13028 15496 13084
rect 15432 13024 15496 13028
rect 15512 13084 15576 13088
rect 15512 13028 15516 13084
rect 15516 13028 15572 13084
rect 15572 13028 15576 13084
rect 15512 13024 15576 13028
rect 15592 13084 15656 13088
rect 15592 13028 15596 13084
rect 15596 13028 15652 13084
rect 15652 13028 15656 13084
rect 15592 13024 15656 13028
rect 20152 13084 20216 13088
rect 20152 13028 20156 13084
rect 20156 13028 20212 13084
rect 20212 13028 20216 13084
rect 20152 13024 20216 13028
rect 20232 13084 20296 13088
rect 20232 13028 20236 13084
rect 20236 13028 20292 13084
rect 20292 13028 20296 13084
rect 20232 13024 20296 13028
rect 20312 13084 20376 13088
rect 20312 13028 20316 13084
rect 20316 13028 20372 13084
rect 20372 13028 20376 13084
rect 20312 13024 20376 13028
rect 20392 13084 20456 13088
rect 20392 13028 20396 13084
rect 20396 13028 20452 13084
rect 20452 13028 20456 13084
rect 20392 13024 20456 13028
rect 24952 13084 25016 13088
rect 24952 13028 24956 13084
rect 24956 13028 25012 13084
rect 25012 13028 25016 13084
rect 24952 13024 25016 13028
rect 25032 13084 25096 13088
rect 25032 13028 25036 13084
rect 25036 13028 25092 13084
rect 25092 13028 25096 13084
rect 25032 13024 25096 13028
rect 25112 13084 25176 13088
rect 25112 13028 25116 13084
rect 25116 13028 25172 13084
rect 25172 13028 25176 13084
rect 25112 13024 25176 13028
rect 25192 13084 25256 13088
rect 25192 13028 25196 13084
rect 25196 13028 25252 13084
rect 25252 13028 25256 13084
rect 25192 13024 25256 13028
rect 3352 12540 3416 12544
rect 3352 12484 3356 12540
rect 3356 12484 3412 12540
rect 3412 12484 3416 12540
rect 3352 12480 3416 12484
rect 3432 12540 3496 12544
rect 3432 12484 3436 12540
rect 3436 12484 3492 12540
rect 3492 12484 3496 12540
rect 3432 12480 3496 12484
rect 3512 12540 3576 12544
rect 3512 12484 3516 12540
rect 3516 12484 3572 12540
rect 3572 12484 3576 12540
rect 3512 12480 3576 12484
rect 3592 12540 3656 12544
rect 3592 12484 3596 12540
rect 3596 12484 3652 12540
rect 3652 12484 3656 12540
rect 3592 12480 3656 12484
rect 8152 12540 8216 12544
rect 8152 12484 8156 12540
rect 8156 12484 8212 12540
rect 8212 12484 8216 12540
rect 8152 12480 8216 12484
rect 8232 12540 8296 12544
rect 8232 12484 8236 12540
rect 8236 12484 8292 12540
rect 8292 12484 8296 12540
rect 8232 12480 8296 12484
rect 8312 12540 8376 12544
rect 8312 12484 8316 12540
rect 8316 12484 8372 12540
rect 8372 12484 8376 12540
rect 8312 12480 8376 12484
rect 8392 12540 8456 12544
rect 8392 12484 8396 12540
rect 8396 12484 8452 12540
rect 8452 12484 8456 12540
rect 8392 12480 8456 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 17752 12540 17816 12544
rect 17752 12484 17756 12540
rect 17756 12484 17812 12540
rect 17812 12484 17816 12540
rect 17752 12480 17816 12484
rect 17832 12540 17896 12544
rect 17832 12484 17836 12540
rect 17836 12484 17892 12540
rect 17892 12484 17896 12540
rect 17832 12480 17896 12484
rect 17912 12540 17976 12544
rect 17912 12484 17916 12540
rect 17916 12484 17972 12540
rect 17972 12484 17976 12540
rect 17912 12480 17976 12484
rect 17992 12540 18056 12544
rect 17992 12484 17996 12540
rect 17996 12484 18052 12540
rect 18052 12484 18056 12540
rect 17992 12480 18056 12484
rect 22552 12540 22616 12544
rect 22552 12484 22556 12540
rect 22556 12484 22612 12540
rect 22612 12484 22616 12540
rect 22552 12480 22616 12484
rect 22632 12540 22696 12544
rect 22632 12484 22636 12540
rect 22636 12484 22692 12540
rect 22692 12484 22696 12540
rect 22632 12480 22696 12484
rect 22712 12540 22776 12544
rect 22712 12484 22716 12540
rect 22716 12484 22772 12540
rect 22772 12484 22776 12540
rect 22712 12480 22776 12484
rect 22792 12540 22856 12544
rect 22792 12484 22796 12540
rect 22796 12484 22852 12540
rect 22852 12484 22856 12540
rect 22792 12480 22856 12484
rect 27352 12540 27416 12544
rect 27352 12484 27356 12540
rect 27356 12484 27412 12540
rect 27412 12484 27416 12540
rect 27352 12480 27416 12484
rect 27432 12540 27496 12544
rect 27432 12484 27436 12540
rect 27436 12484 27492 12540
rect 27492 12484 27496 12540
rect 27432 12480 27496 12484
rect 27512 12540 27576 12544
rect 27512 12484 27516 12540
rect 27516 12484 27572 12540
rect 27572 12484 27576 12540
rect 27512 12480 27576 12484
rect 27592 12540 27656 12544
rect 27592 12484 27596 12540
rect 27596 12484 27652 12540
rect 27652 12484 27656 12540
rect 27592 12480 27656 12484
rect 5752 11996 5816 12000
rect 5752 11940 5756 11996
rect 5756 11940 5812 11996
rect 5812 11940 5816 11996
rect 5752 11936 5816 11940
rect 5832 11996 5896 12000
rect 5832 11940 5836 11996
rect 5836 11940 5892 11996
rect 5892 11940 5896 11996
rect 5832 11936 5896 11940
rect 5912 11996 5976 12000
rect 5912 11940 5916 11996
rect 5916 11940 5972 11996
rect 5972 11940 5976 11996
rect 5912 11936 5976 11940
rect 5992 11996 6056 12000
rect 5992 11940 5996 11996
rect 5996 11940 6052 11996
rect 6052 11940 6056 11996
rect 5992 11936 6056 11940
rect 10552 11996 10616 12000
rect 10552 11940 10556 11996
rect 10556 11940 10612 11996
rect 10612 11940 10616 11996
rect 10552 11936 10616 11940
rect 10632 11996 10696 12000
rect 10632 11940 10636 11996
rect 10636 11940 10692 11996
rect 10692 11940 10696 11996
rect 10632 11936 10696 11940
rect 10712 11996 10776 12000
rect 10712 11940 10716 11996
rect 10716 11940 10772 11996
rect 10772 11940 10776 11996
rect 10712 11936 10776 11940
rect 10792 11996 10856 12000
rect 10792 11940 10796 11996
rect 10796 11940 10852 11996
rect 10852 11940 10856 11996
rect 10792 11936 10856 11940
rect 15352 11996 15416 12000
rect 15352 11940 15356 11996
rect 15356 11940 15412 11996
rect 15412 11940 15416 11996
rect 15352 11936 15416 11940
rect 15432 11996 15496 12000
rect 15432 11940 15436 11996
rect 15436 11940 15492 11996
rect 15492 11940 15496 11996
rect 15432 11936 15496 11940
rect 15512 11996 15576 12000
rect 15512 11940 15516 11996
rect 15516 11940 15572 11996
rect 15572 11940 15576 11996
rect 15512 11936 15576 11940
rect 15592 11996 15656 12000
rect 15592 11940 15596 11996
rect 15596 11940 15652 11996
rect 15652 11940 15656 11996
rect 15592 11936 15656 11940
rect 20152 11996 20216 12000
rect 20152 11940 20156 11996
rect 20156 11940 20212 11996
rect 20212 11940 20216 11996
rect 20152 11936 20216 11940
rect 20232 11996 20296 12000
rect 20232 11940 20236 11996
rect 20236 11940 20292 11996
rect 20292 11940 20296 11996
rect 20232 11936 20296 11940
rect 20312 11996 20376 12000
rect 20312 11940 20316 11996
rect 20316 11940 20372 11996
rect 20372 11940 20376 11996
rect 20312 11936 20376 11940
rect 20392 11996 20456 12000
rect 20392 11940 20396 11996
rect 20396 11940 20452 11996
rect 20452 11940 20456 11996
rect 20392 11936 20456 11940
rect 24952 11996 25016 12000
rect 24952 11940 24956 11996
rect 24956 11940 25012 11996
rect 25012 11940 25016 11996
rect 24952 11936 25016 11940
rect 25032 11996 25096 12000
rect 25032 11940 25036 11996
rect 25036 11940 25092 11996
rect 25092 11940 25096 11996
rect 25032 11936 25096 11940
rect 25112 11996 25176 12000
rect 25112 11940 25116 11996
rect 25116 11940 25172 11996
rect 25172 11940 25176 11996
rect 25112 11936 25176 11940
rect 25192 11996 25256 12000
rect 25192 11940 25196 11996
rect 25196 11940 25252 11996
rect 25252 11940 25256 11996
rect 25192 11936 25256 11940
rect 3352 11452 3416 11456
rect 3352 11396 3356 11452
rect 3356 11396 3412 11452
rect 3412 11396 3416 11452
rect 3352 11392 3416 11396
rect 3432 11452 3496 11456
rect 3432 11396 3436 11452
rect 3436 11396 3492 11452
rect 3492 11396 3496 11452
rect 3432 11392 3496 11396
rect 3512 11452 3576 11456
rect 3512 11396 3516 11452
rect 3516 11396 3572 11452
rect 3572 11396 3576 11452
rect 3512 11392 3576 11396
rect 3592 11452 3656 11456
rect 3592 11396 3596 11452
rect 3596 11396 3652 11452
rect 3652 11396 3656 11452
rect 3592 11392 3656 11396
rect 8152 11452 8216 11456
rect 8152 11396 8156 11452
rect 8156 11396 8212 11452
rect 8212 11396 8216 11452
rect 8152 11392 8216 11396
rect 8232 11452 8296 11456
rect 8232 11396 8236 11452
rect 8236 11396 8292 11452
rect 8292 11396 8296 11452
rect 8232 11392 8296 11396
rect 8312 11452 8376 11456
rect 8312 11396 8316 11452
rect 8316 11396 8372 11452
rect 8372 11396 8376 11452
rect 8312 11392 8376 11396
rect 8392 11452 8456 11456
rect 8392 11396 8396 11452
rect 8396 11396 8452 11452
rect 8452 11396 8456 11452
rect 8392 11392 8456 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 17752 11452 17816 11456
rect 17752 11396 17756 11452
rect 17756 11396 17812 11452
rect 17812 11396 17816 11452
rect 17752 11392 17816 11396
rect 17832 11452 17896 11456
rect 17832 11396 17836 11452
rect 17836 11396 17892 11452
rect 17892 11396 17896 11452
rect 17832 11392 17896 11396
rect 17912 11452 17976 11456
rect 17912 11396 17916 11452
rect 17916 11396 17972 11452
rect 17972 11396 17976 11452
rect 17912 11392 17976 11396
rect 17992 11452 18056 11456
rect 17992 11396 17996 11452
rect 17996 11396 18052 11452
rect 18052 11396 18056 11452
rect 17992 11392 18056 11396
rect 22552 11452 22616 11456
rect 22552 11396 22556 11452
rect 22556 11396 22612 11452
rect 22612 11396 22616 11452
rect 22552 11392 22616 11396
rect 22632 11452 22696 11456
rect 22632 11396 22636 11452
rect 22636 11396 22692 11452
rect 22692 11396 22696 11452
rect 22632 11392 22696 11396
rect 22712 11452 22776 11456
rect 22712 11396 22716 11452
rect 22716 11396 22772 11452
rect 22772 11396 22776 11452
rect 22712 11392 22776 11396
rect 22792 11452 22856 11456
rect 22792 11396 22796 11452
rect 22796 11396 22852 11452
rect 22852 11396 22856 11452
rect 22792 11392 22856 11396
rect 27352 11452 27416 11456
rect 27352 11396 27356 11452
rect 27356 11396 27412 11452
rect 27412 11396 27416 11452
rect 27352 11392 27416 11396
rect 27432 11452 27496 11456
rect 27432 11396 27436 11452
rect 27436 11396 27492 11452
rect 27492 11396 27496 11452
rect 27432 11392 27496 11396
rect 27512 11452 27576 11456
rect 27512 11396 27516 11452
rect 27516 11396 27572 11452
rect 27572 11396 27576 11452
rect 27512 11392 27576 11396
rect 27592 11452 27656 11456
rect 27592 11396 27596 11452
rect 27596 11396 27652 11452
rect 27652 11396 27656 11452
rect 27592 11392 27656 11396
rect 5752 10908 5816 10912
rect 5752 10852 5756 10908
rect 5756 10852 5812 10908
rect 5812 10852 5816 10908
rect 5752 10848 5816 10852
rect 5832 10908 5896 10912
rect 5832 10852 5836 10908
rect 5836 10852 5892 10908
rect 5892 10852 5896 10908
rect 5832 10848 5896 10852
rect 5912 10908 5976 10912
rect 5912 10852 5916 10908
rect 5916 10852 5972 10908
rect 5972 10852 5976 10908
rect 5912 10848 5976 10852
rect 5992 10908 6056 10912
rect 5992 10852 5996 10908
rect 5996 10852 6052 10908
rect 6052 10852 6056 10908
rect 5992 10848 6056 10852
rect 10552 10908 10616 10912
rect 10552 10852 10556 10908
rect 10556 10852 10612 10908
rect 10612 10852 10616 10908
rect 10552 10848 10616 10852
rect 10632 10908 10696 10912
rect 10632 10852 10636 10908
rect 10636 10852 10692 10908
rect 10692 10852 10696 10908
rect 10632 10848 10696 10852
rect 10712 10908 10776 10912
rect 10712 10852 10716 10908
rect 10716 10852 10772 10908
rect 10772 10852 10776 10908
rect 10712 10848 10776 10852
rect 10792 10908 10856 10912
rect 10792 10852 10796 10908
rect 10796 10852 10852 10908
rect 10852 10852 10856 10908
rect 10792 10848 10856 10852
rect 15352 10908 15416 10912
rect 15352 10852 15356 10908
rect 15356 10852 15412 10908
rect 15412 10852 15416 10908
rect 15352 10848 15416 10852
rect 15432 10908 15496 10912
rect 15432 10852 15436 10908
rect 15436 10852 15492 10908
rect 15492 10852 15496 10908
rect 15432 10848 15496 10852
rect 15512 10908 15576 10912
rect 15512 10852 15516 10908
rect 15516 10852 15572 10908
rect 15572 10852 15576 10908
rect 15512 10848 15576 10852
rect 15592 10908 15656 10912
rect 15592 10852 15596 10908
rect 15596 10852 15652 10908
rect 15652 10852 15656 10908
rect 15592 10848 15656 10852
rect 20152 10908 20216 10912
rect 20152 10852 20156 10908
rect 20156 10852 20212 10908
rect 20212 10852 20216 10908
rect 20152 10848 20216 10852
rect 20232 10908 20296 10912
rect 20232 10852 20236 10908
rect 20236 10852 20292 10908
rect 20292 10852 20296 10908
rect 20232 10848 20296 10852
rect 20312 10908 20376 10912
rect 20312 10852 20316 10908
rect 20316 10852 20372 10908
rect 20372 10852 20376 10908
rect 20312 10848 20376 10852
rect 20392 10908 20456 10912
rect 20392 10852 20396 10908
rect 20396 10852 20452 10908
rect 20452 10852 20456 10908
rect 20392 10848 20456 10852
rect 24952 10908 25016 10912
rect 24952 10852 24956 10908
rect 24956 10852 25012 10908
rect 25012 10852 25016 10908
rect 24952 10848 25016 10852
rect 25032 10908 25096 10912
rect 25032 10852 25036 10908
rect 25036 10852 25092 10908
rect 25092 10852 25096 10908
rect 25032 10848 25096 10852
rect 25112 10908 25176 10912
rect 25112 10852 25116 10908
rect 25116 10852 25172 10908
rect 25172 10852 25176 10908
rect 25112 10848 25176 10852
rect 25192 10908 25256 10912
rect 25192 10852 25196 10908
rect 25196 10852 25252 10908
rect 25252 10852 25256 10908
rect 25192 10848 25256 10852
rect 3352 10364 3416 10368
rect 3352 10308 3356 10364
rect 3356 10308 3412 10364
rect 3412 10308 3416 10364
rect 3352 10304 3416 10308
rect 3432 10364 3496 10368
rect 3432 10308 3436 10364
rect 3436 10308 3492 10364
rect 3492 10308 3496 10364
rect 3432 10304 3496 10308
rect 3512 10364 3576 10368
rect 3512 10308 3516 10364
rect 3516 10308 3572 10364
rect 3572 10308 3576 10364
rect 3512 10304 3576 10308
rect 3592 10364 3656 10368
rect 3592 10308 3596 10364
rect 3596 10308 3652 10364
rect 3652 10308 3656 10364
rect 3592 10304 3656 10308
rect 8152 10364 8216 10368
rect 8152 10308 8156 10364
rect 8156 10308 8212 10364
rect 8212 10308 8216 10364
rect 8152 10304 8216 10308
rect 8232 10364 8296 10368
rect 8232 10308 8236 10364
rect 8236 10308 8292 10364
rect 8292 10308 8296 10364
rect 8232 10304 8296 10308
rect 8312 10364 8376 10368
rect 8312 10308 8316 10364
rect 8316 10308 8372 10364
rect 8372 10308 8376 10364
rect 8312 10304 8376 10308
rect 8392 10364 8456 10368
rect 8392 10308 8396 10364
rect 8396 10308 8452 10364
rect 8452 10308 8456 10364
rect 8392 10304 8456 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 17752 10364 17816 10368
rect 17752 10308 17756 10364
rect 17756 10308 17812 10364
rect 17812 10308 17816 10364
rect 17752 10304 17816 10308
rect 17832 10364 17896 10368
rect 17832 10308 17836 10364
rect 17836 10308 17892 10364
rect 17892 10308 17896 10364
rect 17832 10304 17896 10308
rect 17912 10364 17976 10368
rect 17912 10308 17916 10364
rect 17916 10308 17972 10364
rect 17972 10308 17976 10364
rect 17912 10304 17976 10308
rect 17992 10364 18056 10368
rect 17992 10308 17996 10364
rect 17996 10308 18052 10364
rect 18052 10308 18056 10364
rect 17992 10304 18056 10308
rect 22552 10364 22616 10368
rect 22552 10308 22556 10364
rect 22556 10308 22612 10364
rect 22612 10308 22616 10364
rect 22552 10304 22616 10308
rect 22632 10364 22696 10368
rect 22632 10308 22636 10364
rect 22636 10308 22692 10364
rect 22692 10308 22696 10364
rect 22632 10304 22696 10308
rect 22712 10364 22776 10368
rect 22712 10308 22716 10364
rect 22716 10308 22772 10364
rect 22772 10308 22776 10364
rect 22712 10304 22776 10308
rect 22792 10364 22856 10368
rect 22792 10308 22796 10364
rect 22796 10308 22852 10364
rect 22852 10308 22856 10364
rect 22792 10304 22856 10308
rect 27352 10364 27416 10368
rect 27352 10308 27356 10364
rect 27356 10308 27412 10364
rect 27412 10308 27416 10364
rect 27352 10304 27416 10308
rect 27432 10364 27496 10368
rect 27432 10308 27436 10364
rect 27436 10308 27492 10364
rect 27492 10308 27496 10364
rect 27432 10304 27496 10308
rect 27512 10364 27576 10368
rect 27512 10308 27516 10364
rect 27516 10308 27572 10364
rect 27572 10308 27576 10364
rect 27512 10304 27576 10308
rect 27592 10364 27656 10368
rect 27592 10308 27596 10364
rect 27596 10308 27652 10364
rect 27652 10308 27656 10364
rect 27592 10304 27656 10308
rect 5752 9820 5816 9824
rect 5752 9764 5756 9820
rect 5756 9764 5812 9820
rect 5812 9764 5816 9820
rect 5752 9760 5816 9764
rect 5832 9820 5896 9824
rect 5832 9764 5836 9820
rect 5836 9764 5892 9820
rect 5892 9764 5896 9820
rect 5832 9760 5896 9764
rect 5912 9820 5976 9824
rect 5912 9764 5916 9820
rect 5916 9764 5972 9820
rect 5972 9764 5976 9820
rect 5912 9760 5976 9764
rect 5992 9820 6056 9824
rect 5992 9764 5996 9820
rect 5996 9764 6052 9820
rect 6052 9764 6056 9820
rect 5992 9760 6056 9764
rect 10552 9820 10616 9824
rect 10552 9764 10556 9820
rect 10556 9764 10612 9820
rect 10612 9764 10616 9820
rect 10552 9760 10616 9764
rect 10632 9820 10696 9824
rect 10632 9764 10636 9820
rect 10636 9764 10692 9820
rect 10692 9764 10696 9820
rect 10632 9760 10696 9764
rect 10712 9820 10776 9824
rect 10712 9764 10716 9820
rect 10716 9764 10772 9820
rect 10772 9764 10776 9820
rect 10712 9760 10776 9764
rect 10792 9820 10856 9824
rect 10792 9764 10796 9820
rect 10796 9764 10852 9820
rect 10852 9764 10856 9820
rect 10792 9760 10856 9764
rect 15352 9820 15416 9824
rect 15352 9764 15356 9820
rect 15356 9764 15412 9820
rect 15412 9764 15416 9820
rect 15352 9760 15416 9764
rect 15432 9820 15496 9824
rect 15432 9764 15436 9820
rect 15436 9764 15492 9820
rect 15492 9764 15496 9820
rect 15432 9760 15496 9764
rect 15512 9820 15576 9824
rect 15512 9764 15516 9820
rect 15516 9764 15572 9820
rect 15572 9764 15576 9820
rect 15512 9760 15576 9764
rect 15592 9820 15656 9824
rect 15592 9764 15596 9820
rect 15596 9764 15652 9820
rect 15652 9764 15656 9820
rect 15592 9760 15656 9764
rect 20152 9820 20216 9824
rect 20152 9764 20156 9820
rect 20156 9764 20212 9820
rect 20212 9764 20216 9820
rect 20152 9760 20216 9764
rect 20232 9820 20296 9824
rect 20232 9764 20236 9820
rect 20236 9764 20292 9820
rect 20292 9764 20296 9820
rect 20232 9760 20296 9764
rect 20312 9820 20376 9824
rect 20312 9764 20316 9820
rect 20316 9764 20372 9820
rect 20372 9764 20376 9820
rect 20312 9760 20376 9764
rect 20392 9820 20456 9824
rect 20392 9764 20396 9820
rect 20396 9764 20452 9820
rect 20452 9764 20456 9820
rect 20392 9760 20456 9764
rect 24952 9820 25016 9824
rect 24952 9764 24956 9820
rect 24956 9764 25012 9820
rect 25012 9764 25016 9820
rect 24952 9760 25016 9764
rect 25032 9820 25096 9824
rect 25032 9764 25036 9820
rect 25036 9764 25092 9820
rect 25092 9764 25096 9820
rect 25032 9760 25096 9764
rect 25112 9820 25176 9824
rect 25112 9764 25116 9820
rect 25116 9764 25172 9820
rect 25172 9764 25176 9820
rect 25112 9760 25176 9764
rect 25192 9820 25256 9824
rect 25192 9764 25196 9820
rect 25196 9764 25252 9820
rect 25252 9764 25256 9820
rect 25192 9760 25256 9764
rect 3352 9276 3416 9280
rect 3352 9220 3356 9276
rect 3356 9220 3412 9276
rect 3412 9220 3416 9276
rect 3352 9216 3416 9220
rect 3432 9276 3496 9280
rect 3432 9220 3436 9276
rect 3436 9220 3492 9276
rect 3492 9220 3496 9276
rect 3432 9216 3496 9220
rect 3512 9276 3576 9280
rect 3512 9220 3516 9276
rect 3516 9220 3572 9276
rect 3572 9220 3576 9276
rect 3512 9216 3576 9220
rect 3592 9276 3656 9280
rect 3592 9220 3596 9276
rect 3596 9220 3652 9276
rect 3652 9220 3656 9276
rect 3592 9216 3656 9220
rect 8152 9276 8216 9280
rect 8152 9220 8156 9276
rect 8156 9220 8212 9276
rect 8212 9220 8216 9276
rect 8152 9216 8216 9220
rect 8232 9276 8296 9280
rect 8232 9220 8236 9276
rect 8236 9220 8292 9276
rect 8292 9220 8296 9276
rect 8232 9216 8296 9220
rect 8312 9276 8376 9280
rect 8312 9220 8316 9276
rect 8316 9220 8372 9276
rect 8372 9220 8376 9276
rect 8312 9216 8376 9220
rect 8392 9276 8456 9280
rect 8392 9220 8396 9276
rect 8396 9220 8452 9276
rect 8452 9220 8456 9276
rect 8392 9216 8456 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 17752 9276 17816 9280
rect 17752 9220 17756 9276
rect 17756 9220 17812 9276
rect 17812 9220 17816 9276
rect 17752 9216 17816 9220
rect 17832 9276 17896 9280
rect 17832 9220 17836 9276
rect 17836 9220 17892 9276
rect 17892 9220 17896 9276
rect 17832 9216 17896 9220
rect 17912 9276 17976 9280
rect 17912 9220 17916 9276
rect 17916 9220 17972 9276
rect 17972 9220 17976 9276
rect 17912 9216 17976 9220
rect 17992 9276 18056 9280
rect 17992 9220 17996 9276
rect 17996 9220 18052 9276
rect 18052 9220 18056 9276
rect 17992 9216 18056 9220
rect 22552 9276 22616 9280
rect 22552 9220 22556 9276
rect 22556 9220 22612 9276
rect 22612 9220 22616 9276
rect 22552 9216 22616 9220
rect 22632 9276 22696 9280
rect 22632 9220 22636 9276
rect 22636 9220 22692 9276
rect 22692 9220 22696 9276
rect 22632 9216 22696 9220
rect 22712 9276 22776 9280
rect 22712 9220 22716 9276
rect 22716 9220 22772 9276
rect 22772 9220 22776 9276
rect 22712 9216 22776 9220
rect 22792 9276 22856 9280
rect 22792 9220 22796 9276
rect 22796 9220 22852 9276
rect 22852 9220 22856 9276
rect 22792 9216 22856 9220
rect 27352 9276 27416 9280
rect 27352 9220 27356 9276
rect 27356 9220 27412 9276
rect 27412 9220 27416 9276
rect 27352 9216 27416 9220
rect 27432 9276 27496 9280
rect 27432 9220 27436 9276
rect 27436 9220 27492 9276
rect 27492 9220 27496 9276
rect 27432 9216 27496 9220
rect 27512 9276 27576 9280
rect 27512 9220 27516 9276
rect 27516 9220 27572 9276
rect 27572 9220 27576 9276
rect 27512 9216 27576 9220
rect 27592 9276 27656 9280
rect 27592 9220 27596 9276
rect 27596 9220 27652 9276
rect 27652 9220 27656 9276
rect 27592 9216 27656 9220
rect 5752 8732 5816 8736
rect 5752 8676 5756 8732
rect 5756 8676 5812 8732
rect 5812 8676 5816 8732
rect 5752 8672 5816 8676
rect 5832 8732 5896 8736
rect 5832 8676 5836 8732
rect 5836 8676 5892 8732
rect 5892 8676 5896 8732
rect 5832 8672 5896 8676
rect 5912 8732 5976 8736
rect 5912 8676 5916 8732
rect 5916 8676 5972 8732
rect 5972 8676 5976 8732
rect 5912 8672 5976 8676
rect 5992 8732 6056 8736
rect 5992 8676 5996 8732
rect 5996 8676 6052 8732
rect 6052 8676 6056 8732
rect 5992 8672 6056 8676
rect 10552 8732 10616 8736
rect 10552 8676 10556 8732
rect 10556 8676 10612 8732
rect 10612 8676 10616 8732
rect 10552 8672 10616 8676
rect 10632 8732 10696 8736
rect 10632 8676 10636 8732
rect 10636 8676 10692 8732
rect 10692 8676 10696 8732
rect 10632 8672 10696 8676
rect 10712 8732 10776 8736
rect 10712 8676 10716 8732
rect 10716 8676 10772 8732
rect 10772 8676 10776 8732
rect 10712 8672 10776 8676
rect 10792 8732 10856 8736
rect 10792 8676 10796 8732
rect 10796 8676 10852 8732
rect 10852 8676 10856 8732
rect 10792 8672 10856 8676
rect 15352 8732 15416 8736
rect 15352 8676 15356 8732
rect 15356 8676 15412 8732
rect 15412 8676 15416 8732
rect 15352 8672 15416 8676
rect 15432 8732 15496 8736
rect 15432 8676 15436 8732
rect 15436 8676 15492 8732
rect 15492 8676 15496 8732
rect 15432 8672 15496 8676
rect 15512 8732 15576 8736
rect 15512 8676 15516 8732
rect 15516 8676 15572 8732
rect 15572 8676 15576 8732
rect 15512 8672 15576 8676
rect 15592 8732 15656 8736
rect 15592 8676 15596 8732
rect 15596 8676 15652 8732
rect 15652 8676 15656 8732
rect 15592 8672 15656 8676
rect 20152 8732 20216 8736
rect 20152 8676 20156 8732
rect 20156 8676 20212 8732
rect 20212 8676 20216 8732
rect 20152 8672 20216 8676
rect 20232 8732 20296 8736
rect 20232 8676 20236 8732
rect 20236 8676 20292 8732
rect 20292 8676 20296 8732
rect 20232 8672 20296 8676
rect 20312 8732 20376 8736
rect 20312 8676 20316 8732
rect 20316 8676 20372 8732
rect 20372 8676 20376 8732
rect 20312 8672 20376 8676
rect 20392 8732 20456 8736
rect 20392 8676 20396 8732
rect 20396 8676 20452 8732
rect 20452 8676 20456 8732
rect 20392 8672 20456 8676
rect 24952 8732 25016 8736
rect 24952 8676 24956 8732
rect 24956 8676 25012 8732
rect 25012 8676 25016 8732
rect 24952 8672 25016 8676
rect 25032 8732 25096 8736
rect 25032 8676 25036 8732
rect 25036 8676 25092 8732
rect 25092 8676 25096 8732
rect 25032 8672 25096 8676
rect 25112 8732 25176 8736
rect 25112 8676 25116 8732
rect 25116 8676 25172 8732
rect 25172 8676 25176 8732
rect 25112 8672 25176 8676
rect 25192 8732 25256 8736
rect 25192 8676 25196 8732
rect 25196 8676 25252 8732
rect 25252 8676 25256 8732
rect 25192 8672 25256 8676
rect 3352 8188 3416 8192
rect 3352 8132 3356 8188
rect 3356 8132 3412 8188
rect 3412 8132 3416 8188
rect 3352 8128 3416 8132
rect 3432 8188 3496 8192
rect 3432 8132 3436 8188
rect 3436 8132 3492 8188
rect 3492 8132 3496 8188
rect 3432 8128 3496 8132
rect 3512 8188 3576 8192
rect 3512 8132 3516 8188
rect 3516 8132 3572 8188
rect 3572 8132 3576 8188
rect 3512 8128 3576 8132
rect 3592 8188 3656 8192
rect 3592 8132 3596 8188
rect 3596 8132 3652 8188
rect 3652 8132 3656 8188
rect 3592 8128 3656 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 8312 8188 8376 8192
rect 8312 8132 8316 8188
rect 8316 8132 8372 8188
rect 8372 8132 8376 8188
rect 8312 8128 8376 8132
rect 8392 8188 8456 8192
rect 8392 8132 8396 8188
rect 8396 8132 8452 8188
rect 8452 8132 8456 8188
rect 8392 8128 8456 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 17752 8188 17816 8192
rect 17752 8132 17756 8188
rect 17756 8132 17812 8188
rect 17812 8132 17816 8188
rect 17752 8128 17816 8132
rect 17832 8188 17896 8192
rect 17832 8132 17836 8188
rect 17836 8132 17892 8188
rect 17892 8132 17896 8188
rect 17832 8128 17896 8132
rect 17912 8188 17976 8192
rect 17912 8132 17916 8188
rect 17916 8132 17972 8188
rect 17972 8132 17976 8188
rect 17912 8128 17976 8132
rect 17992 8188 18056 8192
rect 17992 8132 17996 8188
rect 17996 8132 18052 8188
rect 18052 8132 18056 8188
rect 17992 8128 18056 8132
rect 22552 8188 22616 8192
rect 22552 8132 22556 8188
rect 22556 8132 22612 8188
rect 22612 8132 22616 8188
rect 22552 8128 22616 8132
rect 22632 8188 22696 8192
rect 22632 8132 22636 8188
rect 22636 8132 22692 8188
rect 22692 8132 22696 8188
rect 22632 8128 22696 8132
rect 22712 8188 22776 8192
rect 22712 8132 22716 8188
rect 22716 8132 22772 8188
rect 22772 8132 22776 8188
rect 22712 8128 22776 8132
rect 22792 8188 22856 8192
rect 22792 8132 22796 8188
rect 22796 8132 22852 8188
rect 22852 8132 22856 8188
rect 22792 8128 22856 8132
rect 27352 8188 27416 8192
rect 27352 8132 27356 8188
rect 27356 8132 27412 8188
rect 27412 8132 27416 8188
rect 27352 8128 27416 8132
rect 27432 8188 27496 8192
rect 27432 8132 27436 8188
rect 27436 8132 27492 8188
rect 27492 8132 27496 8188
rect 27432 8128 27496 8132
rect 27512 8188 27576 8192
rect 27512 8132 27516 8188
rect 27516 8132 27572 8188
rect 27572 8132 27576 8188
rect 27512 8128 27576 8132
rect 27592 8188 27656 8192
rect 27592 8132 27596 8188
rect 27596 8132 27652 8188
rect 27652 8132 27656 8188
rect 27592 8128 27656 8132
rect 5752 7644 5816 7648
rect 5752 7588 5756 7644
rect 5756 7588 5812 7644
rect 5812 7588 5816 7644
rect 5752 7584 5816 7588
rect 5832 7644 5896 7648
rect 5832 7588 5836 7644
rect 5836 7588 5892 7644
rect 5892 7588 5896 7644
rect 5832 7584 5896 7588
rect 5912 7644 5976 7648
rect 5912 7588 5916 7644
rect 5916 7588 5972 7644
rect 5972 7588 5976 7644
rect 5912 7584 5976 7588
rect 5992 7644 6056 7648
rect 5992 7588 5996 7644
rect 5996 7588 6052 7644
rect 6052 7588 6056 7644
rect 5992 7584 6056 7588
rect 10552 7644 10616 7648
rect 10552 7588 10556 7644
rect 10556 7588 10612 7644
rect 10612 7588 10616 7644
rect 10552 7584 10616 7588
rect 10632 7644 10696 7648
rect 10632 7588 10636 7644
rect 10636 7588 10692 7644
rect 10692 7588 10696 7644
rect 10632 7584 10696 7588
rect 10712 7644 10776 7648
rect 10712 7588 10716 7644
rect 10716 7588 10772 7644
rect 10772 7588 10776 7644
rect 10712 7584 10776 7588
rect 10792 7644 10856 7648
rect 10792 7588 10796 7644
rect 10796 7588 10852 7644
rect 10852 7588 10856 7644
rect 10792 7584 10856 7588
rect 15352 7644 15416 7648
rect 15352 7588 15356 7644
rect 15356 7588 15412 7644
rect 15412 7588 15416 7644
rect 15352 7584 15416 7588
rect 15432 7644 15496 7648
rect 15432 7588 15436 7644
rect 15436 7588 15492 7644
rect 15492 7588 15496 7644
rect 15432 7584 15496 7588
rect 15512 7644 15576 7648
rect 15512 7588 15516 7644
rect 15516 7588 15572 7644
rect 15572 7588 15576 7644
rect 15512 7584 15576 7588
rect 15592 7644 15656 7648
rect 15592 7588 15596 7644
rect 15596 7588 15652 7644
rect 15652 7588 15656 7644
rect 15592 7584 15656 7588
rect 20152 7644 20216 7648
rect 20152 7588 20156 7644
rect 20156 7588 20212 7644
rect 20212 7588 20216 7644
rect 20152 7584 20216 7588
rect 20232 7644 20296 7648
rect 20232 7588 20236 7644
rect 20236 7588 20292 7644
rect 20292 7588 20296 7644
rect 20232 7584 20296 7588
rect 20312 7644 20376 7648
rect 20312 7588 20316 7644
rect 20316 7588 20372 7644
rect 20372 7588 20376 7644
rect 20312 7584 20376 7588
rect 20392 7644 20456 7648
rect 20392 7588 20396 7644
rect 20396 7588 20452 7644
rect 20452 7588 20456 7644
rect 20392 7584 20456 7588
rect 24952 7644 25016 7648
rect 24952 7588 24956 7644
rect 24956 7588 25012 7644
rect 25012 7588 25016 7644
rect 24952 7584 25016 7588
rect 25032 7644 25096 7648
rect 25032 7588 25036 7644
rect 25036 7588 25092 7644
rect 25092 7588 25096 7644
rect 25032 7584 25096 7588
rect 25112 7644 25176 7648
rect 25112 7588 25116 7644
rect 25116 7588 25172 7644
rect 25172 7588 25176 7644
rect 25112 7584 25176 7588
rect 25192 7644 25256 7648
rect 25192 7588 25196 7644
rect 25196 7588 25252 7644
rect 25252 7588 25256 7644
rect 25192 7584 25256 7588
rect 3352 7100 3416 7104
rect 3352 7044 3356 7100
rect 3356 7044 3412 7100
rect 3412 7044 3416 7100
rect 3352 7040 3416 7044
rect 3432 7100 3496 7104
rect 3432 7044 3436 7100
rect 3436 7044 3492 7100
rect 3492 7044 3496 7100
rect 3432 7040 3496 7044
rect 3512 7100 3576 7104
rect 3512 7044 3516 7100
rect 3516 7044 3572 7100
rect 3572 7044 3576 7100
rect 3512 7040 3576 7044
rect 3592 7100 3656 7104
rect 3592 7044 3596 7100
rect 3596 7044 3652 7100
rect 3652 7044 3656 7100
rect 3592 7040 3656 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 8312 7100 8376 7104
rect 8312 7044 8316 7100
rect 8316 7044 8372 7100
rect 8372 7044 8376 7100
rect 8312 7040 8376 7044
rect 8392 7100 8456 7104
rect 8392 7044 8396 7100
rect 8396 7044 8452 7100
rect 8452 7044 8456 7100
rect 8392 7040 8456 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 17752 7100 17816 7104
rect 17752 7044 17756 7100
rect 17756 7044 17812 7100
rect 17812 7044 17816 7100
rect 17752 7040 17816 7044
rect 17832 7100 17896 7104
rect 17832 7044 17836 7100
rect 17836 7044 17892 7100
rect 17892 7044 17896 7100
rect 17832 7040 17896 7044
rect 17912 7100 17976 7104
rect 17912 7044 17916 7100
rect 17916 7044 17972 7100
rect 17972 7044 17976 7100
rect 17912 7040 17976 7044
rect 17992 7100 18056 7104
rect 17992 7044 17996 7100
rect 17996 7044 18052 7100
rect 18052 7044 18056 7100
rect 17992 7040 18056 7044
rect 22552 7100 22616 7104
rect 22552 7044 22556 7100
rect 22556 7044 22612 7100
rect 22612 7044 22616 7100
rect 22552 7040 22616 7044
rect 22632 7100 22696 7104
rect 22632 7044 22636 7100
rect 22636 7044 22692 7100
rect 22692 7044 22696 7100
rect 22632 7040 22696 7044
rect 22712 7100 22776 7104
rect 22712 7044 22716 7100
rect 22716 7044 22772 7100
rect 22772 7044 22776 7100
rect 22712 7040 22776 7044
rect 22792 7100 22856 7104
rect 22792 7044 22796 7100
rect 22796 7044 22852 7100
rect 22852 7044 22856 7100
rect 22792 7040 22856 7044
rect 27352 7100 27416 7104
rect 27352 7044 27356 7100
rect 27356 7044 27412 7100
rect 27412 7044 27416 7100
rect 27352 7040 27416 7044
rect 27432 7100 27496 7104
rect 27432 7044 27436 7100
rect 27436 7044 27492 7100
rect 27492 7044 27496 7100
rect 27432 7040 27496 7044
rect 27512 7100 27576 7104
rect 27512 7044 27516 7100
rect 27516 7044 27572 7100
rect 27572 7044 27576 7100
rect 27512 7040 27576 7044
rect 27592 7100 27656 7104
rect 27592 7044 27596 7100
rect 27596 7044 27652 7100
rect 27652 7044 27656 7100
rect 27592 7040 27656 7044
rect 5752 6556 5816 6560
rect 5752 6500 5756 6556
rect 5756 6500 5812 6556
rect 5812 6500 5816 6556
rect 5752 6496 5816 6500
rect 5832 6556 5896 6560
rect 5832 6500 5836 6556
rect 5836 6500 5892 6556
rect 5892 6500 5896 6556
rect 5832 6496 5896 6500
rect 5912 6556 5976 6560
rect 5912 6500 5916 6556
rect 5916 6500 5972 6556
rect 5972 6500 5976 6556
rect 5912 6496 5976 6500
rect 5992 6556 6056 6560
rect 5992 6500 5996 6556
rect 5996 6500 6052 6556
rect 6052 6500 6056 6556
rect 5992 6496 6056 6500
rect 10552 6556 10616 6560
rect 10552 6500 10556 6556
rect 10556 6500 10612 6556
rect 10612 6500 10616 6556
rect 10552 6496 10616 6500
rect 10632 6556 10696 6560
rect 10632 6500 10636 6556
rect 10636 6500 10692 6556
rect 10692 6500 10696 6556
rect 10632 6496 10696 6500
rect 10712 6556 10776 6560
rect 10712 6500 10716 6556
rect 10716 6500 10772 6556
rect 10772 6500 10776 6556
rect 10712 6496 10776 6500
rect 10792 6556 10856 6560
rect 10792 6500 10796 6556
rect 10796 6500 10852 6556
rect 10852 6500 10856 6556
rect 10792 6496 10856 6500
rect 15352 6556 15416 6560
rect 15352 6500 15356 6556
rect 15356 6500 15412 6556
rect 15412 6500 15416 6556
rect 15352 6496 15416 6500
rect 15432 6556 15496 6560
rect 15432 6500 15436 6556
rect 15436 6500 15492 6556
rect 15492 6500 15496 6556
rect 15432 6496 15496 6500
rect 15512 6556 15576 6560
rect 15512 6500 15516 6556
rect 15516 6500 15572 6556
rect 15572 6500 15576 6556
rect 15512 6496 15576 6500
rect 15592 6556 15656 6560
rect 15592 6500 15596 6556
rect 15596 6500 15652 6556
rect 15652 6500 15656 6556
rect 15592 6496 15656 6500
rect 20152 6556 20216 6560
rect 20152 6500 20156 6556
rect 20156 6500 20212 6556
rect 20212 6500 20216 6556
rect 20152 6496 20216 6500
rect 20232 6556 20296 6560
rect 20232 6500 20236 6556
rect 20236 6500 20292 6556
rect 20292 6500 20296 6556
rect 20232 6496 20296 6500
rect 20312 6556 20376 6560
rect 20312 6500 20316 6556
rect 20316 6500 20372 6556
rect 20372 6500 20376 6556
rect 20312 6496 20376 6500
rect 20392 6556 20456 6560
rect 20392 6500 20396 6556
rect 20396 6500 20452 6556
rect 20452 6500 20456 6556
rect 20392 6496 20456 6500
rect 24952 6556 25016 6560
rect 24952 6500 24956 6556
rect 24956 6500 25012 6556
rect 25012 6500 25016 6556
rect 24952 6496 25016 6500
rect 25032 6556 25096 6560
rect 25032 6500 25036 6556
rect 25036 6500 25092 6556
rect 25092 6500 25096 6556
rect 25032 6496 25096 6500
rect 25112 6556 25176 6560
rect 25112 6500 25116 6556
rect 25116 6500 25172 6556
rect 25172 6500 25176 6556
rect 25112 6496 25176 6500
rect 25192 6556 25256 6560
rect 25192 6500 25196 6556
rect 25196 6500 25252 6556
rect 25252 6500 25256 6556
rect 25192 6496 25256 6500
rect 3352 6012 3416 6016
rect 3352 5956 3356 6012
rect 3356 5956 3412 6012
rect 3412 5956 3416 6012
rect 3352 5952 3416 5956
rect 3432 6012 3496 6016
rect 3432 5956 3436 6012
rect 3436 5956 3492 6012
rect 3492 5956 3496 6012
rect 3432 5952 3496 5956
rect 3512 6012 3576 6016
rect 3512 5956 3516 6012
rect 3516 5956 3572 6012
rect 3572 5956 3576 6012
rect 3512 5952 3576 5956
rect 3592 6012 3656 6016
rect 3592 5956 3596 6012
rect 3596 5956 3652 6012
rect 3652 5956 3656 6012
rect 3592 5952 3656 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 8312 6012 8376 6016
rect 8312 5956 8316 6012
rect 8316 5956 8372 6012
rect 8372 5956 8376 6012
rect 8312 5952 8376 5956
rect 8392 6012 8456 6016
rect 8392 5956 8396 6012
rect 8396 5956 8452 6012
rect 8452 5956 8456 6012
rect 8392 5952 8456 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 17752 6012 17816 6016
rect 17752 5956 17756 6012
rect 17756 5956 17812 6012
rect 17812 5956 17816 6012
rect 17752 5952 17816 5956
rect 17832 6012 17896 6016
rect 17832 5956 17836 6012
rect 17836 5956 17892 6012
rect 17892 5956 17896 6012
rect 17832 5952 17896 5956
rect 17912 6012 17976 6016
rect 17912 5956 17916 6012
rect 17916 5956 17972 6012
rect 17972 5956 17976 6012
rect 17912 5952 17976 5956
rect 17992 6012 18056 6016
rect 17992 5956 17996 6012
rect 17996 5956 18052 6012
rect 18052 5956 18056 6012
rect 17992 5952 18056 5956
rect 22552 6012 22616 6016
rect 22552 5956 22556 6012
rect 22556 5956 22612 6012
rect 22612 5956 22616 6012
rect 22552 5952 22616 5956
rect 22632 6012 22696 6016
rect 22632 5956 22636 6012
rect 22636 5956 22692 6012
rect 22692 5956 22696 6012
rect 22632 5952 22696 5956
rect 22712 6012 22776 6016
rect 22712 5956 22716 6012
rect 22716 5956 22772 6012
rect 22772 5956 22776 6012
rect 22712 5952 22776 5956
rect 22792 6012 22856 6016
rect 22792 5956 22796 6012
rect 22796 5956 22852 6012
rect 22852 5956 22856 6012
rect 22792 5952 22856 5956
rect 27352 6012 27416 6016
rect 27352 5956 27356 6012
rect 27356 5956 27412 6012
rect 27412 5956 27416 6012
rect 27352 5952 27416 5956
rect 27432 6012 27496 6016
rect 27432 5956 27436 6012
rect 27436 5956 27492 6012
rect 27492 5956 27496 6012
rect 27432 5952 27496 5956
rect 27512 6012 27576 6016
rect 27512 5956 27516 6012
rect 27516 5956 27572 6012
rect 27572 5956 27576 6012
rect 27512 5952 27576 5956
rect 27592 6012 27656 6016
rect 27592 5956 27596 6012
rect 27596 5956 27652 6012
rect 27652 5956 27656 6012
rect 27592 5952 27656 5956
rect 5752 5468 5816 5472
rect 5752 5412 5756 5468
rect 5756 5412 5812 5468
rect 5812 5412 5816 5468
rect 5752 5408 5816 5412
rect 5832 5468 5896 5472
rect 5832 5412 5836 5468
rect 5836 5412 5892 5468
rect 5892 5412 5896 5468
rect 5832 5408 5896 5412
rect 5912 5468 5976 5472
rect 5912 5412 5916 5468
rect 5916 5412 5972 5468
rect 5972 5412 5976 5468
rect 5912 5408 5976 5412
rect 5992 5468 6056 5472
rect 5992 5412 5996 5468
rect 5996 5412 6052 5468
rect 6052 5412 6056 5468
rect 5992 5408 6056 5412
rect 10552 5468 10616 5472
rect 10552 5412 10556 5468
rect 10556 5412 10612 5468
rect 10612 5412 10616 5468
rect 10552 5408 10616 5412
rect 10632 5468 10696 5472
rect 10632 5412 10636 5468
rect 10636 5412 10692 5468
rect 10692 5412 10696 5468
rect 10632 5408 10696 5412
rect 10712 5468 10776 5472
rect 10712 5412 10716 5468
rect 10716 5412 10772 5468
rect 10772 5412 10776 5468
rect 10712 5408 10776 5412
rect 10792 5468 10856 5472
rect 10792 5412 10796 5468
rect 10796 5412 10852 5468
rect 10852 5412 10856 5468
rect 10792 5408 10856 5412
rect 15352 5468 15416 5472
rect 15352 5412 15356 5468
rect 15356 5412 15412 5468
rect 15412 5412 15416 5468
rect 15352 5408 15416 5412
rect 15432 5468 15496 5472
rect 15432 5412 15436 5468
rect 15436 5412 15492 5468
rect 15492 5412 15496 5468
rect 15432 5408 15496 5412
rect 15512 5468 15576 5472
rect 15512 5412 15516 5468
rect 15516 5412 15572 5468
rect 15572 5412 15576 5468
rect 15512 5408 15576 5412
rect 15592 5468 15656 5472
rect 15592 5412 15596 5468
rect 15596 5412 15652 5468
rect 15652 5412 15656 5468
rect 15592 5408 15656 5412
rect 20152 5468 20216 5472
rect 20152 5412 20156 5468
rect 20156 5412 20212 5468
rect 20212 5412 20216 5468
rect 20152 5408 20216 5412
rect 20232 5468 20296 5472
rect 20232 5412 20236 5468
rect 20236 5412 20292 5468
rect 20292 5412 20296 5468
rect 20232 5408 20296 5412
rect 20312 5468 20376 5472
rect 20312 5412 20316 5468
rect 20316 5412 20372 5468
rect 20372 5412 20376 5468
rect 20312 5408 20376 5412
rect 20392 5468 20456 5472
rect 20392 5412 20396 5468
rect 20396 5412 20452 5468
rect 20452 5412 20456 5468
rect 20392 5408 20456 5412
rect 24952 5468 25016 5472
rect 24952 5412 24956 5468
rect 24956 5412 25012 5468
rect 25012 5412 25016 5468
rect 24952 5408 25016 5412
rect 25032 5468 25096 5472
rect 25032 5412 25036 5468
rect 25036 5412 25092 5468
rect 25092 5412 25096 5468
rect 25032 5408 25096 5412
rect 25112 5468 25176 5472
rect 25112 5412 25116 5468
rect 25116 5412 25172 5468
rect 25172 5412 25176 5468
rect 25112 5408 25176 5412
rect 25192 5468 25256 5472
rect 25192 5412 25196 5468
rect 25196 5412 25252 5468
rect 25252 5412 25256 5468
rect 25192 5408 25256 5412
rect 3352 4924 3416 4928
rect 3352 4868 3356 4924
rect 3356 4868 3412 4924
rect 3412 4868 3416 4924
rect 3352 4864 3416 4868
rect 3432 4924 3496 4928
rect 3432 4868 3436 4924
rect 3436 4868 3492 4924
rect 3492 4868 3496 4924
rect 3432 4864 3496 4868
rect 3512 4924 3576 4928
rect 3512 4868 3516 4924
rect 3516 4868 3572 4924
rect 3572 4868 3576 4924
rect 3512 4864 3576 4868
rect 3592 4924 3656 4928
rect 3592 4868 3596 4924
rect 3596 4868 3652 4924
rect 3652 4868 3656 4924
rect 3592 4864 3656 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 8312 4924 8376 4928
rect 8312 4868 8316 4924
rect 8316 4868 8372 4924
rect 8372 4868 8376 4924
rect 8312 4864 8376 4868
rect 8392 4924 8456 4928
rect 8392 4868 8396 4924
rect 8396 4868 8452 4924
rect 8452 4868 8456 4924
rect 8392 4864 8456 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 17752 4924 17816 4928
rect 17752 4868 17756 4924
rect 17756 4868 17812 4924
rect 17812 4868 17816 4924
rect 17752 4864 17816 4868
rect 17832 4924 17896 4928
rect 17832 4868 17836 4924
rect 17836 4868 17892 4924
rect 17892 4868 17896 4924
rect 17832 4864 17896 4868
rect 17912 4924 17976 4928
rect 17912 4868 17916 4924
rect 17916 4868 17972 4924
rect 17972 4868 17976 4924
rect 17912 4864 17976 4868
rect 17992 4924 18056 4928
rect 17992 4868 17996 4924
rect 17996 4868 18052 4924
rect 18052 4868 18056 4924
rect 17992 4864 18056 4868
rect 22552 4924 22616 4928
rect 22552 4868 22556 4924
rect 22556 4868 22612 4924
rect 22612 4868 22616 4924
rect 22552 4864 22616 4868
rect 22632 4924 22696 4928
rect 22632 4868 22636 4924
rect 22636 4868 22692 4924
rect 22692 4868 22696 4924
rect 22632 4864 22696 4868
rect 22712 4924 22776 4928
rect 22712 4868 22716 4924
rect 22716 4868 22772 4924
rect 22772 4868 22776 4924
rect 22712 4864 22776 4868
rect 22792 4924 22856 4928
rect 22792 4868 22796 4924
rect 22796 4868 22852 4924
rect 22852 4868 22856 4924
rect 22792 4864 22856 4868
rect 27352 4924 27416 4928
rect 27352 4868 27356 4924
rect 27356 4868 27412 4924
rect 27412 4868 27416 4924
rect 27352 4864 27416 4868
rect 27432 4924 27496 4928
rect 27432 4868 27436 4924
rect 27436 4868 27492 4924
rect 27492 4868 27496 4924
rect 27432 4864 27496 4868
rect 27512 4924 27576 4928
rect 27512 4868 27516 4924
rect 27516 4868 27572 4924
rect 27572 4868 27576 4924
rect 27512 4864 27576 4868
rect 27592 4924 27656 4928
rect 27592 4868 27596 4924
rect 27596 4868 27652 4924
rect 27652 4868 27656 4924
rect 27592 4864 27656 4868
rect 5752 4380 5816 4384
rect 5752 4324 5756 4380
rect 5756 4324 5812 4380
rect 5812 4324 5816 4380
rect 5752 4320 5816 4324
rect 5832 4380 5896 4384
rect 5832 4324 5836 4380
rect 5836 4324 5892 4380
rect 5892 4324 5896 4380
rect 5832 4320 5896 4324
rect 5912 4380 5976 4384
rect 5912 4324 5916 4380
rect 5916 4324 5972 4380
rect 5972 4324 5976 4380
rect 5912 4320 5976 4324
rect 5992 4380 6056 4384
rect 5992 4324 5996 4380
rect 5996 4324 6052 4380
rect 6052 4324 6056 4380
rect 5992 4320 6056 4324
rect 10552 4380 10616 4384
rect 10552 4324 10556 4380
rect 10556 4324 10612 4380
rect 10612 4324 10616 4380
rect 10552 4320 10616 4324
rect 10632 4380 10696 4384
rect 10632 4324 10636 4380
rect 10636 4324 10692 4380
rect 10692 4324 10696 4380
rect 10632 4320 10696 4324
rect 10712 4380 10776 4384
rect 10712 4324 10716 4380
rect 10716 4324 10772 4380
rect 10772 4324 10776 4380
rect 10712 4320 10776 4324
rect 10792 4380 10856 4384
rect 10792 4324 10796 4380
rect 10796 4324 10852 4380
rect 10852 4324 10856 4380
rect 10792 4320 10856 4324
rect 15352 4380 15416 4384
rect 15352 4324 15356 4380
rect 15356 4324 15412 4380
rect 15412 4324 15416 4380
rect 15352 4320 15416 4324
rect 15432 4380 15496 4384
rect 15432 4324 15436 4380
rect 15436 4324 15492 4380
rect 15492 4324 15496 4380
rect 15432 4320 15496 4324
rect 15512 4380 15576 4384
rect 15512 4324 15516 4380
rect 15516 4324 15572 4380
rect 15572 4324 15576 4380
rect 15512 4320 15576 4324
rect 15592 4380 15656 4384
rect 15592 4324 15596 4380
rect 15596 4324 15652 4380
rect 15652 4324 15656 4380
rect 15592 4320 15656 4324
rect 20152 4380 20216 4384
rect 20152 4324 20156 4380
rect 20156 4324 20212 4380
rect 20212 4324 20216 4380
rect 20152 4320 20216 4324
rect 20232 4380 20296 4384
rect 20232 4324 20236 4380
rect 20236 4324 20292 4380
rect 20292 4324 20296 4380
rect 20232 4320 20296 4324
rect 20312 4380 20376 4384
rect 20312 4324 20316 4380
rect 20316 4324 20372 4380
rect 20372 4324 20376 4380
rect 20312 4320 20376 4324
rect 20392 4380 20456 4384
rect 20392 4324 20396 4380
rect 20396 4324 20452 4380
rect 20452 4324 20456 4380
rect 20392 4320 20456 4324
rect 24952 4380 25016 4384
rect 24952 4324 24956 4380
rect 24956 4324 25012 4380
rect 25012 4324 25016 4380
rect 24952 4320 25016 4324
rect 25032 4380 25096 4384
rect 25032 4324 25036 4380
rect 25036 4324 25092 4380
rect 25092 4324 25096 4380
rect 25032 4320 25096 4324
rect 25112 4380 25176 4384
rect 25112 4324 25116 4380
rect 25116 4324 25172 4380
rect 25172 4324 25176 4380
rect 25112 4320 25176 4324
rect 25192 4380 25256 4384
rect 25192 4324 25196 4380
rect 25196 4324 25252 4380
rect 25252 4324 25256 4380
rect 25192 4320 25256 4324
rect 3352 3836 3416 3840
rect 3352 3780 3356 3836
rect 3356 3780 3412 3836
rect 3412 3780 3416 3836
rect 3352 3776 3416 3780
rect 3432 3836 3496 3840
rect 3432 3780 3436 3836
rect 3436 3780 3492 3836
rect 3492 3780 3496 3836
rect 3432 3776 3496 3780
rect 3512 3836 3576 3840
rect 3512 3780 3516 3836
rect 3516 3780 3572 3836
rect 3572 3780 3576 3836
rect 3512 3776 3576 3780
rect 3592 3836 3656 3840
rect 3592 3780 3596 3836
rect 3596 3780 3652 3836
rect 3652 3780 3656 3836
rect 3592 3776 3656 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 8312 3836 8376 3840
rect 8312 3780 8316 3836
rect 8316 3780 8372 3836
rect 8372 3780 8376 3836
rect 8312 3776 8376 3780
rect 8392 3836 8456 3840
rect 8392 3780 8396 3836
rect 8396 3780 8452 3836
rect 8452 3780 8456 3836
rect 8392 3776 8456 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 17752 3836 17816 3840
rect 17752 3780 17756 3836
rect 17756 3780 17812 3836
rect 17812 3780 17816 3836
rect 17752 3776 17816 3780
rect 17832 3836 17896 3840
rect 17832 3780 17836 3836
rect 17836 3780 17892 3836
rect 17892 3780 17896 3836
rect 17832 3776 17896 3780
rect 17912 3836 17976 3840
rect 17912 3780 17916 3836
rect 17916 3780 17972 3836
rect 17972 3780 17976 3836
rect 17912 3776 17976 3780
rect 17992 3836 18056 3840
rect 17992 3780 17996 3836
rect 17996 3780 18052 3836
rect 18052 3780 18056 3836
rect 17992 3776 18056 3780
rect 22552 3836 22616 3840
rect 22552 3780 22556 3836
rect 22556 3780 22612 3836
rect 22612 3780 22616 3836
rect 22552 3776 22616 3780
rect 22632 3836 22696 3840
rect 22632 3780 22636 3836
rect 22636 3780 22692 3836
rect 22692 3780 22696 3836
rect 22632 3776 22696 3780
rect 22712 3836 22776 3840
rect 22712 3780 22716 3836
rect 22716 3780 22772 3836
rect 22772 3780 22776 3836
rect 22712 3776 22776 3780
rect 22792 3836 22856 3840
rect 22792 3780 22796 3836
rect 22796 3780 22852 3836
rect 22852 3780 22856 3836
rect 22792 3776 22856 3780
rect 27352 3836 27416 3840
rect 27352 3780 27356 3836
rect 27356 3780 27412 3836
rect 27412 3780 27416 3836
rect 27352 3776 27416 3780
rect 27432 3836 27496 3840
rect 27432 3780 27436 3836
rect 27436 3780 27492 3836
rect 27492 3780 27496 3836
rect 27432 3776 27496 3780
rect 27512 3836 27576 3840
rect 27512 3780 27516 3836
rect 27516 3780 27572 3836
rect 27572 3780 27576 3836
rect 27512 3776 27576 3780
rect 27592 3836 27656 3840
rect 27592 3780 27596 3836
rect 27596 3780 27652 3836
rect 27652 3780 27656 3836
rect 27592 3776 27656 3780
rect 5752 3292 5816 3296
rect 5752 3236 5756 3292
rect 5756 3236 5812 3292
rect 5812 3236 5816 3292
rect 5752 3232 5816 3236
rect 5832 3292 5896 3296
rect 5832 3236 5836 3292
rect 5836 3236 5892 3292
rect 5892 3236 5896 3292
rect 5832 3232 5896 3236
rect 5912 3292 5976 3296
rect 5912 3236 5916 3292
rect 5916 3236 5972 3292
rect 5972 3236 5976 3292
rect 5912 3232 5976 3236
rect 5992 3292 6056 3296
rect 5992 3236 5996 3292
rect 5996 3236 6052 3292
rect 6052 3236 6056 3292
rect 5992 3232 6056 3236
rect 10552 3292 10616 3296
rect 10552 3236 10556 3292
rect 10556 3236 10612 3292
rect 10612 3236 10616 3292
rect 10552 3232 10616 3236
rect 10632 3292 10696 3296
rect 10632 3236 10636 3292
rect 10636 3236 10692 3292
rect 10692 3236 10696 3292
rect 10632 3232 10696 3236
rect 10712 3292 10776 3296
rect 10712 3236 10716 3292
rect 10716 3236 10772 3292
rect 10772 3236 10776 3292
rect 10712 3232 10776 3236
rect 10792 3292 10856 3296
rect 10792 3236 10796 3292
rect 10796 3236 10852 3292
rect 10852 3236 10856 3292
rect 10792 3232 10856 3236
rect 15352 3292 15416 3296
rect 15352 3236 15356 3292
rect 15356 3236 15412 3292
rect 15412 3236 15416 3292
rect 15352 3232 15416 3236
rect 15432 3292 15496 3296
rect 15432 3236 15436 3292
rect 15436 3236 15492 3292
rect 15492 3236 15496 3292
rect 15432 3232 15496 3236
rect 15512 3292 15576 3296
rect 15512 3236 15516 3292
rect 15516 3236 15572 3292
rect 15572 3236 15576 3292
rect 15512 3232 15576 3236
rect 15592 3292 15656 3296
rect 15592 3236 15596 3292
rect 15596 3236 15652 3292
rect 15652 3236 15656 3292
rect 15592 3232 15656 3236
rect 20152 3292 20216 3296
rect 20152 3236 20156 3292
rect 20156 3236 20212 3292
rect 20212 3236 20216 3292
rect 20152 3232 20216 3236
rect 20232 3292 20296 3296
rect 20232 3236 20236 3292
rect 20236 3236 20292 3292
rect 20292 3236 20296 3292
rect 20232 3232 20296 3236
rect 20312 3292 20376 3296
rect 20312 3236 20316 3292
rect 20316 3236 20372 3292
rect 20372 3236 20376 3292
rect 20312 3232 20376 3236
rect 20392 3292 20456 3296
rect 20392 3236 20396 3292
rect 20396 3236 20452 3292
rect 20452 3236 20456 3292
rect 20392 3232 20456 3236
rect 24952 3292 25016 3296
rect 24952 3236 24956 3292
rect 24956 3236 25012 3292
rect 25012 3236 25016 3292
rect 24952 3232 25016 3236
rect 25032 3292 25096 3296
rect 25032 3236 25036 3292
rect 25036 3236 25092 3292
rect 25092 3236 25096 3292
rect 25032 3232 25096 3236
rect 25112 3292 25176 3296
rect 25112 3236 25116 3292
rect 25116 3236 25172 3292
rect 25172 3236 25176 3292
rect 25112 3232 25176 3236
rect 25192 3292 25256 3296
rect 25192 3236 25196 3292
rect 25196 3236 25252 3292
rect 25252 3236 25256 3292
rect 25192 3232 25256 3236
rect 3352 2748 3416 2752
rect 3352 2692 3356 2748
rect 3356 2692 3412 2748
rect 3412 2692 3416 2748
rect 3352 2688 3416 2692
rect 3432 2748 3496 2752
rect 3432 2692 3436 2748
rect 3436 2692 3492 2748
rect 3492 2692 3496 2748
rect 3432 2688 3496 2692
rect 3512 2748 3576 2752
rect 3512 2692 3516 2748
rect 3516 2692 3572 2748
rect 3572 2692 3576 2748
rect 3512 2688 3576 2692
rect 3592 2748 3656 2752
rect 3592 2692 3596 2748
rect 3596 2692 3652 2748
rect 3652 2692 3656 2748
rect 3592 2688 3656 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 8312 2748 8376 2752
rect 8312 2692 8316 2748
rect 8316 2692 8372 2748
rect 8372 2692 8376 2748
rect 8312 2688 8376 2692
rect 8392 2748 8456 2752
rect 8392 2692 8396 2748
rect 8396 2692 8452 2748
rect 8452 2692 8456 2748
rect 8392 2688 8456 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 17752 2748 17816 2752
rect 17752 2692 17756 2748
rect 17756 2692 17812 2748
rect 17812 2692 17816 2748
rect 17752 2688 17816 2692
rect 17832 2748 17896 2752
rect 17832 2692 17836 2748
rect 17836 2692 17892 2748
rect 17892 2692 17896 2748
rect 17832 2688 17896 2692
rect 17912 2748 17976 2752
rect 17912 2692 17916 2748
rect 17916 2692 17972 2748
rect 17972 2692 17976 2748
rect 17912 2688 17976 2692
rect 17992 2748 18056 2752
rect 17992 2692 17996 2748
rect 17996 2692 18052 2748
rect 18052 2692 18056 2748
rect 17992 2688 18056 2692
rect 22552 2748 22616 2752
rect 22552 2692 22556 2748
rect 22556 2692 22612 2748
rect 22612 2692 22616 2748
rect 22552 2688 22616 2692
rect 22632 2748 22696 2752
rect 22632 2692 22636 2748
rect 22636 2692 22692 2748
rect 22692 2692 22696 2748
rect 22632 2688 22696 2692
rect 22712 2748 22776 2752
rect 22712 2692 22716 2748
rect 22716 2692 22772 2748
rect 22772 2692 22776 2748
rect 22712 2688 22776 2692
rect 22792 2748 22856 2752
rect 22792 2692 22796 2748
rect 22796 2692 22852 2748
rect 22852 2692 22856 2748
rect 22792 2688 22856 2692
rect 27352 2748 27416 2752
rect 27352 2692 27356 2748
rect 27356 2692 27412 2748
rect 27412 2692 27416 2748
rect 27352 2688 27416 2692
rect 27432 2748 27496 2752
rect 27432 2692 27436 2748
rect 27436 2692 27492 2748
rect 27492 2692 27496 2748
rect 27432 2688 27496 2692
rect 27512 2748 27576 2752
rect 27512 2692 27516 2748
rect 27516 2692 27572 2748
rect 27572 2692 27576 2748
rect 27512 2688 27576 2692
rect 27592 2748 27656 2752
rect 27592 2692 27596 2748
rect 27596 2692 27652 2748
rect 27652 2692 27656 2748
rect 27592 2688 27656 2692
rect 5752 2204 5816 2208
rect 5752 2148 5756 2204
rect 5756 2148 5812 2204
rect 5812 2148 5816 2204
rect 5752 2144 5816 2148
rect 5832 2204 5896 2208
rect 5832 2148 5836 2204
rect 5836 2148 5892 2204
rect 5892 2148 5896 2204
rect 5832 2144 5896 2148
rect 5912 2204 5976 2208
rect 5912 2148 5916 2204
rect 5916 2148 5972 2204
rect 5972 2148 5976 2204
rect 5912 2144 5976 2148
rect 5992 2204 6056 2208
rect 5992 2148 5996 2204
rect 5996 2148 6052 2204
rect 6052 2148 6056 2204
rect 5992 2144 6056 2148
rect 10552 2204 10616 2208
rect 10552 2148 10556 2204
rect 10556 2148 10612 2204
rect 10612 2148 10616 2204
rect 10552 2144 10616 2148
rect 10632 2204 10696 2208
rect 10632 2148 10636 2204
rect 10636 2148 10692 2204
rect 10692 2148 10696 2204
rect 10632 2144 10696 2148
rect 10712 2204 10776 2208
rect 10712 2148 10716 2204
rect 10716 2148 10772 2204
rect 10772 2148 10776 2204
rect 10712 2144 10776 2148
rect 10792 2204 10856 2208
rect 10792 2148 10796 2204
rect 10796 2148 10852 2204
rect 10852 2148 10856 2204
rect 10792 2144 10856 2148
rect 15352 2204 15416 2208
rect 15352 2148 15356 2204
rect 15356 2148 15412 2204
rect 15412 2148 15416 2204
rect 15352 2144 15416 2148
rect 15432 2204 15496 2208
rect 15432 2148 15436 2204
rect 15436 2148 15492 2204
rect 15492 2148 15496 2204
rect 15432 2144 15496 2148
rect 15512 2204 15576 2208
rect 15512 2148 15516 2204
rect 15516 2148 15572 2204
rect 15572 2148 15576 2204
rect 15512 2144 15576 2148
rect 15592 2204 15656 2208
rect 15592 2148 15596 2204
rect 15596 2148 15652 2204
rect 15652 2148 15656 2204
rect 15592 2144 15656 2148
rect 20152 2204 20216 2208
rect 20152 2148 20156 2204
rect 20156 2148 20212 2204
rect 20212 2148 20216 2204
rect 20152 2144 20216 2148
rect 20232 2204 20296 2208
rect 20232 2148 20236 2204
rect 20236 2148 20292 2204
rect 20292 2148 20296 2204
rect 20232 2144 20296 2148
rect 20312 2204 20376 2208
rect 20312 2148 20316 2204
rect 20316 2148 20372 2204
rect 20372 2148 20376 2204
rect 20312 2144 20376 2148
rect 20392 2204 20456 2208
rect 20392 2148 20396 2204
rect 20396 2148 20452 2204
rect 20452 2148 20456 2204
rect 20392 2144 20456 2148
rect 24952 2204 25016 2208
rect 24952 2148 24956 2204
rect 24956 2148 25012 2204
rect 25012 2148 25016 2204
rect 24952 2144 25016 2148
rect 25032 2204 25096 2208
rect 25032 2148 25036 2204
rect 25036 2148 25092 2204
rect 25092 2148 25096 2204
rect 25032 2144 25096 2148
rect 25112 2204 25176 2208
rect 25112 2148 25116 2204
rect 25116 2148 25172 2204
rect 25172 2148 25176 2204
rect 25112 2144 25176 2148
rect 25192 2204 25256 2208
rect 25192 2148 25196 2204
rect 25196 2148 25252 2204
rect 25252 2148 25256 2204
rect 25192 2144 25256 2148
<< metal4 >>
rect 3344 27776 3664 27792
rect 3344 27712 3352 27776
rect 3416 27712 3432 27776
rect 3496 27712 3512 27776
rect 3576 27712 3592 27776
rect 3656 27712 3664 27776
rect 3344 26688 3664 27712
rect 3344 26624 3352 26688
rect 3416 26624 3432 26688
rect 3496 26624 3512 26688
rect 3576 26624 3592 26688
rect 3656 26624 3664 26688
rect 3344 25600 3664 26624
rect 3344 25536 3352 25600
rect 3416 25536 3432 25600
rect 3496 25536 3512 25600
rect 3576 25536 3592 25600
rect 3656 25536 3664 25600
rect 3344 24512 3664 25536
rect 3344 24448 3352 24512
rect 3416 24448 3432 24512
rect 3496 24448 3512 24512
rect 3576 24448 3592 24512
rect 3656 24448 3664 24512
rect 3344 23424 3664 24448
rect 3344 23360 3352 23424
rect 3416 23360 3432 23424
rect 3496 23360 3512 23424
rect 3576 23360 3592 23424
rect 3656 23360 3664 23424
rect 3344 22336 3664 23360
rect 3344 22272 3352 22336
rect 3416 22272 3432 22336
rect 3496 22272 3512 22336
rect 3576 22272 3592 22336
rect 3656 22272 3664 22336
rect 3344 21248 3664 22272
rect 3344 21184 3352 21248
rect 3416 21184 3432 21248
rect 3496 21184 3512 21248
rect 3576 21184 3592 21248
rect 3656 21184 3664 21248
rect 3344 20160 3664 21184
rect 3344 20096 3352 20160
rect 3416 20096 3432 20160
rect 3496 20096 3512 20160
rect 3576 20096 3592 20160
rect 3656 20096 3664 20160
rect 3344 19072 3664 20096
rect 3344 19008 3352 19072
rect 3416 19008 3432 19072
rect 3496 19008 3512 19072
rect 3576 19008 3592 19072
rect 3656 19008 3664 19072
rect 3344 17984 3664 19008
rect 3344 17920 3352 17984
rect 3416 17920 3432 17984
rect 3496 17920 3512 17984
rect 3576 17920 3592 17984
rect 3656 17920 3664 17984
rect 3344 16896 3664 17920
rect 3344 16832 3352 16896
rect 3416 16832 3432 16896
rect 3496 16832 3512 16896
rect 3576 16832 3592 16896
rect 3656 16832 3664 16896
rect 3344 15808 3664 16832
rect 3344 15744 3352 15808
rect 3416 15744 3432 15808
rect 3496 15744 3512 15808
rect 3576 15744 3592 15808
rect 3656 15744 3664 15808
rect 3344 14720 3664 15744
rect 3344 14656 3352 14720
rect 3416 14656 3432 14720
rect 3496 14656 3512 14720
rect 3576 14656 3592 14720
rect 3656 14656 3664 14720
rect 3344 13632 3664 14656
rect 3344 13568 3352 13632
rect 3416 13568 3432 13632
rect 3496 13568 3512 13632
rect 3576 13568 3592 13632
rect 3656 13568 3664 13632
rect 3344 12544 3664 13568
rect 3344 12480 3352 12544
rect 3416 12480 3432 12544
rect 3496 12480 3512 12544
rect 3576 12480 3592 12544
rect 3656 12480 3664 12544
rect 3344 11456 3664 12480
rect 3344 11392 3352 11456
rect 3416 11392 3432 11456
rect 3496 11392 3512 11456
rect 3576 11392 3592 11456
rect 3656 11392 3664 11456
rect 3344 10368 3664 11392
rect 3344 10304 3352 10368
rect 3416 10304 3432 10368
rect 3496 10304 3512 10368
rect 3576 10304 3592 10368
rect 3656 10304 3664 10368
rect 3344 9280 3664 10304
rect 3344 9216 3352 9280
rect 3416 9216 3432 9280
rect 3496 9216 3512 9280
rect 3576 9216 3592 9280
rect 3656 9216 3664 9280
rect 3344 8192 3664 9216
rect 3344 8128 3352 8192
rect 3416 8128 3432 8192
rect 3496 8128 3512 8192
rect 3576 8128 3592 8192
rect 3656 8128 3664 8192
rect 3344 7104 3664 8128
rect 3344 7040 3352 7104
rect 3416 7040 3432 7104
rect 3496 7040 3512 7104
rect 3576 7040 3592 7104
rect 3656 7040 3664 7104
rect 3344 6016 3664 7040
rect 3344 5952 3352 6016
rect 3416 5952 3432 6016
rect 3496 5952 3512 6016
rect 3576 5952 3592 6016
rect 3656 5952 3664 6016
rect 3344 4928 3664 5952
rect 3344 4864 3352 4928
rect 3416 4864 3432 4928
rect 3496 4864 3512 4928
rect 3576 4864 3592 4928
rect 3656 4864 3664 4928
rect 3344 3840 3664 4864
rect 3344 3776 3352 3840
rect 3416 3776 3432 3840
rect 3496 3776 3512 3840
rect 3576 3776 3592 3840
rect 3656 3776 3664 3840
rect 3344 2752 3664 3776
rect 3344 2688 3352 2752
rect 3416 2688 3432 2752
rect 3496 2688 3512 2752
rect 3576 2688 3592 2752
rect 3656 2688 3664 2752
rect 3344 2128 3664 2688
rect 5744 27232 6064 27792
rect 5744 27168 5752 27232
rect 5816 27168 5832 27232
rect 5896 27168 5912 27232
rect 5976 27168 5992 27232
rect 6056 27168 6064 27232
rect 5744 26144 6064 27168
rect 5744 26080 5752 26144
rect 5816 26080 5832 26144
rect 5896 26080 5912 26144
rect 5976 26080 5992 26144
rect 6056 26080 6064 26144
rect 5744 25056 6064 26080
rect 5744 24992 5752 25056
rect 5816 24992 5832 25056
rect 5896 24992 5912 25056
rect 5976 24992 5992 25056
rect 6056 24992 6064 25056
rect 5744 23968 6064 24992
rect 5744 23904 5752 23968
rect 5816 23904 5832 23968
rect 5896 23904 5912 23968
rect 5976 23904 5992 23968
rect 6056 23904 6064 23968
rect 5744 22880 6064 23904
rect 5744 22816 5752 22880
rect 5816 22816 5832 22880
rect 5896 22816 5912 22880
rect 5976 22816 5992 22880
rect 6056 22816 6064 22880
rect 5744 21792 6064 22816
rect 5744 21728 5752 21792
rect 5816 21728 5832 21792
rect 5896 21728 5912 21792
rect 5976 21728 5992 21792
rect 6056 21728 6064 21792
rect 5744 20704 6064 21728
rect 5744 20640 5752 20704
rect 5816 20640 5832 20704
rect 5896 20640 5912 20704
rect 5976 20640 5992 20704
rect 6056 20640 6064 20704
rect 5744 19616 6064 20640
rect 5744 19552 5752 19616
rect 5816 19552 5832 19616
rect 5896 19552 5912 19616
rect 5976 19552 5992 19616
rect 6056 19552 6064 19616
rect 5744 18528 6064 19552
rect 5744 18464 5752 18528
rect 5816 18464 5832 18528
rect 5896 18464 5912 18528
rect 5976 18464 5992 18528
rect 6056 18464 6064 18528
rect 5744 17440 6064 18464
rect 5744 17376 5752 17440
rect 5816 17376 5832 17440
rect 5896 17376 5912 17440
rect 5976 17376 5992 17440
rect 6056 17376 6064 17440
rect 5744 16352 6064 17376
rect 5744 16288 5752 16352
rect 5816 16288 5832 16352
rect 5896 16288 5912 16352
rect 5976 16288 5992 16352
rect 6056 16288 6064 16352
rect 5744 15264 6064 16288
rect 5744 15200 5752 15264
rect 5816 15200 5832 15264
rect 5896 15200 5912 15264
rect 5976 15200 5992 15264
rect 6056 15200 6064 15264
rect 5744 14176 6064 15200
rect 5744 14112 5752 14176
rect 5816 14112 5832 14176
rect 5896 14112 5912 14176
rect 5976 14112 5992 14176
rect 6056 14112 6064 14176
rect 5744 13088 6064 14112
rect 5744 13024 5752 13088
rect 5816 13024 5832 13088
rect 5896 13024 5912 13088
rect 5976 13024 5992 13088
rect 6056 13024 6064 13088
rect 5744 12000 6064 13024
rect 5744 11936 5752 12000
rect 5816 11936 5832 12000
rect 5896 11936 5912 12000
rect 5976 11936 5992 12000
rect 6056 11936 6064 12000
rect 5744 10912 6064 11936
rect 5744 10848 5752 10912
rect 5816 10848 5832 10912
rect 5896 10848 5912 10912
rect 5976 10848 5992 10912
rect 6056 10848 6064 10912
rect 5744 9824 6064 10848
rect 5744 9760 5752 9824
rect 5816 9760 5832 9824
rect 5896 9760 5912 9824
rect 5976 9760 5992 9824
rect 6056 9760 6064 9824
rect 5744 8736 6064 9760
rect 5744 8672 5752 8736
rect 5816 8672 5832 8736
rect 5896 8672 5912 8736
rect 5976 8672 5992 8736
rect 6056 8672 6064 8736
rect 5744 7648 6064 8672
rect 5744 7584 5752 7648
rect 5816 7584 5832 7648
rect 5896 7584 5912 7648
rect 5976 7584 5992 7648
rect 6056 7584 6064 7648
rect 5744 6560 6064 7584
rect 5744 6496 5752 6560
rect 5816 6496 5832 6560
rect 5896 6496 5912 6560
rect 5976 6496 5992 6560
rect 6056 6496 6064 6560
rect 5744 5472 6064 6496
rect 5744 5408 5752 5472
rect 5816 5408 5832 5472
rect 5896 5408 5912 5472
rect 5976 5408 5992 5472
rect 6056 5408 6064 5472
rect 5744 4384 6064 5408
rect 5744 4320 5752 4384
rect 5816 4320 5832 4384
rect 5896 4320 5912 4384
rect 5976 4320 5992 4384
rect 6056 4320 6064 4384
rect 5744 3296 6064 4320
rect 5744 3232 5752 3296
rect 5816 3232 5832 3296
rect 5896 3232 5912 3296
rect 5976 3232 5992 3296
rect 6056 3232 6064 3296
rect 5744 2208 6064 3232
rect 5744 2144 5752 2208
rect 5816 2144 5832 2208
rect 5896 2144 5912 2208
rect 5976 2144 5992 2208
rect 6056 2144 6064 2208
rect 5744 2128 6064 2144
rect 8144 27776 8464 27792
rect 8144 27712 8152 27776
rect 8216 27712 8232 27776
rect 8296 27712 8312 27776
rect 8376 27712 8392 27776
rect 8456 27712 8464 27776
rect 8144 26688 8464 27712
rect 8144 26624 8152 26688
rect 8216 26624 8232 26688
rect 8296 26624 8312 26688
rect 8376 26624 8392 26688
rect 8456 26624 8464 26688
rect 8144 25600 8464 26624
rect 8144 25536 8152 25600
rect 8216 25536 8232 25600
rect 8296 25536 8312 25600
rect 8376 25536 8392 25600
rect 8456 25536 8464 25600
rect 8144 24512 8464 25536
rect 8144 24448 8152 24512
rect 8216 24448 8232 24512
rect 8296 24448 8312 24512
rect 8376 24448 8392 24512
rect 8456 24448 8464 24512
rect 8144 23424 8464 24448
rect 8144 23360 8152 23424
rect 8216 23360 8232 23424
rect 8296 23360 8312 23424
rect 8376 23360 8392 23424
rect 8456 23360 8464 23424
rect 8144 22336 8464 23360
rect 8144 22272 8152 22336
rect 8216 22272 8232 22336
rect 8296 22272 8312 22336
rect 8376 22272 8392 22336
rect 8456 22272 8464 22336
rect 8144 21248 8464 22272
rect 8144 21184 8152 21248
rect 8216 21184 8232 21248
rect 8296 21184 8312 21248
rect 8376 21184 8392 21248
rect 8456 21184 8464 21248
rect 8144 20160 8464 21184
rect 8144 20096 8152 20160
rect 8216 20096 8232 20160
rect 8296 20096 8312 20160
rect 8376 20096 8392 20160
rect 8456 20096 8464 20160
rect 8144 19072 8464 20096
rect 8144 19008 8152 19072
rect 8216 19008 8232 19072
rect 8296 19008 8312 19072
rect 8376 19008 8392 19072
rect 8456 19008 8464 19072
rect 8144 17984 8464 19008
rect 8144 17920 8152 17984
rect 8216 17920 8232 17984
rect 8296 17920 8312 17984
rect 8376 17920 8392 17984
rect 8456 17920 8464 17984
rect 8144 16896 8464 17920
rect 8144 16832 8152 16896
rect 8216 16832 8232 16896
rect 8296 16832 8312 16896
rect 8376 16832 8392 16896
rect 8456 16832 8464 16896
rect 8144 15808 8464 16832
rect 8144 15744 8152 15808
rect 8216 15744 8232 15808
rect 8296 15744 8312 15808
rect 8376 15744 8392 15808
rect 8456 15744 8464 15808
rect 8144 14720 8464 15744
rect 8144 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8312 14720
rect 8376 14656 8392 14720
rect 8456 14656 8464 14720
rect 8144 13632 8464 14656
rect 8144 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8312 13632
rect 8376 13568 8392 13632
rect 8456 13568 8464 13632
rect 8144 12544 8464 13568
rect 8144 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8312 12544
rect 8376 12480 8392 12544
rect 8456 12480 8464 12544
rect 8144 11456 8464 12480
rect 8144 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8312 11456
rect 8376 11392 8392 11456
rect 8456 11392 8464 11456
rect 8144 10368 8464 11392
rect 8144 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8312 10368
rect 8376 10304 8392 10368
rect 8456 10304 8464 10368
rect 8144 9280 8464 10304
rect 8144 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8312 9280
rect 8376 9216 8392 9280
rect 8456 9216 8464 9280
rect 8144 8192 8464 9216
rect 8144 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8312 8192
rect 8376 8128 8392 8192
rect 8456 8128 8464 8192
rect 8144 7104 8464 8128
rect 8144 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8312 7104
rect 8376 7040 8392 7104
rect 8456 7040 8464 7104
rect 8144 6016 8464 7040
rect 8144 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8312 6016
rect 8376 5952 8392 6016
rect 8456 5952 8464 6016
rect 8144 4928 8464 5952
rect 8144 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8312 4928
rect 8376 4864 8392 4928
rect 8456 4864 8464 4928
rect 8144 3840 8464 4864
rect 8144 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8312 3840
rect 8376 3776 8392 3840
rect 8456 3776 8464 3840
rect 8144 2752 8464 3776
rect 8144 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8312 2752
rect 8376 2688 8392 2752
rect 8456 2688 8464 2752
rect 8144 2128 8464 2688
rect 10544 27232 10864 27792
rect 10544 27168 10552 27232
rect 10616 27168 10632 27232
rect 10696 27168 10712 27232
rect 10776 27168 10792 27232
rect 10856 27168 10864 27232
rect 10544 26144 10864 27168
rect 10544 26080 10552 26144
rect 10616 26080 10632 26144
rect 10696 26080 10712 26144
rect 10776 26080 10792 26144
rect 10856 26080 10864 26144
rect 10544 25056 10864 26080
rect 10544 24992 10552 25056
rect 10616 24992 10632 25056
rect 10696 24992 10712 25056
rect 10776 24992 10792 25056
rect 10856 24992 10864 25056
rect 10544 23968 10864 24992
rect 10544 23904 10552 23968
rect 10616 23904 10632 23968
rect 10696 23904 10712 23968
rect 10776 23904 10792 23968
rect 10856 23904 10864 23968
rect 10544 22880 10864 23904
rect 10544 22816 10552 22880
rect 10616 22816 10632 22880
rect 10696 22816 10712 22880
rect 10776 22816 10792 22880
rect 10856 22816 10864 22880
rect 10544 21792 10864 22816
rect 10544 21728 10552 21792
rect 10616 21728 10632 21792
rect 10696 21728 10712 21792
rect 10776 21728 10792 21792
rect 10856 21728 10864 21792
rect 10544 20704 10864 21728
rect 10544 20640 10552 20704
rect 10616 20640 10632 20704
rect 10696 20640 10712 20704
rect 10776 20640 10792 20704
rect 10856 20640 10864 20704
rect 10544 19616 10864 20640
rect 10544 19552 10552 19616
rect 10616 19552 10632 19616
rect 10696 19552 10712 19616
rect 10776 19552 10792 19616
rect 10856 19552 10864 19616
rect 10544 18528 10864 19552
rect 10544 18464 10552 18528
rect 10616 18464 10632 18528
rect 10696 18464 10712 18528
rect 10776 18464 10792 18528
rect 10856 18464 10864 18528
rect 10544 17440 10864 18464
rect 10544 17376 10552 17440
rect 10616 17376 10632 17440
rect 10696 17376 10712 17440
rect 10776 17376 10792 17440
rect 10856 17376 10864 17440
rect 10544 16352 10864 17376
rect 10544 16288 10552 16352
rect 10616 16288 10632 16352
rect 10696 16288 10712 16352
rect 10776 16288 10792 16352
rect 10856 16288 10864 16352
rect 10544 15264 10864 16288
rect 10544 15200 10552 15264
rect 10616 15200 10632 15264
rect 10696 15200 10712 15264
rect 10776 15200 10792 15264
rect 10856 15200 10864 15264
rect 10544 14176 10864 15200
rect 10544 14112 10552 14176
rect 10616 14112 10632 14176
rect 10696 14112 10712 14176
rect 10776 14112 10792 14176
rect 10856 14112 10864 14176
rect 10544 13088 10864 14112
rect 10544 13024 10552 13088
rect 10616 13024 10632 13088
rect 10696 13024 10712 13088
rect 10776 13024 10792 13088
rect 10856 13024 10864 13088
rect 10544 12000 10864 13024
rect 10544 11936 10552 12000
rect 10616 11936 10632 12000
rect 10696 11936 10712 12000
rect 10776 11936 10792 12000
rect 10856 11936 10864 12000
rect 10544 10912 10864 11936
rect 10544 10848 10552 10912
rect 10616 10848 10632 10912
rect 10696 10848 10712 10912
rect 10776 10848 10792 10912
rect 10856 10848 10864 10912
rect 10544 9824 10864 10848
rect 10544 9760 10552 9824
rect 10616 9760 10632 9824
rect 10696 9760 10712 9824
rect 10776 9760 10792 9824
rect 10856 9760 10864 9824
rect 10544 8736 10864 9760
rect 10544 8672 10552 8736
rect 10616 8672 10632 8736
rect 10696 8672 10712 8736
rect 10776 8672 10792 8736
rect 10856 8672 10864 8736
rect 10544 7648 10864 8672
rect 10544 7584 10552 7648
rect 10616 7584 10632 7648
rect 10696 7584 10712 7648
rect 10776 7584 10792 7648
rect 10856 7584 10864 7648
rect 10544 6560 10864 7584
rect 10544 6496 10552 6560
rect 10616 6496 10632 6560
rect 10696 6496 10712 6560
rect 10776 6496 10792 6560
rect 10856 6496 10864 6560
rect 10544 5472 10864 6496
rect 10544 5408 10552 5472
rect 10616 5408 10632 5472
rect 10696 5408 10712 5472
rect 10776 5408 10792 5472
rect 10856 5408 10864 5472
rect 10544 4384 10864 5408
rect 10544 4320 10552 4384
rect 10616 4320 10632 4384
rect 10696 4320 10712 4384
rect 10776 4320 10792 4384
rect 10856 4320 10864 4384
rect 10544 3296 10864 4320
rect 10544 3232 10552 3296
rect 10616 3232 10632 3296
rect 10696 3232 10712 3296
rect 10776 3232 10792 3296
rect 10856 3232 10864 3296
rect 10544 2208 10864 3232
rect 10544 2144 10552 2208
rect 10616 2144 10632 2208
rect 10696 2144 10712 2208
rect 10776 2144 10792 2208
rect 10856 2144 10864 2208
rect 10544 2128 10864 2144
rect 12944 27776 13264 27792
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 15344 27232 15664 27792
rect 15344 27168 15352 27232
rect 15416 27168 15432 27232
rect 15496 27168 15512 27232
rect 15576 27168 15592 27232
rect 15656 27168 15664 27232
rect 15344 26144 15664 27168
rect 15344 26080 15352 26144
rect 15416 26080 15432 26144
rect 15496 26080 15512 26144
rect 15576 26080 15592 26144
rect 15656 26080 15664 26144
rect 15344 25056 15664 26080
rect 15344 24992 15352 25056
rect 15416 24992 15432 25056
rect 15496 24992 15512 25056
rect 15576 24992 15592 25056
rect 15656 24992 15664 25056
rect 15344 23968 15664 24992
rect 15344 23904 15352 23968
rect 15416 23904 15432 23968
rect 15496 23904 15512 23968
rect 15576 23904 15592 23968
rect 15656 23904 15664 23968
rect 15344 22880 15664 23904
rect 15344 22816 15352 22880
rect 15416 22816 15432 22880
rect 15496 22816 15512 22880
rect 15576 22816 15592 22880
rect 15656 22816 15664 22880
rect 15344 21792 15664 22816
rect 15344 21728 15352 21792
rect 15416 21728 15432 21792
rect 15496 21728 15512 21792
rect 15576 21728 15592 21792
rect 15656 21728 15664 21792
rect 15344 20704 15664 21728
rect 15344 20640 15352 20704
rect 15416 20640 15432 20704
rect 15496 20640 15512 20704
rect 15576 20640 15592 20704
rect 15656 20640 15664 20704
rect 15344 19616 15664 20640
rect 15344 19552 15352 19616
rect 15416 19552 15432 19616
rect 15496 19552 15512 19616
rect 15576 19552 15592 19616
rect 15656 19552 15664 19616
rect 15344 18528 15664 19552
rect 15344 18464 15352 18528
rect 15416 18464 15432 18528
rect 15496 18464 15512 18528
rect 15576 18464 15592 18528
rect 15656 18464 15664 18528
rect 15344 17440 15664 18464
rect 15344 17376 15352 17440
rect 15416 17376 15432 17440
rect 15496 17376 15512 17440
rect 15576 17376 15592 17440
rect 15656 17376 15664 17440
rect 15344 16352 15664 17376
rect 15344 16288 15352 16352
rect 15416 16288 15432 16352
rect 15496 16288 15512 16352
rect 15576 16288 15592 16352
rect 15656 16288 15664 16352
rect 15344 15264 15664 16288
rect 15344 15200 15352 15264
rect 15416 15200 15432 15264
rect 15496 15200 15512 15264
rect 15576 15200 15592 15264
rect 15656 15200 15664 15264
rect 15344 14176 15664 15200
rect 15344 14112 15352 14176
rect 15416 14112 15432 14176
rect 15496 14112 15512 14176
rect 15576 14112 15592 14176
rect 15656 14112 15664 14176
rect 15344 13088 15664 14112
rect 15344 13024 15352 13088
rect 15416 13024 15432 13088
rect 15496 13024 15512 13088
rect 15576 13024 15592 13088
rect 15656 13024 15664 13088
rect 15344 12000 15664 13024
rect 15344 11936 15352 12000
rect 15416 11936 15432 12000
rect 15496 11936 15512 12000
rect 15576 11936 15592 12000
rect 15656 11936 15664 12000
rect 15344 10912 15664 11936
rect 15344 10848 15352 10912
rect 15416 10848 15432 10912
rect 15496 10848 15512 10912
rect 15576 10848 15592 10912
rect 15656 10848 15664 10912
rect 15344 9824 15664 10848
rect 15344 9760 15352 9824
rect 15416 9760 15432 9824
rect 15496 9760 15512 9824
rect 15576 9760 15592 9824
rect 15656 9760 15664 9824
rect 15344 8736 15664 9760
rect 15344 8672 15352 8736
rect 15416 8672 15432 8736
rect 15496 8672 15512 8736
rect 15576 8672 15592 8736
rect 15656 8672 15664 8736
rect 15344 7648 15664 8672
rect 15344 7584 15352 7648
rect 15416 7584 15432 7648
rect 15496 7584 15512 7648
rect 15576 7584 15592 7648
rect 15656 7584 15664 7648
rect 15344 6560 15664 7584
rect 15344 6496 15352 6560
rect 15416 6496 15432 6560
rect 15496 6496 15512 6560
rect 15576 6496 15592 6560
rect 15656 6496 15664 6560
rect 15344 5472 15664 6496
rect 15344 5408 15352 5472
rect 15416 5408 15432 5472
rect 15496 5408 15512 5472
rect 15576 5408 15592 5472
rect 15656 5408 15664 5472
rect 15344 4384 15664 5408
rect 15344 4320 15352 4384
rect 15416 4320 15432 4384
rect 15496 4320 15512 4384
rect 15576 4320 15592 4384
rect 15656 4320 15664 4384
rect 15344 3296 15664 4320
rect 15344 3232 15352 3296
rect 15416 3232 15432 3296
rect 15496 3232 15512 3296
rect 15576 3232 15592 3296
rect 15656 3232 15664 3296
rect 15344 2208 15664 3232
rect 15344 2144 15352 2208
rect 15416 2144 15432 2208
rect 15496 2144 15512 2208
rect 15576 2144 15592 2208
rect 15656 2144 15664 2208
rect 15344 2128 15664 2144
rect 17744 27776 18064 27792
rect 17744 27712 17752 27776
rect 17816 27712 17832 27776
rect 17896 27712 17912 27776
rect 17976 27712 17992 27776
rect 18056 27712 18064 27776
rect 17744 26688 18064 27712
rect 17744 26624 17752 26688
rect 17816 26624 17832 26688
rect 17896 26624 17912 26688
rect 17976 26624 17992 26688
rect 18056 26624 18064 26688
rect 17744 25600 18064 26624
rect 17744 25536 17752 25600
rect 17816 25536 17832 25600
rect 17896 25536 17912 25600
rect 17976 25536 17992 25600
rect 18056 25536 18064 25600
rect 17744 24512 18064 25536
rect 17744 24448 17752 24512
rect 17816 24448 17832 24512
rect 17896 24448 17912 24512
rect 17976 24448 17992 24512
rect 18056 24448 18064 24512
rect 17744 23424 18064 24448
rect 17744 23360 17752 23424
rect 17816 23360 17832 23424
rect 17896 23360 17912 23424
rect 17976 23360 17992 23424
rect 18056 23360 18064 23424
rect 17744 22336 18064 23360
rect 17744 22272 17752 22336
rect 17816 22272 17832 22336
rect 17896 22272 17912 22336
rect 17976 22272 17992 22336
rect 18056 22272 18064 22336
rect 17744 21248 18064 22272
rect 17744 21184 17752 21248
rect 17816 21184 17832 21248
rect 17896 21184 17912 21248
rect 17976 21184 17992 21248
rect 18056 21184 18064 21248
rect 17744 20160 18064 21184
rect 17744 20096 17752 20160
rect 17816 20096 17832 20160
rect 17896 20096 17912 20160
rect 17976 20096 17992 20160
rect 18056 20096 18064 20160
rect 17744 19072 18064 20096
rect 17744 19008 17752 19072
rect 17816 19008 17832 19072
rect 17896 19008 17912 19072
rect 17976 19008 17992 19072
rect 18056 19008 18064 19072
rect 17744 17984 18064 19008
rect 17744 17920 17752 17984
rect 17816 17920 17832 17984
rect 17896 17920 17912 17984
rect 17976 17920 17992 17984
rect 18056 17920 18064 17984
rect 17744 16896 18064 17920
rect 17744 16832 17752 16896
rect 17816 16832 17832 16896
rect 17896 16832 17912 16896
rect 17976 16832 17992 16896
rect 18056 16832 18064 16896
rect 17744 15808 18064 16832
rect 17744 15744 17752 15808
rect 17816 15744 17832 15808
rect 17896 15744 17912 15808
rect 17976 15744 17992 15808
rect 18056 15744 18064 15808
rect 17744 14720 18064 15744
rect 17744 14656 17752 14720
rect 17816 14656 17832 14720
rect 17896 14656 17912 14720
rect 17976 14656 17992 14720
rect 18056 14656 18064 14720
rect 17744 13632 18064 14656
rect 17744 13568 17752 13632
rect 17816 13568 17832 13632
rect 17896 13568 17912 13632
rect 17976 13568 17992 13632
rect 18056 13568 18064 13632
rect 17744 12544 18064 13568
rect 17744 12480 17752 12544
rect 17816 12480 17832 12544
rect 17896 12480 17912 12544
rect 17976 12480 17992 12544
rect 18056 12480 18064 12544
rect 17744 11456 18064 12480
rect 17744 11392 17752 11456
rect 17816 11392 17832 11456
rect 17896 11392 17912 11456
rect 17976 11392 17992 11456
rect 18056 11392 18064 11456
rect 17744 10368 18064 11392
rect 17744 10304 17752 10368
rect 17816 10304 17832 10368
rect 17896 10304 17912 10368
rect 17976 10304 17992 10368
rect 18056 10304 18064 10368
rect 17744 9280 18064 10304
rect 17744 9216 17752 9280
rect 17816 9216 17832 9280
rect 17896 9216 17912 9280
rect 17976 9216 17992 9280
rect 18056 9216 18064 9280
rect 17744 8192 18064 9216
rect 17744 8128 17752 8192
rect 17816 8128 17832 8192
rect 17896 8128 17912 8192
rect 17976 8128 17992 8192
rect 18056 8128 18064 8192
rect 17744 7104 18064 8128
rect 17744 7040 17752 7104
rect 17816 7040 17832 7104
rect 17896 7040 17912 7104
rect 17976 7040 17992 7104
rect 18056 7040 18064 7104
rect 17744 6016 18064 7040
rect 17744 5952 17752 6016
rect 17816 5952 17832 6016
rect 17896 5952 17912 6016
rect 17976 5952 17992 6016
rect 18056 5952 18064 6016
rect 17744 4928 18064 5952
rect 17744 4864 17752 4928
rect 17816 4864 17832 4928
rect 17896 4864 17912 4928
rect 17976 4864 17992 4928
rect 18056 4864 18064 4928
rect 17744 3840 18064 4864
rect 17744 3776 17752 3840
rect 17816 3776 17832 3840
rect 17896 3776 17912 3840
rect 17976 3776 17992 3840
rect 18056 3776 18064 3840
rect 17744 2752 18064 3776
rect 17744 2688 17752 2752
rect 17816 2688 17832 2752
rect 17896 2688 17912 2752
rect 17976 2688 17992 2752
rect 18056 2688 18064 2752
rect 17744 2128 18064 2688
rect 20144 27232 20464 27792
rect 20144 27168 20152 27232
rect 20216 27168 20232 27232
rect 20296 27168 20312 27232
rect 20376 27168 20392 27232
rect 20456 27168 20464 27232
rect 20144 26144 20464 27168
rect 20144 26080 20152 26144
rect 20216 26080 20232 26144
rect 20296 26080 20312 26144
rect 20376 26080 20392 26144
rect 20456 26080 20464 26144
rect 20144 25056 20464 26080
rect 20144 24992 20152 25056
rect 20216 24992 20232 25056
rect 20296 24992 20312 25056
rect 20376 24992 20392 25056
rect 20456 24992 20464 25056
rect 20144 23968 20464 24992
rect 20144 23904 20152 23968
rect 20216 23904 20232 23968
rect 20296 23904 20312 23968
rect 20376 23904 20392 23968
rect 20456 23904 20464 23968
rect 20144 22880 20464 23904
rect 20144 22816 20152 22880
rect 20216 22816 20232 22880
rect 20296 22816 20312 22880
rect 20376 22816 20392 22880
rect 20456 22816 20464 22880
rect 20144 21792 20464 22816
rect 20144 21728 20152 21792
rect 20216 21728 20232 21792
rect 20296 21728 20312 21792
rect 20376 21728 20392 21792
rect 20456 21728 20464 21792
rect 20144 20704 20464 21728
rect 20144 20640 20152 20704
rect 20216 20640 20232 20704
rect 20296 20640 20312 20704
rect 20376 20640 20392 20704
rect 20456 20640 20464 20704
rect 20144 19616 20464 20640
rect 20144 19552 20152 19616
rect 20216 19552 20232 19616
rect 20296 19552 20312 19616
rect 20376 19552 20392 19616
rect 20456 19552 20464 19616
rect 20144 18528 20464 19552
rect 20144 18464 20152 18528
rect 20216 18464 20232 18528
rect 20296 18464 20312 18528
rect 20376 18464 20392 18528
rect 20456 18464 20464 18528
rect 20144 17440 20464 18464
rect 20144 17376 20152 17440
rect 20216 17376 20232 17440
rect 20296 17376 20312 17440
rect 20376 17376 20392 17440
rect 20456 17376 20464 17440
rect 20144 16352 20464 17376
rect 20144 16288 20152 16352
rect 20216 16288 20232 16352
rect 20296 16288 20312 16352
rect 20376 16288 20392 16352
rect 20456 16288 20464 16352
rect 20144 15264 20464 16288
rect 20144 15200 20152 15264
rect 20216 15200 20232 15264
rect 20296 15200 20312 15264
rect 20376 15200 20392 15264
rect 20456 15200 20464 15264
rect 20144 14176 20464 15200
rect 20144 14112 20152 14176
rect 20216 14112 20232 14176
rect 20296 14112 20312 14176
rect 20376 14112 20392 14176
rect 20456 14112 20464 14176
rect 20144 13088 20464 14112
rect 20144 13024 20152 13088
rect 20216 13024 20232 13088
rect 20296 13024 20312 13088
rect 20376 13024 20392 13088
rect 20456 13024 20464 13088
rect 20144 12000 20464 13024
rect 20144 11936 20152 12000
rect 20216 11936 20232 12000
rect 20296 11936 20312 12000
rect 20376 11936 20392 12000
rect 20456 11936 20464 12000
rect 20144 10912 20464 11936
rect 20144 10848 20152 10912
rect 20216 10848 20232 10912
rect 20296 10848 20312 10912
rect 20376 10848 20392 10912
rect 20456 10848 20464 10912
rect 20144 9824 20464 10848
rect 20144 9760 20152 9824
rect 20216 9760 20232 9824
rect 20296 9760 20312 9824
rect 20376 9760 20392 9824
rect 20456 9760 20464 9824
rect 20144 8736 20464 9760
rect 20144 8672 20152 8736
rect 20216 8672 20232 8736
rect 20296 8672 20312 8736
rect 20376 8672 20392 8736
rect 20456 8672 20464 8736
rect 20144 7648 20464 8672
rect 20144 7584 20152 7648
rect 20216 7584 20232 7648
rect 20296 7584 20312 7648
rect 20376 7584 20392 7648
rect 20456 7584 20464 7648
rect 20144 6560 20464 7584
rect 20144 6496 20152 6560
rect 20216 6496 20232 6560
rect 20296 6496 20312 6560
rect 20376 6496 20392 6560
rect 20456 6496 20464 6560
rect 20144 5472 20464 6496
rect 20144 5408 20152 5472
rect 20216 5408 20232 5472
rect 20296 5408 20312 5472
rect 20376 5408 20392 5472
rect 20456 5408 20464 5472
rect 20144 4384 20464 5408
rect 20144 4320 20152 4384
rect 20216 4320 20232 4384
rect 20296 4320 20312 4384
rect 20376 4320 20392 4384
rect 20456 4320 20464 4384
rect 20144 3296 20464 4320
rect 20144 3232 20152 3296
rect 20216 3232 20232 3296
rect 20296 3232 20312 3296
rect 20376 3232 20392 3296
rect 20456 3232 20464 3296
rect 20144 2208 20464 3232
rect 20144 2144 20152 2208
rect 20216 2144 20232 2208
rect 20296 2144 20312 2208
rect 20376 2144 20392 2208
rect 20456 2144 20464 2208
rect 20144 2128 20464 2144
rect 22544 27776 22864 27792
rect 22544 27712 22552 27776
rect 22616 27712 22632 27776
rect 22696 27712 22712 27776
rect 22776 27712 22792 27776
rect 22856 27712 22864 27776
rect 22544 26688 22864 27712
rect 22544 26624 22552 26688
rect 22616 26624 22632 26688
rect 22696 26624 22712 26688
rect 22776 26624 22792 26688
rect 22856 26624 22864 26688
rect 22544 25600 22864 26624
rect 22544 25536 22552 25600
rect 22616 25536 22632 25600
rect 22696 25536 22712 25600
rect 22776 25536 22792 25600
rect 22856 25536 22864 25600
rect 22544 24512 22864 25536
rect 22544 24448 22552 24512
rect 22616 24448 22632 24512
rect 22696 24448 22712 24512
rect 22776 24448 22792 24512
rect 22856 24448 22864 24512
rect 22544 23424 22864 24448
rect 22544 23360 22552 23424
rect 22616 23360 22632 23424
rect 22696 23360 22712 23424
rect 22776 23360 22792 23424
rect 22856 23360 22864 23424
rect 22544 22336 22864 23360
rect 22544 22272 22552 22336
rect 22616 22272 22632 22336
rect 22696 22272 22712 22336
rect 22776 22272 22792 22336
rect 22856 22272 22864 22336
rect 22544 21248 22864 22272
rect 22544 21184 22552 21248
rect 22616 21184 22632 21248
rect 22696 21184 22712 21248
rect 22776 21184 22792 21248
rect 22856 21184 22864 21248
rect 22544 20160 22864 21184
rect 22544 20096 22552 20160
rect 22616 20096 22632 20160
rect 22696 20096 22712 20160
rect 22776 20096 22792 20160
rect 22856 20096 22864 20160
rect 22544 19072 22864 20096
rect 22544 19008 22552 19072
rect 22616 19008 22632 19072
rect 22696 19008 22712 19072
rect 22776 19008 22792 19072
rect 22856 19008 22864 19072
rect 22544 17984 22864 19008
rect 22544 17920 22552 17984
rect 22616 17920 22632 17984
rect 22696 17920 22712 17984
rect 22776 17920 22792 17984
rect 22856 17920 22864 17984
rect 22544 16896 22864 17920
rect 22544 16832 22552 16896
rect 22616 16832 22632 16896
rect 22696 16832 22712 16896
rect 22776 16832 22792 16896
rect 22856 16832 22864 16896
rect 22544 15808 22864 16832
rect 22544 15744 22552 15808
rect 22616 15744 22632 15808
rect 22696 15744 22712 15808
rect 22776 15744 22792 15808
rect 22856 15744 22864 15808
rect 22544 14720 22864 15744
rect 22544 14656 22552 14720
rect 22616 14656 22632 14720
rect 22696 14656 22712 14720
rect 22776 14656 22792 14720
rect 22856 14656 22864 14720
rect 22544 13632 22864 14656
rect 22544 13568 22552 13632
rect 22616 13568 22632 13632
rect 22696 13568 22712 13632
rect 22776 13568 22792 13632
rect 22856 13568 22864 13632
rect 22544 12544 22864 13568
rect 22544 12480 22552 12544
rect 22616 12480 22632 12544
rect 22696 12480 22712 12544
rect 22776 12480 22792 12544
rect 22856 12480 22864 12544
rect 22544 11456 22864 12480
rect 22544 11392 22552 11456
rect 22616 11392 22632 11456
rect 22696 11392 22712 11456
rect 22776 11392 22792 11456
rect 22856 11392 22864 11456
rect 22544 10368 22864 11392
rect 22544 10304 22552 10368
rect 22616 10304 22632 10368
rect 22696 10304 22712 10368
rect 22776 10304 22792 10368
rect 22856 10304 22864 10368
rect 22544 9280 22864 10304
rect 22544 9216 22552 9280
rect 22616 9216 22632 9280
rect 22696 9216 22712 9280
rect 22776 9216 22792 9280
rect 22856 9216 22864 9280
rect 22544 8192 22864 9216
rect 22544 8128 22552 8192
rect 22616 8128 22632 8192
rect 22696 8128 22712 8192
rect 22776 8128 22792 8192
rect 22856 8128 22864 8192
rect 22544 7104 22864 8128
rect 22544 7040 22552 7104
rect 22616 7040 22632 7104
rect 22696 7040 22712 7104
rect 22776 7040 22792 7104
rect 22856 7040 22864 7104
rect 22544 6016 22864 7040
rect 22544 5952 22552 6016
rect 22616 5952 22632 6016
rect 22696 5952 22712 6016
rect 22776 5952 22792 6016
rect 22856 5952 22864 6016
rect 22544 4928 22864 5952
rect 22544 4864 22552 4928
rect 22616 4864 22632 4928
rect 22696 4864 22712 4928
rect 22776 4864 22792 4928
rect 22856 4864 22864 4928
rect 22544 3840 22864 4864
rect 22544 3776 22552 3840
rect 22616 3776 22632 3840
rect 22696 3776 22712 3840
rect 22776 3776 22792 3840
rect 22856 3776 22864 3840
rect 22544 2752 22864 3776
rect 22544 2688 22552 2752
rect 22616 2688 22632 2752
rect 22696 2688 22712 2752
rect 22776 2688 22792 2752
rect 22856 2688 22864 2752
rect 22544 2128 22864 2688
rect 24944 27232 25264 27792
rect 24944 27168 24952 27232
rect 25016 27168 25032 27232
rect 25096 27168 25112 27232
rect 25176 27168 25192 27232
rect 25256 27168 25264 27232
rect 24944 26144 25264 27168
rect 24944 26080 24952 26144
rect 25016 26080 25032 26144
rect 25096 26080 25112 26144
rect 25176 26080 25192 26144
rect 25256 26080 25264 26144
rect 24944 25056 25264 26080
rect 24944 24992 24952 25056
rect 25016 24992 25032 25056
rect 25096 24992 25112 25056
rect 25176 24992 25192 25056
rect 25256 24992 25264 25056
rect 24944 23968 25264 24992
rect 24944 23904 24952 23968
rect 25016 23904 25032 23968
rect 25096 23904 25112 23968
rect 25176 23904 25192 23968
rect 25256 23904 25264 23968
rect 24944 22880 25264 23904
rect 24944 22816 24952 22880
rect 25016 22816 25032 22880
rect 25096 22816 25112 22880
rect 25176 22816 25192 22880
rect 25256 22816 25264 22880
rect 24944 21792 25264 22816
rect 24944 21728 24952 21792
rect 25016 21728 25032 21792
rect 25096 21728 25112 21792
rect 25176 21728 25192 21792
rect 25256 21728 25264 21792
rect 24944 20704 25264 21728
rect 24944 20640 24952 20704
rect 25016 20640 25032 20704
rect 25096 20640 25112 20704
rect 25176 20640 25192 20704
rect 25256 20640 25264 20704
rect 24944 19616 25264 20640
rect 24944 19552 24952 19616
rect 25016 19552 25032 19616
rect 25096 19552 25112 19616
rect 25176 19552 25192 19616
rect 25256 19552 25264 19616
rect 24944 18528 25264 19552
rect 24944 18464 24952 18528
rect 25016 18464 25032 18528
rect 25096 18464 25112 18528
rect 25176 18464 25192 18528
rect 25256 18464 25264 18528
rect 24944 17440 25264 18464
rect 24944 17376 24952 17440
rect 25016 17376 25032 17440
rect 25096 17376 25112 17440
rect 25176 17376 25192 17440
rect 25256 17376 25264 17440
rect 24944 16352 25264 17376
rect 24944 16288 24952 16352
rect 25016 16288 25032 16352
rect 25096 16288 25112 16352
rect 25176 16288 25192 16352
rect 25256 16288 25264 16352
rect 24944 15264 25264 16288
rect 24944 15200 24952 15264
rect 25016 15200 25032 15264
rect 25096 15200 25112 15264
rect 25176 15200 25192 15264
rect 25256 15200 25264 15264
rect 24944 14176 25264 15200
rect 24944 14112 24952 14176
rect 25016 14112 25032 14176
rect 25096 14112 25112 14176
rect 25176 14112 25192 14176
rect 25256 14112 25264 14176
rect 24944 13088 25264 14112
rect 24944 13024 24952 13088
rect 25016 13024 25032 13088
rect 25096 13024 25112 13088
rect 25176 13024 25192 13088
rect 25256 13024 25264 13088
rect 24944 12000 25264 13024
rect 24944 11936 24952 12000
rect 25016 11936 25032 12000
rect 25096 11936 25112 12000
rect 25176 11936 25192 12000
rect 25256 11936 25264 12000
rect 24944 10912 25264 11936
rect 24944 10848 24952 10912
rect 25016 10848 25032 10912
rect 25096 10848 25112 10912
rect 25176 10848 25192 10912
rect 25256 10848 25264 10912
rect 24944 9824 25264 10848
rect 24944 9760 24952 9824
rect 25016 9760 25032 9824
rect 25096 9760 25112 9824
rect 25176 9760 25192 9824
rect 25256 9760 25264 9824
rect 24944 8736 25264 9760
rect 24944 8672 24952 8736
rect 25016 8672 25032 8736
rect 25096 8672 25112 8736
rect 25176 8672 25192 8736
rect 25256 8672 25264 8736
rect 24944 7648 25264 8672
rect 24944 7584 24952 7648
rect 25016 7584 25032 7648
rect 25096 7584 25112 7648
rect 25176 7584 25192 7648
rect 25256 7584 25264 7648
rect 24944 6560 25264 7584
rect 24944 6496 24952 6560
rect 25016 6496 25032 6560
rect 25096 6496 25112 6560
rect 25176 6496 25192 6560
rect 25256 6496 25264 6560
rect 24944 5472 25264 6496
rect 24944 5408 24952 5472
rect 25016 5408 25032 5472
rect 25096 5408 25112 5472
rect 25176 5408 25192 5472
rect 25256 5408 25264 5472
rect 24944 4384 25264 5408
rect 24944 4320 24952 4384
rect 25016 4320 25032 4384
rect 25096 4320 25112 4384
rect 25176 4320 25192 4384
rect 25256 4320 25264 4384
rect 24944 3296 25264 4320
rect 24944 3232 24952 3296
rect 25016 3232 25032 3296
rect 25096 3232 25112 3296
rect 25176 3232 25192 3296
rect 25256 3232 25264 3296
rect 24944 2208 25264 3232
rect 24944 2144 24952 2208
rect 25016 2144 25032 2208
rect 25096 2144 25112 2208
rect 25176 2144 25192 2208
rect 25256 2144 25264 2208
rect 24944 2128 25264 2144
rect 27344 27776 27664 27792
rect 27344 27712 27352 27776
rect 27416 27712 27432 27776
rect 27496 27712 27512 27776
rect 27576 27712 27592 27776
rect 27656 27712 27664 27776
rect 27344 26688 27664 27712
rect 27344 26624 27352 26688
rect 27416 26624 27432 26688
rect 27496 26624 27512 26688
rect 27576 26624 27592 26688
rect 27656 26624 27664 26688
rect 27344 25600 27664 26624
rect 27344 25536 27352 25600
rect 27416 25536 27432 25600
rect 27496 25536 27512 25600
rect 27576 25536 27592 25600
rect 27656 25536 27664 25600
rect 27344 24512 27664 25536
rect 27344 24448 27352 24512
rect 27416 24448 27432 24512
rect 27496 24448 27512 24512
rect 27576 24448 27592 24512
rect 27656 24448 27664 24512
rect 27344 23424 27664 24448
rect 27344 23360 27352 23424
rect 27416 23360 27432 23424
rect 27496 23360 27512 23424
rect 27576 23360 27592 23424
rect 27656 23360 27664 23424
rect 27344 22336 27664 23360
rect 27344 22272 27352 22336
rect 27416 22272 27432 22336
rect 27496 22272 27512 22336
rect 27576 22272 27592 22336
rect 27656 22272 27664 22336
rect 27344 21248 27664 22272
rect 27344 21184 27352 21248
rect 27416 21184 27432 21248
rect 27496 21184 27512 21248
rect 27576 21184 27592 21248
rect 27656 21184 27664 21248
rect 27344 20160 27664 21184
rect 27344 20096 27352 20160
rect 27416 20096 27432 20160
rect 27496 20096 27512 20160
rect 27576 20096 27592 20160
rect 27656 20096 27664 20160
rect 27344 19072 27664 20096
rect 27344 19008 27352 19072
rect 27416 19008 27432 19072
rect 27496 19008 27512 19072
rect 27576 19008 27592 19072
rect 27656 19008 27664 19072
rect 27344 17984 27664 19008
rect 27344 17920 27352 17984
rect 27416 17920 27432 17984
rect 27496 17920 27512 17984
rect 27576 17920 27592 17984
rect 27656 17920 27664 17984
rect 27344 16896 27664 17920
rect 27344 16832 27352 16896
rect 27416 16832 27432 16896
rect 27496 16832 27512 16896
rect 27576 16832 27592 16896
rect 27656 16832 27664 16896
rect 27344 15808 27664 16832
rect 27344 15744 27352 15808
rect 27416 15744 27432 15808
rect 27496 15744 27512 15808
rect 27576 15744 27592 15808
rect 27656 15744 27664 15808
rect 27344 14720 27664 15744
rect 27344 14656 27352 14720
rect 27416 14656 27432 14720
rect 27496 14656 27512 14720
rect 27576 14656 27592 14720
rect 27656 14656 27664 14720
rect 27344 13632 27664 14656
rect 27344 13568 27352 13632
rect 27416 13568 27432 13632
rect 27496 13568 27512 13632
rect 27576 13568 27592 13632
rect 27656 13568 27664 13632
rect 27344 12544 27664 13568
rect 27344 12480 27352 12544
rect 27416 12480 27432 12544
rect 27496 12480 27512 12544
rect 27576 12480 27592 12544
rect 27656 12480 27664 12544
rect 27344 11456 27664 12480
rect 27344 11392 27352 11456
rect 27416 11392 27432 11456
rect 27496 11392 27512 11456
rect 27576 11392 27592 11456
rect 27656 11392 27664 11456
rect 27344 10368 27664 11392
rect 27344 10304 27352 10368
rect 27416 10304 27432 10368
rect 27496 10304 27512 10368
rect 27576 10304 27592 10368
rect 27656 10304 27664 10368
rect 27344 9280 27664 10304
rect 27344 9216 27352 9280
rect 27416 9216 27432 9280
rect 27496 9216 27512 9280
rect 27576 9216 27592 9280
rect 27656 9216 27664 9280
rect 27344 8192 27664 9216
rect 27344 8128 27352 8192
rect 27416 8128 27432 8192
rect 27496 8128 27512 8192
rect 27576 8128 27592 8192
rect 27656 8128 27664 8192
rect 27344 7104 27664 8128
rect 27344 7040 27352 7104
rect 27416 7040 27432 7104
rect 27496 7040 27512 7104
rect 27576 7040 27592 7104
rect 27656 7040 27664 7104
rect 27344 6016 27664 7040
rect 27344 5952 27352 6016
rect 27416 5952 27432 6016
rect 27496 5952 27512 6016
rect 27576 5952 27592 6016
rect 27656 5952 27664 6016
rect 27344 4928 27664 5952
rect 27344 4864 27352 4928
rect 27416 4864 27432 4928
rect 27496 4864 27512 4928
rect 27576 4864 27592 4928
rect 27656 4864 27664 4928
rect 27344 3840 27664 4864
rect 27344 3776 27352 3840
rect 27416 3776 27432 3840
rect 27496 3776 27512 3840
rect 27576 3776 27592 3840
rect 27656 3776 27664 3840
rect 27344 2752 27664 3776
rect 27344 2688 27352 2752
rect 27416 2688 27432 2752
rect 27496 2688 27512 2752
rect 27576 2688 27592 2752
rect 27656 2688 27664 2752
rect 27344 2128 27664 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__150__S pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 22908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__S
timestamp 1670032574
transform -1 0 21896 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__S
timestamp 1670032574
transform 1 0 24564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__S
timestamp 1670032574
transform 1 0 24104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__S
timestamp 1670032574
transform 1 0 22816 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__S
timestamp 1670032574
transform 1 0 24012 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__S
timestamp 1670032574
transform 1 0 24380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__S
timestamp 1670032574
transform 1 0 24012 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__S
timestamp 1670032574
transform 1 0 24288 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__S
timestamp 1670032574
transform -1 0 23092 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__B
timestamp 1670032574
transform 1 0 18860 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1670032574
transform 1 0 17940 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1670032574
transform 1 0 8464 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1670032574
transform -1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1670032574
transform 1 0 7084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1670032574
transform 1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A
timestamp 1670032574
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1670032574
transform 1 0 12236 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1670032574
transform -1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1670032574
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A
timestamp 1670032574
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1670032574
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1670032574
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__S
timestamp 1670032574
transform 1 0 25024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__S
timestamp 1670032574
transform 1 0 26588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__S
timestamp 1670032574
transform 1 0 27508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__S
timestamp 1670032574
transform 1 0 26588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__S
timestamp 1670032574
transform 1 0 26588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__S
timestamp 1670032574
transform 1 0 26588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__S
timestamp 1670032574
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__S
timestamp 1670032574
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__S
timestamp 1670032574
transform 1 0 3864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__S
timestamp 1670032574
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__S
timestamp 1670032574
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__S
timestamp 1670032574
transform 1 0 3772 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A2
timestamp 1670032574
transform 1 0 18308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__B1
timestamp 1670032574
transform 1 0 18124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A
timestamp 1670032574
transform 1 0 9752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__B1
timestamp 1670032574
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__B1
timestamp 1670032574
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__B1
timestamp 1670032574
transform 1 0 5244 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__B1
timestamp 1670032574
transform 1 0 5980 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__C1
timestamp 1670032574
transform -1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A2
timestamp 1670032574
transform 1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__RESET_B
timestamp 1670032574
transform -1 0 26128 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__RESET_B
timestamp 1670032574
transform 1 0 3864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__RESET_B
timestamp 1670032574
transform 1 0 3864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__RESET_B
timestamp 1670032574
transform 1 0 3312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__RESET_B
timestamp 1670032574
transform 1 0 23092 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__RESET_B
timestamp 1670032574
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__RESET_B
timestamp 1670032574
transform 1 0 4508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__RESET_B
timestamp 1670032574
transform 1 0 11592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__RESET_B
timestamp 1670032574
transform 1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__SET_B
timestamp 1670032574
transform 1 0 12696 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1670032574
transform 1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_clk_A
timestamp 1670032574
transform 1 0 9844 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_clk_A
timestamp 1670032574
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_clk_A
timestamp 1670032574
transform -1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_clk_A
timestamp 1670032574
transform -1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_clk_A
timestamp 1670032574
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_clk_A
timestamp 1670032574
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_clk_A
timestamp 1670032574
transform 1 0 20608 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_clk_A
timestamp 1670032574
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref_A
timestamp 1670032574
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref_A
timestamp 1670032574
transform 1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref_A
timestamp 1670032574
transform 1 0 8188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref_A
timestamp 1670032574
transform 1 0 12420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref_A
timestamp 1670032574
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref_A
timestamp 1670032574
transform 1 0 12604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref_A
timestamp 1670032574
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref_A
timestamp 1670032574
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref_A
timestamp 1670032574
transform 1 0 13800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref_A
timestamp 1670032574
transform 1 0 12972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref_A
timestamp 1670032574
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref_A
timestamp 1670032574
transform 1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref_A
timestamp 1670032574
transform 1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref_A
timestamp 1670032574
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref_A
timestamp 1670032574
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref_A
timestamp 1670032574
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref_A
timestamp 1670032574
transform 1 0 11592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref_A
timestamp 1670032574
transform 1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref_A
timestamp 1670032574
transform 1 0 10304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref_A
timestamp 1670032574
transform 1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref_A
timestamp 1670032574
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref_A
timestamp 1670032574
transform 1 0 11960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref_A
timestamp 1670032574
transform 1 0 12604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref_A
timestamp 1670032574
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref_A
timestamp 1670032574
transform 1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref_A
timestamp 1670032574
transform 1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref_A
timestamp 1670032574
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref_A
timestamp 1670032574
transform 1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref_A
timestamp 1670032574
transform 1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref_A
timestamp 1670032574
transform 1 0 11592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref_A
timestamp 1670032574
transform 1 0 11132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dac.vdac_single.einvp_batch\[0\].vref_A
timestamp 1670032574
transform 1 0 5152 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_dcdc_TE
timestamp 1670032574
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout22_A
timestamp 1670032574
transform 1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout23_A
timestamp 1670032574
transform -1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout25_A
timestamp 1670032574
transform -1 0 19872 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout27_A
timestamp 1670032574
transform 1 0 17020 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1670032574
transform -1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1670032574
transform -1 0 19504 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1670032574
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1670032574
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1670032574
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1670032574
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1670032574
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1670032574
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1670032574
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1670032574
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1670032574
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1670032574
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121
timestamp 1670032574
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1670032574
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1670032574
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1670032574
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1670032574
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1670032574
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_181 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_189
timestamp 1670032574
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1670032574
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 1670032574
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_200
timestamp 1670032574
transform 1 0 19504 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_212
timestamp 1670032574
transform 1 0 20608 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1670032574
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1670032574
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1670032574
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1670032574
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_265
timestamp 1670032574
transform 1 0 25484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1670032574
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1670032574
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1670032574
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 1670032574
transform 1 0 28520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1670032574
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1670032574
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1670032574
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_29
timestamp 1670032574
transform 1 0 3772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_41
timestamp 1670032574
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1670032574
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1670032574
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1670032574
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1670032574
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1670032574
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1670032574
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1670032574
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1670032574
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1670032574
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1670032574
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1670032574
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1670032574
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1670032574
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1670032574
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_181
timestamp 1670032574
transform 1 0 17756 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_189
timestamp 1670032574
transform 1 0 18492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_201
timestamp 1670032574
transform 1 0 19596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_204
timestamp 1670032574
transform 1 0 19872 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1670032574
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1670032574
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_229
timestamp 1670032574
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_250
timestamp 1670032574
transform 1 0 24104 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1670032574
transform 1 0 24840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_262
timestamp 1670032574
transform 1 0 25208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1670032574
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1670032574
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1670032574
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1670032574
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1670032574
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1670032574
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1670032574
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_32
timestamp 1670032574
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_44
timestamp 1670032574
transform 1 0 5152 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_56
timestamp 1670032574
transform 1 0 6256 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_68
timestamp 1670032574
transform 1 0 7360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1670032574
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1670032574
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1670032574
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1670032574
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1670032574
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1670032574
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1670032574
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1670032574
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1670032574
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1670032574
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp 1670032574
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1670032574
transform 1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1670032574
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp 1670032574
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1670032574
transform 1 0 21160 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_240
timestamp 1670032574
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1670032574
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_257
timestamp 1670032574
transform 1 0 24748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_278
timestamp 1670032574
transform 1 0 26680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_285
timestamp 1670032574
transform 1 0 27324 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_293
timestamp 1670032574
transform 1 0 28060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1670032574
transform 1 0 28520 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1670032574
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1670032574
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1670032574
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1670032574
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1670032574
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1670032574
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1670032574
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1670032574
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1670032574
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1670032574
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1670032574
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1670032574
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1670032574
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1670032574
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1670032574
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1670032574
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1670032574
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1670032574
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1670032574
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1670032574
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_212
timestamp 1670032574
transform 1 0 20608 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1670032574
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_230
timestamp 1670032574
transform 1 0 22264 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_238
timestamp 1670032574
transform 1 0 23000 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_243
timestamp 1670032574
transform 1 0 23460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_255
timestamp 1670032574
transform 1 0 24564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_261
timestamp 1670032574
transform 1 0 25116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_265
timestamp 1670032574
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1670032574
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp 1670032574
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1670032574
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1670032574
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_15
timestamp 1670032574
transform 1 0 2484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_23
timestamp 1670032574
transform 1 0 3220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1670032574
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1670032574
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1670032574
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1670032574
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1670032574
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1670032574
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1670032574
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1670032574
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1670032574
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_101
timestamp 1670032574
transform 1 0 10396 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1670032574
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_108
timestamp 1670032574
transform 1 0 11040 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_111
timestamp 1670032574
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_123
timestamp 1670032574
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1670032574
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1670032574
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1670032574
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1670032574
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1670032574
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1670032574
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1670032574
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1670032574
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1670032574
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1670032574
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp 1670032574
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_226
timestamp 1670032574
transform 1 0 21896 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_237
timestamp 1670032574
transform 1 0 22908 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1670032574
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1670032574
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1670032574
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_277
timestamp 1670032574
transform 1 0 26588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1670032574
transform 1 0 28520 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1670032574
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1670032574
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1670032574
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1670032574
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1670032574
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1670032574
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1670032574
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1670032574
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1670032574
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1670032574
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_97
timestamp 1670032574
transform 1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1670032574
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1670032574
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1670032574
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_116
timestamp 1670032574
transform 1 0 11776 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_120
timestamp 1670032574
transform 1 0 12144 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_132
timestamp 1670032574
transform 1 0 13248 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_144
timestamp 1670032574
transform 1 0 14352 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_156
timestamp 1670032574
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1670032574
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1670032574
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_189
timestamp 1670032574
transform 1 0 18492 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1670032574
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1670032574
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1670032574
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_239
timestamp 1670032574
transform 1 0 23092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_251
timestamp 1670032574
transform 1 0 24196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_263
timestamp 1670032574
transform 1 0 25300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1670032574
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1670032574
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1670032574
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1670032574
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1670032574
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1670032574
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1670032574
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1670032574
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1670032574
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_53
timestamp 1670032574
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp 1670032574
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1670032574
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_72
timestamp 1670032574
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1670032574
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_90
timestamp 1670032574
transform 1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_95
timestamp 1670032574
transform 1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1670032574
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1670032574
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_116
timestamp 1670032574
transform 1 0 11776 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_123
timestamp 1670032574
transform 1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_127
timestamp 1670032574
transform 1 0 12788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1670032574
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1670032574
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1670032574
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1670032574
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1670032574
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1670032574
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1670032574
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 1670032574
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_202
timestamp 1670032574
transform 1 0 19688 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_214
timestamp 1670032574
transform 1 0 20792 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_226
timestamp 1670032574
transform 1 0 21896 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_238
timestamp 1670032574
transform 1 0 23000 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1670032574
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1670032574
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_257
timestamp 1670032574
transform 1 0 24748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_268
timestamp 1670032574
transform 1 0 25760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1670032574
transform 1 0 26496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1670032574
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1670032574
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1670032574
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1670032574
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 1670032574
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_37
timestamp 1670032574
transform 1 0 4508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_42
timestamp 1670032574
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_46
timestamp 1670032574
transform 1 0 5336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1670032574
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 1670032574
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1670032574
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_72
timestamp 1670032574
transform 1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_79
timestamp 1670032574
transform 1 0 8372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_85
timestamp 1670032574
transform 1 0 8924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1670032574
transform 1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_95
timestamp 1670032574
transform 1 0 9844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1670032574
transform 1 0 10488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1670032574
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1670032574
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_119
timestamp 1670032574
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_126
timestamp 1670032574
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp 1670032574
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1670032574
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1670032574
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1670032574
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1670032574
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1670032574
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1670032574
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_193
timestamp 1670032574
transform 1 0 18860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1670032574
transform 1 0 19412 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1670032574
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_216
timestamp 1670032574
transform 1 0 20976 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1670032574
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1670032574
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_232
timestamp 1670032574
transform 1 0 22448 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_244
timestamp 1670032574
transform 1 0 23552 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_256
timestamp 1670032574
transform 1 0 24656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1670032574
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp 1670032574
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1670032574
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1670032574
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1670032574
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1670032574
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1670032574
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1670032574
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1670032574
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_51
timestamp 1670032574
transform 1 0 5796 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_58
timestamp 1670032574
transform 1 0 6440 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1670032574
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_72
timestamp 1670032574
transform 1 0 7728 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1670032574
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1670032574
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1670032574
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_95
timestamp 1670032574
transform 1 0 9844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1670032574
transform 1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1670032574
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1670032574
transform 1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 1670032574
transform 1 0 12420 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_127
timestamp 1670032574
transform 1 0 12788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1670032574
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1670032574
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1670032574
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1670032574
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_177
timestamp 1670032574
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_185
timestamp 1670032574
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_191
timestamp 1670032574
transform 1 0 18676 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1670032574
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1670032574
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1670032574
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1670032574
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_219
timestamp 1670032574
transform 1 0 21252 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1670032574
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1670032574
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp 1670032574
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_261
timestamp 1670032574
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1670032574
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_277
timestamp 1670032574
transform 1 0 26588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_281
timestamp 1670032574
transform 1 0 26956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_285
timestamp 1670032574
transform 1 0 27324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_289
timestamp 1670032574
transform 1 0 27692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_293
timestamp 1670032574
transform 1 0 28060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1670032574
transform 1 0 28520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1670032574
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_8
timestamp 1670032574
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1670032574
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1670032574
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_44
timestamp 1670032574
transform 1 0 5152 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1670032574
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1670032574
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1670032574
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_72
timestamp 1670032574
transform 1 0 7728 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_84
timestamp 1670032574
transform 1 0 8832 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_92
timestamp 1670032574
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_97
timestamp 1670032574
transform 1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1670032574
transform 1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1670032574
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1670032574
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_116
timestamp 1670032574
transform 1 0 11776 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_128
timestamp 1670032574
transform 1 0 12880 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1670032574
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_140
timestamp 1670032574
transform 1 0 13984 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_152
timestamp 1670032574
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1670032574
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1670032574
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_177
timestamp 1670032574
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_201
timestamp 1670032574
transform 1 0 19596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_213
timestamp 1670032574
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1670032574
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_225
timestamp 1670032574
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_233
timestamp 1670032574
transform 1 0 22540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_245
timestamp 1670032574
transform 1 0 23644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_257
timestamp 1670032574
transform 1 0 24748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1670032574
transform 1 0 25852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1670032574
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1670032574
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1670032574
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1670032574
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1670032574
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1670032574
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_32
timestamp 1670032574
transform 1 0 4048 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_44
timestamp 1670032574
transform 1 0 5152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1670032574
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1670032574
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_72
timestamp 1670032574
transform 1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1670032574
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1670032574
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1670032574
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_96
timestamp 1670032574
transform 1 0 9936 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_108
timestamp 1670032574
transform 1 0 11040 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1670032574
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_126
timestamp 1670032574
transform 1 0 12696 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1670032574
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1670032574
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1670032574
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_147
timestamp 1670032574
transform 1 0 14628 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_151
timestamp 1670032574
transform 1 0 14996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_163
timestamp 1670032574
transform 1 0 16100 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_175
timestamp 1670032574
transform 1 0 17204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1670032574
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1670032574
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1670032574
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp 1670032574
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1670032574
transform 1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_234
timestamp 1670032574
transform 1 0 22632 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1670032574
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1670032574
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1670032574
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1670032574
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1670032574
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_289
timestamp 1670032574
transform 1 0 27692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1670032574
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1670032574
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_14
timestamp 1670032574
transform 1 0 2392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_25
timestamp 1670032574
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_29
timestamp 1670032574
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_41
timestamp 1670032574
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1670032574
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1670032574
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_63
timestamp 1670032574
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1670032574
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1670032574
transform 1 0 8464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_87
timestamp 1670032574
transform 1 0 9108 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_91
timestamp 1670032574
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1670032574
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1670032574
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1670032574
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1670032574
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_124
timestamp 1670032574
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_131
timestamp 1670032574
transform 1 0 13156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_138
timestamp 1670032574
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_145
timestamp 1670032574
transform 1 0 14444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1670032574
transform 1 0 15088 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_156
timestamp 1670032574
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1670032574
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_181
timestamp 1670032574
transform 1 0 17756 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1670032574
transform 1 0 18032 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_206
timestamp 1670032574
transform 1 0 20056 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1670032574
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_225
timestamp 1670032574
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_230
timestamp 1670032574
transform 1 0 22264 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_235
timestamp 1670032574
transform 1 0 22724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_247
timestamp 1670032574
transform 1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_252
timestamp 1670032574
transform 1 0 24288 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_263
timestamp 1670032574
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_275
timestamp 1670032574
transform 1 0 26404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1670032574
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp 1670032574
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1670032574
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1670032574
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1670032574
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1670032574
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1670032574
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_33
timestamp 1670032574
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_39
timestamp 1670032574
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_51
timestamp 1670032574
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_63
timestamp 1670032574
transform 1 0 6900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1670032574
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1670032574
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1670032574
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1670032574
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_93
timestamp 1670032574
transform 1 0 9660 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_105
timestamp 1670032574
transform 1 0 10764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_113
timestamp 1670032574
transform 1 0 11500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_119
timestamp 1670032574
transform 1 0 12052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1670032574
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1670032574
transform 1 0 12788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_131
timestamp 1670032574
transform 1 0 13156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1670032574
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1670032574
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_147
timestamp 1670032574
transform 1 0 14628 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_151
timestamp 1670032574
transform 1 0 14996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_163
timestamp 1670032574
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_175
timestamp 1670032574
transform 1 0 17204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1670032574
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1670032574
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1670032574
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1670032574
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1670032574
transform 1 0 21436 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_242
timestamp 1670032574
transform 1 0 23368 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1670032574
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_253
timestamp 1670032574
transform 1 0 24380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_274
timestamp 1670032574
transform 1 0 26312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_296
timestamp 1670032574
transform 1 0 28336 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1670032574
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1670032574
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_27
timestamp 1670032574
transform 1 0 3588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_33
timestamp 1670032574
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_39
timestamp 1670032574
transform 1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1670032574
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1670032574
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1670032574
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_69
timestamp 1670032574
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_77
timestamp 1670032574
transform 1 0 8188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1670032574
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1670032574
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1670032574
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_99
timestamp 1670032574
transform 1 0 10212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_107
timestamp 1670032574
transform 1 0 10948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1670032574
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1670032574
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_119
timestamp 1670032574
transform 1 0 12052 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1670032574
transform 1 0 12420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1670032574
transform 1 0 13248 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_136
timestamp 1670032574
transform 1 0 13616 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_148
timestamp 1670032574
transform 1 0 14720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1670032574
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1670032574
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 1670032574
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_184
timestamp 1670032574
transform 1 0 18032 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_196
timestamp 1670032574
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1670032574
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1670032574
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1670032574
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1670032574
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_249
timestamp 1670032574
transform 1 0 24012 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_255
timestamp 1670032574
transform 1 0 24564 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_259
timestamp 1670032574
transform 1 0 24932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1670032574
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1670032574
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_281
timestamp 1670032574
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_285
timestamp 1670032574
transform 1 0 27324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_293
timestamp 1670032574
transform 1 0 28060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1670032574
transform 1 0 28520 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1670032574
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1670032574
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1670032574
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1670032574
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1670032574
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_39
timestamp 1670032574
transform 1 0 4692 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_46
timestamp 1670032574
transform 1 0 5336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_56
timestamp 1670032574
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1670032574
transform 1 0 6900 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_67
timestamp 1670032574
transform 1 0 7268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1670032574
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1670032574
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1670032574
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_92
timestamp 1670032574
transform 1 0 9568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_99
timestamp 1670032574
transform 1 0 10212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1670032574
transform 1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1670032574
transform 1 0 12604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1670032574
transform 1 0 13248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1670032574
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1670032574
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_153
timestamp 1670032574
transform 1 0 15180 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_182
timestamp 1670032574
transform 1 0 17848 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1670032574
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1670032574
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_205
timestamp 1670032574
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_226
timestamp 1670032574
transform 1 0 21896 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_238
timestamp 1670032574
transform 1 0 23000 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1670032574
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1670032574
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1670032574
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1670032574
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1670032574
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1670032574
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1670032574
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1670032574
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_27
timestamp 1670032574
transform 1 0 3588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_33
timestamp 1670032574
transform 1 0 4140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_39
timestamp 1670032574
transform 1 0 4692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 1670032574
transform 1 0 5336 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1670032574
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1670032574
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1670032574
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1670032574
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_97
timestamp 1670032574
transform 1 0 10028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1670032574
transform 1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1670032574
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1670032574
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_120
timestamp 1670032574
transform 1 0 12144 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_126
timestamp 1670032574
transform 1 0 12696 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1670032574
transform 1 0 13248 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_136
timestamp 1670032574
transform 1 0 13616 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_148
timestamp 1670032574
transform 1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1670032574
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1670032574
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1670032574
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 1670032574
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_201
timestamp 1670032574
transform 1 0 19596 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_209
timestamp 1670032574
transform 1 0 20332 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_214
timestamp 1670032574
transform 1 0 20792 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1670032574
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1670032574
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_233
timestamp 1670032574
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_238
timestamp 1670032574
transform 1 0 23000 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1670032574
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1670032574
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_273
timestamp 1670032574
transform 1 0 26220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1670032574
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_281
timestamp 1670032574
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1670032574
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1670032574
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1670032574
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1670032574
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1670032574
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1670032574
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_39
timestamp 1670032574
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1670032574
transform 1 0 5796 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_61
timestamp 1670032574
transform 1 0 6716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1670032574
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_75
timestamp 1670032574
transform 1 0 8004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1670032574
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1670032574
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1670032574
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_96
timestamp 1670032574
transform 1 0 9936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_101
timestamp 1670032574
transform 1 0 10396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1670032574
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_113
timestamp 1670032574
transform 1 0 11500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1670032574
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1670032574
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1670032574
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1670032574
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_153
timestamp 1670032574
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1670032574
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_185
timestamp 1670032574
transform 1 0 18124 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1670032574
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1670032574
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1670032574
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_221
timestamp 1670032574
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_229
timestamp 1670032574
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1670032574
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1670032574
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_265
timestamp 1670032574
transform 1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_273
timestamp 1670032574
transform 1 0 26220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_296
timestamp 1670032574
transform 1 0 28336 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1670032574
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_35
timestamp 1670032574
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1670032574
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1670032574
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1670032574
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp 1670032574
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1670032574
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1670032574
transform 1 0 7544 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_74
timestamp 1670032574
transform 1 0 7912 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_86
timestamp 1670032574
transform 1 0 9016 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_98
timestamp 1670032574
transform 1 0 10120 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1670032574
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1670032574
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_125
timestamp 1670032574
transform 1 0 12604 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1670032574
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1670032574
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_140
timestamp 1670032574
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_152
timestamp 1670032574
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1670032574
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1670032574
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_185
timestamp 1670032574
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_189
timestamp 1670032574
transform 1 0 18492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_201
timestamp 1670032574
transform 1 0 19596 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1670032574
transform 1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1670032574
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1670032574
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1670032574
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_237
timestamp 1670032574
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_246
timestamp 1670032574
transform 1 0 23736 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_258
timestamp 1670032574
transform 1 0 24840 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_270
timestamp 1670032574
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1670032574
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_281
timestamp 1670032574
transform 1 0 26956 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_285
timestamp 1670032574
transform 1 0 27324 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_293
timestamp 1670032574
transform 1 0 28060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp 1670032574
transform 1 0 28520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1670032574
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_8
timestamp 1670032574
transform 1 0 1840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_21
timestamp 1670032574
transform 1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1670032574
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1670032574
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_32
timestamp 1670032574
transform 1 0 4048 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_44
timestamp 1670032574
transform 1 0 5152 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_50
timestamp 1670032574
transform 1 0 5704 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1670032574
transform 1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_58
timestamp 1670032574
transform 1 0 6440 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_65
timestamp 1670032574
transform 1 0 7084 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_72
timestamp 1670032574
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1670032574
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1670032574
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_96
timestamp 1670032574
transform 1 0 9936 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1670032574
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_112
timestamp 1670032574
transform 1 0 11408 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_120
timestamp 1670032574
transform 1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1670032574
transform 1 0 12788 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1670032574
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1670032574
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1670032574
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_153
timestamp 1670032574
transform 1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_163
timestamp 1670032574
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_175
timestamp 1670032574
transform 1 0 17204 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_182
timestamp 1670032574
transform 1 0 17848 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1670032574
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1670032574
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_225
timestamp 1670032574
transform 1 0 21804 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_237
timestamp 1670032574
transform 1 0 22908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1670032574
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_253
timestamp 1670032574
transform 1 0 24380 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1670032574
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1670032574
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1670032574
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1670032574
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1670032574
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_24
timestamp 1670032574
transform 1 0 3312 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_28
timestamp 1670032574
transform 1 0 3680 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1670032574
transform 1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_41
timestamp 1670032574
transform 1 0 4876 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_47
timestamp 1670032574
transform 1 0 5428 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1670032574
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1670032574
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1670032574
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_70
timestamp 1670032574
transform 1 0 7544 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_83
timestamp 1670032574
transform 1 0 8740 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1670032574
transform 1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_100
timestamp 1670032574
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1670032574
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1670032574
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_124
timestamp 1670032574
transform 1 0 12512 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_136
timestamp 1670032574
transform 1 0 13616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1670032574
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1670032574
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1670032574
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_177
timestamp 1670032574
transform 1 0 17388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_189
timestamp 1670032574
transform 1 0 18492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_201
timestamp 1670032574
transform 1 0 19596 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_214
timestamp 1670032574
transform 1 0 20792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1670032574
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_225
timestamp 1670032574
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_231
timestamp 1670032574
transform 1 0 22356 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_243
timestamp 1670032574
transform 1 0 23460 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_251
timestamp 1670032574
transform 1 0 24196 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_273
timestamp 1670032574
transform 1 0 26220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1670032574
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1670032574
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1670032574
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1670032574
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1670032574
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1670032574
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1670032574
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1670032574
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_37
timestamp 1670032574
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_44
timestamp 1670032574
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_56
timestamp 1670032574
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_68
timestamp 1670032574
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_80
timestamp 1670032574
transform 1 0 8464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1670032574
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1670032574
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_106
timestamp 1670032574
transform 1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_114
timestamp 1670032574
transform 1 0 11592 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_126
timestamp 1670032574
transform 1 0 12696 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1670032574
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1670032574
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1670032574
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1670032574
transform 1 0 14444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_152
timestamp 1670032574
transform 1 0 15088 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_157
timestamp 1670032574
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1670032574
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_168
timestamp 1670032574
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_179
timestamp 1670032574
transform 1 0 17572 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1670032574
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1670032574
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1670032574
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_209
timestamp 1670032574
transform 1 0 20332 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1670032574
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_234
timestamp 1670032574
transform 1 0 22632 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1670032574
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_253
timestamp 1670032574
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_262
timestamp 1670032574
transform 1 0 25208 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_274
timestamp 1670032574
transform 1 0 26312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1670032574
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1670032574
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1670032574
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1670032574
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1670032574
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1670032574
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1670032574
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1670032574
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_64
timestamp 1670032574
transform 1 0 6992 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_76
timestamp 1670032574
transform 1 0 8096 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_88
timestamp 1670032574
transform 1 0 9200 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_100
timestamp 1670032574
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1670032574
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_128
timestamp 1670032574
transform 1 0 12880 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_137
timestamp 1670032574
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_143
timestamp 1670032574
transform 1 0 14260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1670032574
transform 1 0 14996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1670032574
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1670032574
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1670032574
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1670032574
transform 1 0 17204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_179
timestamp 1670032574
transform 1 0 17572 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_208
timestamp 1670032574
transform 1 0 20240 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_216
timestamp 1670032574
transform 1 0 20976 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1670032574
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_225
timestamp 1670032574
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_230
timestamp 1670032574
transform 1 0 22264 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_252
timestamp 1670032574
transform 1 0 24288 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_260
timestamp 1670032574
transform 1 0 25024 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_272
timestamp 1670032574
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_281
timestamp 1670032574
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_285
timestamp 1670032574
transform 1 0 27324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_293
timestamp 1670032574
transform 1 0 28060 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_298
timestamp 1670032574
transform 1 0 28520 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1670032574
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1670032574
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1670032574
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1670032574
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_38
timestamp 1670032574
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_42
timestamp 1670032574
transform 1 0 4968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_49
timestamp 1670032574
transform 1 0 5612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1670032574
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_63
timestamp 1670032574
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1670032574
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1670032574
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1670032574
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1670032574
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1670032574
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1670032574
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1670032574
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1670032574
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1670032574
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1670032574
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_173
timestamp 1670032574
transform 1 0 17020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 1670032574
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1670032574
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1670032574
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1670032574
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_221
timestamp 1670032574
transform 1 0 21436 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_229
timestamp 1670032574
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_241
timestamp 1670032574
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1670032574
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1670032574
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1670032574
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1670032574
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1670032574
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1670032574
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1670032574
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_15
timestamp 1670032574
transform 1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_21
timestamp 1670032574
transform 1 0 3036 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_42
timestamp 1670032574
transform 1 0 4968 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_48
timestamp 1670032574
transform 1 0 5520 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1670032574
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1670032574
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1670032574
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_67
timestamp 1670032574
transform 1 0 7268 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_90
timestamp 1670032574
transform 1 0 9384 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1670032574
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1670032574
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1670032574
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 1670032574
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_128
timestamp 1670032574
transform 1 0 12880 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_140
timestamp 1670032574
transform 1 0 13984 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_152
timestamp 1670032574
transform 1 0 15088 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1670032574
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1670032574
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_175
timestamp 1670032574
transform 1 0 17204 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_187
timestamp 1670032574
transform 1 0 18308 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_194
timestamp 1670032574
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_200
timestamp 1670032574
transform 1 0 19504 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 1670032574
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1670032574
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_225
timestamp 1670032574
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_232
timestamp 1670032574
transform 1 0 22448 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_244
timestamp 1670032574
transform 1 0 23552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_252
timestamp 1670032574
transform 1 0 24288 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_255
timestamp 1670032574
transform 1 0 24564 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_266
timestamp 1670032574
transform 1 0 25576 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1670032574
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1670032574
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1670032574
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1670032574
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1670032574
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1670032574
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1670032574
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1670032574
transform 1 0 7084 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_69
timestamp 1670032574
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1670032574
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1670032574
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_92
timestamp 1670032574
transform 1 0 9568 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1670032574
transform 1 0 10304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1670032574
transform 1 0 12236 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_125
timestamp 1670032574
transform 1 0 12604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1670032574
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1670032574
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1670032574
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1670032574
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1670032574
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1670032574
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1670032574
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1670032574
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1670032574
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1670032574
transform 1 0 20608 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_234
timestamp 1670032574
transform 1 0 22632 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1670032574
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_253
timestamp 1670032574
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_274
timestamp 1670032574
transform 1 0 26312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1670032574
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1670032574
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1670032574
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_27
timestamp 1670032574
transform 1 0 3588 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1670032574
transform 1 0 4416 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1670032574
transform 1 0 5060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1670032574
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1670032574
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1670032574
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_69
timestamp 1670032574
transform 1 0 7452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_77
timestamp 1670032574
transform 1 0 8188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_85
timestamp 1670032574
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1670032574
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1670032574
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1670032574
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_134
timestamp 1670032574
transform 1 0 13432 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_146
timestamp 1670032574
transform 1 0 14536 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_156
timestamp 1670032574
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1670032574
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1670032574
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_185
timestamp 1670032574
transform 1 0 18124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_197
timestamp 1670032574
transform 1 0 19228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_209
timestamp 1670032574
transform 1 0 20332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1670032574
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_225
timestamp 1670032574
transform 1 0 21804 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_229
timestamp 1670032574
transform 1 0 22172 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_241
timestamp 1670032574
transform 1 0 23276 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_253
timestamp 1670032574
transform 1 0 24380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_259
timestamp 1670032574
transform 1 0 24932 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_263
timestamp 1670032574
transform 1 0 25300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_275
timestamp 1670032574
transform 1 0 26404 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1670032574
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1670032574
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_292
timestamp 1670032574
transform 1 0 27968 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 1670032574
transform 1 0 28520 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1670032574
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1670032574
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1670032574
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1670032574
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1670032574
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1670032574
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_65
timestamp 1670032574
transform 1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1670032574
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1670032574
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1670032574
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 1670032574
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_122
timestamp 1670032574
transform 1 0 12328 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 1670032574
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1670032574
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1670032574
transform 1 0 14904 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_174
timestamp 1670032574
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1670032574
transform 1 0 17940 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1670032574
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_197
timestamp 1670032574
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_202
timestamp 1670032574
transform 1 0 19688 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_214
timestamp 1670032574
transform 1 0 20792 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_222
timestamp 1670032574
transform 1 0 21528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_244
timestamp 1670032574
transform 1 0 23552 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_248
timestamp 1670032574
transform 1 0 23920 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1670032574
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1670032574
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_263
timestamp 1670032574
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_275
timestamp 1670032574
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_287
timestamp 1670032574
transform 1 0 27508 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_293
timestamp 1670032574
transform 1 0 28060 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp 1670032574
transform 1 0 28520 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1670032574
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_8
timestamp 1670032574
transform 1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_21
timestamp 1670032574
transform 1 0 3036 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_25
timestamp 1670032574
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_37
timestamp 1670032574
transform 1 0 4508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_48
timestamp 1670032574
transform 1 0 5520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_52
timestamp 1670032574
transform 1 0 5888 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1670032574
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1670032574
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_69
timestamp 1670032574
transform 1 0 7452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_90
timestamp 1670032574
transform 1 0 9384 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1670032574
transform 1 0 10120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_102
timestamp 1670032574
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1670032574
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1670032574
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_116
timestamp 1670032574
transform 1 0 11776 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_124
timestamp 1670032574
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_128
timestamp 1670032574
transform 1 0 12880 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_151
timestamp 1670032574
transform 1 0 14996 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1670032574
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1670032574
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_173
timestamp 1670032574
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_179
timestamp 1670032574
transform 1 0 17572 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_185
timestamp 1670032574
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_193
timestamp 1670032574
transform 1 0 18860 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_199
timestamp 1670032574
transform 1 0 19412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1670032574
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 1670032574
transform 1 0 20700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1670032574
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1670032574
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_237
timestamp 1670032574
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_241
timestamp 1670032574
transform 1 0 23276 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_263
timestamp 1670032574
transform 1 0 25300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1670032574
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1670032574
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1670032574
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1670032574
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1670032574
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1670032574
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1670032574
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1670032574
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_44
timestamp 1670032574
transform 1 0 5152 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_53
timestamp 1670032574
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_61
timestamp 1670032574
transform 1 0 6716 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 1670032574
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1670032574
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1670032574
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1670032574
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1670032574
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1670032574
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1670032574
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1670032574
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1670032574
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_168
timestamp 1670032574
transform 1 0 16560 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_176
timestamp 1670032574
transform 1 0 17296 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1670032574
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1670032574
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1670032574
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1670032574
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1670032574
transform 1 0 20424 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_214
timestamp 1670032574
transform 1 0 20792 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_222
timestamp 1670032574
transform 1 0 21528 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_234
timestamp 1670032574
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1670032574
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_253
timestamp 1670032574
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_257
timestamp 1670032574
transform 1 0 24748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_269
timestamp 1670032574
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_273
timestamp 1670032574
transform 1 0 26220 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1670032574
transform 1 0 28152 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_298
timestamp 1670032574
transform 1 0 28520 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1670032574
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1670032574
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1670032574
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1670032574
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1670032574
transform 1 0 4784 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1670032574
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1670032574
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_65
timestamp 1670032574
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_88
timestamp 1670032574
transform 1 0 9200 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_100
timestamp 1670032574
transform 1 0 10304 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1670032574
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1670032574
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1670032574
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1670032574
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1670032574
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1670032574
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1670032574
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1670032574
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_193
timestamp 1670032574
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1670032574
transform 1 0 19596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1670032574
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1670032574
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1670032574
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_249
timestamp 1670032574
transform 1 0 24012 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_254
timestamp 1670032574
transform 1 0 24472 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_266
timestamp 1670032574
transform 1 0 25576 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1670032574
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1670032574
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_281
timestamp 1670032574
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_291
timestamp 1670032574
transform 1 0 27876 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1670032574
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1670032574
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1670032574
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1670032574
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_41
timestamp 1670032574
transform 1 0 4876 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_62
timestamp 1670032574
transform 1 0 6808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp 1670032574
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1670032574
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1670032574
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1670032574
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1670032574
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1670032574
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1670032574
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1670032574
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1670032574
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1670032574
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1670032574
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_177
timestamp 1670032574
transform 1 0 17388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_185
timestamp 1670032574
transform 1 0 18124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1670032574
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1670032574
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1670032574
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_209
timestamp 1670032574
transform 1 0 20332 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_220
timestamp 1670032574
transform 1 0 21344 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_232
timestamp 1670032574
transform 1 0 22448 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_244
timestamp 1670032574
transform 1 0 23552 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1670032574
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_253
timestamp 1670032574
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_263
timestamp 1670032574
transform 1 0 25300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_275
timestamp 1670032574
transform 1 0 26404 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_287
timestamp 1670032574
transform 1 0 27508 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_293
timestamp 1670032574
transform 1 0 28060 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_298
timestamp 1670032574
transform 1 0 28520 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1670032574
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1670032574
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1670032574
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1670032574
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1670032574
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1670032574
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1670032574
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1670032574
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1670032574
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1670032574
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1670032574
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1670032574
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1670032574
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1670032574
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1670032574
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1670032574
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1670032574
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1670032574
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1670032574
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_201
timestamp 1670032574
transform 1 0 19596 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_213
timestamp 1670032574
transform 1 0 20700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1670032574
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1670032574
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_237
timestamp 1670032574
transform 1 0 22908 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1670032574
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1670032574
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1670032574
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1670032574
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1670032574
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1670032574
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1670032574
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_17
timestamp 1670032574
transform 1 0 2668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1670032574
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1670032574
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1670032574
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1670032574
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1670032574
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1670032574
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1670032574
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1670032574
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1670032574
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1670032574
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1670032574
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1670032574
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1670032574
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1670032574
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1670032574
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_165
timestamp 1670032574
transform 1 0 16284 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_180
timestamp 1670032574
transform 1 0 17664 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1670032574
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1670032574
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1670032574
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1670032574
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_229
timestamp 1670032574
transform 1 0 22172 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_241
timestamp 1670032574
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1670032574
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1670032574
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_265
timestamp 1670032574
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_271
timestamp 1670032574
transform 1 0 26036 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_292
timestamp 1670032574
transform 1 0 27968 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 1670032574
transform 1 0 28520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1670032574
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1670032574
transform 1 0 2116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_16
timestamp 1670032574
transform 1 0 2576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_27
timestamp 1670032574
transform 1 0 3588 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_31
timestamp 1670032574
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_43
timestamp 1670032574
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1670032574
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1670032574
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1670032574
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1670032574
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1670032574
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1670032574
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1670032574
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1670032574
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1670032574
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1670032574
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1670032574
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1670032574
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1670032574
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp 1670032574
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_190
timestamp 1670032574
transform 1 0 18584 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_202
timestamp 1670032574
transform 1 0 19688 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1670032574
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1670032574
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_225
timestamp 1670032574
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_235
timestamp 1670032574
transform 1 0 22724 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_239
timestamp 1670032574
transform 1 0 23092 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_251
timestamp 1670032574
transform 1 0 24196 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_263
timestamp 1670032574
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_275
timestamp 1670032574
transform 1 0 26404 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1670032574
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_281
timestamp 1670032574
transform 1 0 26956 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_291
timestamp 1670032574
transform 1 0 27876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1670032574
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1670032574
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_29
timestamp 1670032574
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_39
timestamp 1670032574
transform 1 0 4692 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_43
timestamp 1670032574
transform 1 0 5060 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_55
timestamp 1670032574
transform 1 0 6164 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_67
timestamp 1670032574
transform 1 0 7268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1670032574
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1670032574
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1670032574
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1670032574
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1670032574
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1670032574
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1670032574
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1670032574
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1670032574
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1670032574
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_165
timestamp 1670032574
transform 1 0 16284 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_174
timestamp 1670032574
transform 1 0 17112 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_186
timestamp 1670032574
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1670032574
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_197
timestamp 1670032574
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_214
timestamp 1670032574
transform 1 0 20792 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_226
timestamp 1670032574
transform 1 0 21896 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_230
timestamp 1670032574
transform 1 0 22264 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_242
timestamp 1670032574
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1670032574
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1670032574
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1670032574
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_269
timestamp 1670032574
transform 1 0 25852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_272
timestamp 1670032574
transform 1 0 26128 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_294
timestamp 1670032574
transform 1 0 28152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_298
timestamp 1670032574
transform 1 0 28520 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1670032574
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1670032574
transform 1 0 1748 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_28
timestamp 1670032574
transform 1 0 3680 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_40
timestamp 1670032574
transform 1 0 4784 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1670032574
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1670032574
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1670032574
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1670032574
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1670032574
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1670032574
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1670032574
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1670032574
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1670032574
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1670032574
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1670032574
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1670032574
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1670032574
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1670032574
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1670032574
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_193
timestamp 1670032574
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1670032574
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_225
timestamp 1670032574
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_246
timestamp 1670032574
transform 1 0 23736 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_251
timestamp 1670032574
transform 1 0 24196 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_263
timestamp 1670032574
transform 1 0 25300 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_269
timestamp 1670032574
transform 1 0 25852 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1670032574
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_281
timestamp 1670032574
transform 1 0 26956 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_285
timestamp 1670032574
transform 1 0 27324 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_293
timestamp 1670032574
transform 1 0 28060 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1670032574
transform 1 0 28520 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1670032574
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1670032574
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1670032574
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1670032574
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1670032574
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1670032574
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1670032574
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1670032574
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1670032574
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1670032574
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1670032574
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1670032574
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1670032574
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1670032574
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1670032574
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1670032574
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1670032574
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1670032574
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1670032574
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1670032574
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1670032574
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1670032574
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_205
timestamp 1670032574
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1670032574
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_221
timestamp 1670032574
transform 1 0 21436 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_229
timestamp 1670032574
transform 1 0 22172 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1670032574
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1670032574
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_261
timestamp 1670032574
transform 1 0 25116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_283
timestamp 1670032574
transform 1 0 27140 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_294
timestamp 1670032574
transform 1 0 28152 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_298
timestamp 1670032574
transform 1 0 28520 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 1670032574
transform 1 0 1380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1670032574
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1670032574
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1670032574
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1670032574
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1670032574
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1670032574
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1670032574
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1670032574
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1670032574
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1670032574
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1670032574
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1670032574
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1670032574
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1670032574
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1670032574
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1670032574
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1670032574
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1670032574
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1670032574
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1670032574
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1670032574
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1670032574
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1670032574
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1670032574
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_250
timestamp 1670032574
transform 1 0 24104 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1670032574
transform 1 0 25208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_266
timestamp 1670032574
transform 1 0 25576 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1670032574
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1670032574
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1670032574
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1670032574
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1670032574
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1670032574
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1670032574
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1670032574
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1670032574
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1670032574
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1670032574
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1670032574
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1670032574
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1670032574
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1670032574
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1670032574
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1670032574
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1670032574
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1670032574
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1670032574
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1670032574
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1670032574
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1670032574
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1670032574
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1670032574
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1670032574
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1670032574
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1670032574
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1670032574
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1670032574
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1670032574
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1670032574
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1670032574
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1670032574
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_289
timestamp 1670032574
transform 1 0 27692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1670032574
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1670032574
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1670032574
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1670032574
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1670032574
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1670032574
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1670032574
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1670032574
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1670032574
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1670032574
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1670032574
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1670032574
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1670032574
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1670032574
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1670032574
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1670032574
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1670032574
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1670032574
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1670032574
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1670032574
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1670032574
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1670032574
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1670032574
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1670032574
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1670032574
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1670032574
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1670032574
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1670032574
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1670032574
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1670032574
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1670032574
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1670032574
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_293
timestamp 1670032574
transform 1 0 28060 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_298
timestamp 1670032574
transform 1 0 28520 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1670032574
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1670032574
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1670032574
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1670032574
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1670032574
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1670032574
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1670032574
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1670032574
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1670032574
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1670032574
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1670032574
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1670032574
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1670032574
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1670032574
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1670032574
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1670032574
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1670032574
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1670032574
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1670032574
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1670032574
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1670032574
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1670032574
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1670032574
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1670032574
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1670032574
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1670032574
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1670032574
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1670032574
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1670032574
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1670032574
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp 1670032574
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1670032574
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1670032574
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1670032574
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1670032574
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1670032574
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1670032574
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1670032574
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1670032574
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1670032574
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1670032574
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1670032574
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1670032574
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1670032574
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1670032574
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1670032574
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1670032574
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1670032574
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1670032574
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1670032574
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1670032574
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1670032574
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1670032574
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1670032574
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1670032574
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1670032574
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1670032574
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1670032574
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1670032574
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1670032574
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1670032574
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1670032574
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1670032574
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1670032574
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1670032574
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1670032574
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1670032574
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1670032574
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1670032574
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1670032574
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1670032574
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1670032574
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1670032574
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1670032574
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1670032574
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1670032574
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1670032574
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1670032574
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1670032574
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1670032574
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1670032574
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1670032574
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1670032574
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1670032574
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1670032574
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1670032574
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1670032574
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1670032574
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1670032574
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1670032574
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1670032574
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1670032574
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1670032574
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1670032574
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp 1670032574
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1670032574
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1670032574
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1670032574
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1670032574
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1670032574
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1670032574
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1670032574
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1670032574
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1670032574
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1670032574
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1670032574
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1670032574
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1670032574
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1670032574
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1670032574
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1670032574
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1670032574
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1670032574
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1670032574
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1670032574
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1670032574
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1670032574
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1670032574
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1670032574
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1670032574
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1670032574
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1670032574
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1670032574
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1670032574
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1670032574
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1670032574
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1670032574
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1670032574
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1670032574
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1670032574
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1670032574
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1670032574
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1670032574
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1670032574
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1670032574
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1670032574
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1670032574
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1670032574
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1670032574
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1670032574
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1670032574
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1670032574
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1670032574
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1670032574
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1670032574
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1670032574
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1670032574
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1670032574
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1670032574
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1670032574
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1670032574
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1670032574
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1670032574
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1670032574
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1670032574
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1670032574
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1670032574
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1670032574
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1670032574
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_293
timestamp 1670032574
transform 1 0 28060 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_298
timestamp 1670032574
transform 1 0 28520 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1670032574
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1670032574
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1670032574
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1670032574
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1670032574
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1670032574
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1670032574
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1670032574
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1670032574
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1670032574
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1670032574
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1670032574
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1670032574
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1670032574
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1670032574
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1670032574
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1670032574
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1670032574
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1670032574
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1670032574
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1670032574
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1670032574
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1670032574
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1670032574
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1670032574
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1670032574
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1670032574
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1670032574
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1670032574
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1670032574
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1670032574
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1670032574
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_3
timestamp 1670032574
transform 1 0 1380 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_8
timestamp 1670032574
transform 1 0 1840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1670032574
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1670032574
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1670032574
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp 1670032574
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_57
timestamp 1670032574
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_69
timestamp 1670032574
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1670032574
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1670032574
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1670032574
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp 1670032574
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_113
timestamp 1670032574
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_125
timestamp 1670032574
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1670032574
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1670032574
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1670032574
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1670032574
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_169
timestamp 1670032574
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_181
timestamp 1670032574
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1670032574
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1670032574
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1670032574
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp 1670032574
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1670032574
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1670032574
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1670032574
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1670032574
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1670032574
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_277
timestamp 1670032574
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_281
timestamp 1670032574
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_293
timestamp 1670032574
transform 1 0 28060 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_298
timestamp 1670032574
transform 1 0 28520 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1670032574
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1670032574
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1670032574
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1670032574
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1670032574
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1670032574
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1670032574
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1670032574
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1670032574
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1670032574
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1670032574
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1670032574
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1670032574
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1670032574
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1670032574
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1670032574
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1670032574
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1670032574
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1670032574
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1670032574
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1670032574
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1670032574
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1670032574
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1670032574
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1670032574
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1670032574
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1670032574
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1670032574
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1670032574
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1670032574
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1670032574
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1670032574
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1670032574
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1670032574
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1670032574
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1670032574
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1670032574
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1670032574
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1670032574
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1670032574
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1670032574
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1670032574
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1670032574
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1670032574
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1670032574
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1670032574
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1670032574
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1670032574
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1670032574
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1670032574
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1670032574
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1670032574
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1670032574
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1670032574
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1670032574
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1670032574
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1670032574
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1670032574
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1670032574
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1670032574
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1670032574
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1670032574
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1670032574
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1670032574
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1670032574
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1670032574
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1670032574
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1670032574
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1670032574
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1670032574
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1670032574
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1670032574
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1670032574
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1670032574
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1670032574
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1670032574
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1670032574
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1670032574
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1670032574
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1670032574
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1670032574
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1670032574
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1670032574
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1670032574
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1670032574
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1670032574
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1670032574
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1670032574
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1670032574
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1670032574
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1670032574
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1670032574
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1670032574
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1670032574
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1670032574
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1670032574
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1670032574
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1670032574
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1670032574
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1670032574
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1670032574
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1670032574
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1670032574
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1670032574
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1670032574
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1670032574
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1670032574
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1670032574
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1670032574
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1670032574
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1670032574
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1670032574
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1670032574
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1670032574
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1670032574
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1670032574
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1670032574
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1670032574
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1670032574
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1670032574
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1670032574
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1670032574
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1670032574
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1670032574
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1670032574
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1670032574
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1670032574
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1670032574
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1670032574
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1670032574
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1670032574
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1670032574
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1670032574
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1670032574
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1670032574
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1670032574
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1670032574
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1670032574
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1670032574
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1670032574
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1670032574
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1670032574
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1670032574
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1670032574
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1670032574
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1670032574
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1670032574
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1670032574
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1670032574
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1670032574
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1670032574
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1670032574
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1670032574
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1670032574
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1670032574
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1670032574
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1670032574
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1670032574
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1670032574
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1670032574
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1670032574
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1670032574
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1670032574
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1670032574
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1670032574
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1670032574
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1670032574
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1670032574
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1670032574
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1670032574
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1670032574
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1670032574
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1670032574
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1670032574
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1670032574
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1670032574
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1670032574
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1670032574
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1670032574
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1670032574
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1670032574
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1670032574
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1670032574
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1670032574
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1670032574
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1670032574
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1670032574
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1670032574
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1670032574
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1670032574
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1670032574
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1670032574
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1670032574
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1670032574
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1670032574
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1670032574
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1670032574
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1670032574
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1670032574
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1670032574
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1670032574
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1670032574
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1670032574
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1670032574
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1670032574
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1670032574
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1670032574
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1670032574
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1670032574
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1670032574
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1670032574
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1670032574
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1670032574
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1670032574
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1670032574
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1670032574
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1670032574
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1670032574
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1670032574
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1670032574
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1670032574
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1670032574
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1670032574
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1670032574
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1670032574
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1670032574
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1670032574
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1670032574
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1670032574
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1670032574
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1670032574
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1670032574
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1670032574
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1670032574
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1670032574
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1670032574
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1670032574
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1670032574
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1670032574
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1670032574
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1670032574
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1670032574
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1670032574
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1670032574
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1670032574
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1670032574
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1670032574
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1670032574
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1670032574
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1670032574
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1670032574
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1670032574
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1670032574
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1670032574
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1670032574
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1670032574
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1670032574
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1670032574
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1670032574
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1670032574
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1670032574
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1670032574
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1670032574
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1670032574
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1670032574
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1670032574
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1670032574
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1670032574
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1670032574
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1670032574
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1670032574
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1670032574
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1670032574
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1670032574
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1670032574
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1670032574
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1670032574
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1670032574
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1670032574
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1670032574
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1670032574
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1670032574
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1670032574
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1670032574
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1670032574
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1670032574
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1670032574
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1670032574
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1670032574
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1670032574
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1670032574
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1670032574
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1670032574
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1670032574
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1670032574
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1670032574
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1670032574
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1670032574
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1670032574
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1670032574
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1670032574
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1670032574
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1670032574
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1670032574
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1670032574
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1670032574
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1670032574
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1670032574
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1670032574
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1670032574
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1670032574
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1670032574
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1670032574
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1670032574
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1670032574
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1670032574
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1670032574
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1670032574
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1670032574
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1670032574
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1670032574
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1670032574
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1670032574
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1670032574
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1670032574
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1670032574
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1670032574
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1670032574
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1670032574
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1670032574
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1670032574
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1670032574
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1670032574
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1670032574
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1670032574
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1670032574
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1670032574
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1670032574
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_4  _143_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 16744 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__or3b_1  _144_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 17388 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _145_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 15548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _146_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 14444 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _147_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 17296 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _148_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 17572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _149_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 21620 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _150_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 23092 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _151_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _152_
timestamp 1670032574
transform 1 0 22080 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1670032574
transform -1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _154_
timestamp 1670032574
transform -1 0 25760 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1670032574
transform -1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _156_
timestamp 1670032574
transform -1 0 25300 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1670032574
transform -1 0 24932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _158_
timestamp 1670032574
transform -1 0 24012 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1670032574
transform -1 0 23736 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp 1670032574
transform -1 0 25484 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1670032574
transform -1 0 25208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp 1670032574
transform -1 0 25576 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1670032574
transform -1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _164_
timestamp 1670032574
transform 1 0 24472 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1670032574
transform -1 0 24748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 1670032574
transform 1 0 24472 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1670032574
transform 1 0 23920 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _168_
timestamp 1670032574
transform 1 0 21896 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1670032574
transform -1 0 22264 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _170_
timestamp 1670032574
transform 1 0 19964 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1670032574
transform -1 0 20332 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _172_
timestamp 1670032574
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1670032574
transform -1 0 17112 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _174_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 22816 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _175_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 22264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _176_
timestamp 1670032574
transform -1 0 22172 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _177_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 21344 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _178_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 20424 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _179_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 18308 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _180_
timestamp 1670032574
transform -1 0 18860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _181_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 17572 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _182_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 17940 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _183_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 19320 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _184_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 18308 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _185_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 19872 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _186_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 19320 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _187_
timestamp 1670032574
transform -1 0 21436 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _188_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 21436 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _189_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 20792 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1670032574
transform -1 0 22448 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _191_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 21896 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _192_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 20792 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1670032574
transform 1 0 22448 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _194_
timestamp 1670032574
transform -1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _195_
timestamp 1670032574
transform -1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _196_
timestamp 1670032574
transform 1 0 20976 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _197_
timestamp 1670032574
transform -1 0 22356 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _198_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 22816 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _199_
timestamp 1670032574
transform 1 0 20332 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1670032574
transform 1 0 20516 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _201_
timestamp 1670032574
transform -1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _202_
timestamp 1670032574
transform -1 0 21620 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _203_
timestamp 1670032574
transform -1 0 19780 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _204_
timestamp 1670032574
transform 1 0 21896 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _205_
timestamp 1670032574
transform 1 0 19964 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1670032574
transform -1 0 22172 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _207_
timestamp 1670032574
transform -1 0 19504 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _208_
timestamp 1670032574
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _209_
timestamp 1670032574
transform 1 0 20884 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _210_
timestamp 1670032574
transform 1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _211_
timestamp 1670032574
transform -1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _212_
timestamp 1670032574
transform 1 0 19504 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _213_
timestamp 1670032574
transform 1 0 18216 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1670032574
transform 1 0 18216 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _215_
timestamp 1670032574
transform 1 0 17112 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _216_
timestamp 1670032574
transform -1 0 17940 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1670032574
transform 1 0 16284 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _218_
timestamp 1670032574
transform -1 0 6716 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _219_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 6440 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1670032574
transform -1 0 7268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1670032574
transform 1 0 4600 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _222_
timestamp 1670032574
transform 1 0 5152 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _223_
timestamp 1670032574
transform -1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _224_
timestamp 1670032574
transform 1 0 6808 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _225_
timestamp 1670032574
transform 1 0 8280 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1670032574
transform 1 0 10120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _227_
timestamp 1670032574
transform 1 0 4692 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _228_
timestamp 1670032574
transform 1 0 5520 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1670032574
transform 1 0 7268 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _230_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 11132 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1670032574
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _232_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 18124 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _233_
timestamp 1670032574
transform 1 0 5060 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _234_
timestamp 1670032574
transform 1 0 5612 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _235_
timestamp 1670032574
transform 1 0 6440 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _236_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 6992 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _237_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 8464 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _238_
timestamp 1670032574
transform -1 0 16376 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _239_
timestamp 1670032574
transform -1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _240_
timestamp 1670032574
transform 1 0 8648 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _241_
timestamp 1670032574
transform 1 0 9384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _242_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 5612 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _243_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 6900 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1670032574
transform 1 0 10488 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _245_
timestamp 1670032574
transform 1 0 11684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _246_
timestamp 1670032574
transform 1 0 9292 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _247_
timestamp 1670032574
transform 1 0 11040 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _248_
timestamp 1670032574
transform 1 0 11592 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1670032574
transform -1 0 12144 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _250_
timestamp 1670032574
transform -1 0 7084 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _251_
timestamp 1670032574
transform -1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _252_
timestamp 1670032574
transform 1 0 6624 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1670032574
transform -1 0 7544 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _254_
timestamp 1670032574
transform 1 0 11500 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _255_
timestamp 1670032574
transform 1 0 12972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _256_
timestamp 1670032574
transform 1 0 12696 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1670032574
transform -1 0 13616 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _258_
timestamp 1670032574
transform -1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1670032574
transform 1 0 25392 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1670032574
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _261_
timestamp 1670032574
transform 1 0 27232 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1670032574
transform 1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _263_
timestamp 1670032574
transform 1 0 27232 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1670032574
transform 1 0 27048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _265_
timestamp 1670032574
transform 1 0 27232 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1670032574
transform 1 0 27048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _267_
timestamp 1670032574
transform 1 0 27232 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1670032574
transform 1 0 27048 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _269_
timestamp 1670032574
transform 1 0 27232 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1670032574
transform 1 0 27048 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _271_
timestamp 1670032574
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 1670032574
transform -1 0 26772 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1670032574
transform 1 0 27048 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1670032574
transform 1 0 26496 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1670032574
transform 1 0 27048 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1670032574
transform 1 0 26496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _277_
timestamp 1670032574
transform -1 0 24104 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp 1670032574
transform 1 0 23920 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _279_
timestamp 1670032574
transform 1 0 25944 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1670032574
transform 1 0 25668 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _281_
timestamp 1670032574
transform 1 0 27324 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1670032574
transform 1 0 27048 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _283_
timestamp 1670032574
transform -1 0 11040 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _284_
timestamp 1670032574
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _285_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 9108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_4  _286_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 11040 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp 1670032574
transform 1 0 2484 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1670032574
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _289_
timestamp 1670032574
transform 1 0 2576 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1670032574
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _291_
timestamp 1670032574
transform 1 0 2208 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1670032574
transform 1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1670032574
transform 1 0 2208 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1670032574
transform -1 0 2484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1670032574
transform 1 0 3864 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1670032574
transform 1 0 2392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1670032574
transform 1 0 2760 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1670032574
transform 1 0 2300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1670032574
transform -1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _300_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _301_
timestamp 1670032574
transform -1 0 16100 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _302_
timestamp 1670032574
transform -1 0 15088 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _303_
timestamp 1670032574
transform -1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _304_
timestamp 1670032574
transform -1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _305_
timestamp 1670032574
transform -1 0 9752 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _306_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 3772 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _307_
timestamp 1670032574
transform 1 0 3864 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _308_
timestamp 1670032574
transform 1 0 3680 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _309_
timestamp 1670032574
transform 1 0 5244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _310_
timestamp 1670032574
transform 1 0 4048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _311_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 16192 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _312_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 12236 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _313_
timestamp 1670032574
transform 1 0 9660 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _314_
timestamp 1670032574
transform -1 0 8188 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _315_
timestamp 1670032574
transform -1 0 8096 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _316_
timestamp 1670032574
transform -1 0 8004 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _317_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 14168 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _318_
timestamp 1670032574
transform 1 0 12420 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _319_
timestamp 1670032574
transform 1 0 15732 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _320_
timestamp 1670032574
transform 1 0 17572 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _321_
timestamp 1670032574
transform -1 0 15732 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _322_
timestamp 1670032574
transform 1 0 16744 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _323_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 15088 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _324_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _325_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 24840 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1670032574
transform 1 0 26680 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 1670032574
transform 1 0 26588 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _328_
timestamp 1670032574
transform 1 0 26496 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _329_
timestamp 1670032574
transform 1 0 26496 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _330_
timestamp 1670032574
transform 1 0 26588 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _331_
timestamp 1670032574
transform 1 0 26588 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _332_
timestamp 1670032574
transform 1 0 26312 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1670032574
transform 1 0 26128 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _334_
timestamp 1670032574
transform 1 0 22356 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _335_
timestamp 1670032574
transform 1 0 25300 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _336_
timestamp 1670032574
transform 1 0 26312 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _337_
timestamp 1670032574
transform 1 0 1656 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _338_
timestamp 1670032574
transform 1 0 1656 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 1670032574
transform 1 0 1472 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _340_
timestamp 1670032574
transform -1 0 3312 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _341_
timestamp 1670032574
transform 1 0 1748 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _342_
timestamp 1670032574
transform 1 0 1840 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _343_
timestamp 1670032574
transform 1 0 19320 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _344_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 19596 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _345_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 18768 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _346_
timestamp 1670032574
transform 1 0 22356 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _347_
timestamp 1670032574
transform 1 0 21528 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _348_
timestamp 1670032574
transform 1 0 20056 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _349_
timestamp 1670032574
transform 1 0 19964 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _350_
timestamp 1670032574
transform 1 0 22448 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _351_
timestamp 1670032574
transform 1 0 21712 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _352_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 18124 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _353_
timestamp 1670032574
transform 1 0 19780 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _354_
timestamp 1670032574
transform 1 0 17756 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _355_
timestamp 1670032574
transform 1 0 15180 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _356_
timestamp 1670032574
transform 1 0 22264 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _357_
timestamp 1670032574
transform 1 0 21344 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _358_
timestamp 1670032574
transform -1 0 26588 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _359_
timestamp 1670032574
transform -1 0 26312 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _360_
timestamp 1670032574
transform -1 0 24196 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _361_
timestamp 1670032574
transform -1 0 26220 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _362_
timestamp 1670032574
transform -1 0 26312 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _363_
timestamp 1670032574
transform 1 0 23460 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _364_
timestamp 1670032574
transform 1 0 23276 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _365_
timestamp 1670032574
transform -1 0 23736 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _366_
timestamp 1670032574
transform 1 0 19136 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _367_
timestamp 1670032574
transform -1 0 18584 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _368_
timestamp 1670032574
transform 1 0 9016 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _369_
timestamp 1670032574
transform -1 0 4324 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _370_
timestamp 1670032574
transform 1 0 3128 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _371_
timestamp 1670032574
transform -1 0 3588 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _372_
timestamp 1670032574
transform 1 0 4968 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _373_
timestamp 1670032574
transform -1 0 4784 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _374_
timestamp 1670032574
transform 1 0 11592 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _375_
timestamp 1670032574
transform 1 0 10488 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _376_
timestamp 1670032574
transform 1 0 7544 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _377_
timestamp 1670032574
transform 1 0 7544 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _378_
timestamp 1670032574
transform 1 0 7360 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _379_
timestamp 1670032574
transform -1 0 14996 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _380_
timestamp 1670032574
transform 1 0 15732 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _381_
timestamp 1670032574
transform 1 0 14904 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _382_
timestamp 1670032574
transform -1 0 19596 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 14168 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1670032574
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1670032574
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1670032574
transform -1 0 7084 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1670032574
transform 1 0 10396 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1670032574
transform 1 0 18216 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1670032574
transform 1 0 20792 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1670032574
transform 1 0 20792 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1670032574
transform 1 0 20792 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 12788 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref
timestamp 1670032574
transform 1 0 13340 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1670032574
transform 1 0 6624 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1670032574
transform -1 0 7360 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1670032574
transform 1 0 7268 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref
timestamp 1670032574
transform 1 0 7544 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1670032574
transform 1 0 9752 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1670032574
transform 1 0 12788 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1670032574
transform -1 0 10856 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1670032574
transform 1 0 13432 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1670032574
transform -1 0 10212 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1670032574
transform -1 0 13248 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1670032574
transform 1 0 9108 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1670032574
transform 1 0 12788 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1670032574
transform 1 0 4232 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1670032574
transform 1 0 13340 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1670032574
transform 1 0 4876 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1670032574
transform 1 0 13984 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1670032574
transform 1 0 4232 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1670032574
transform -1 0 13800 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1670032574
transform 1 0 4232 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1670032574
transform -1 0 13800 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1670032574
transform 1 0 4876 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1670032574
transform 1 0 12696 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1670032574
transform 1 0 4876 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1670032574
transform 1 0 14628 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1670032574
transform 1 0 4232 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref
timestamp 1670032574
transform -1 0 14628 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1670032574
transform 1 0 4232 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1670032574
transform -1 0 14628 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1670032574
transform 1 0 6624 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1670032574
transform 1 0 10672 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1670032574
transform 1 0 7268 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1670032574
transform 1 0 11316 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1670032574
transform -1 0 7084 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1670032574
transform -1 0 11132 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1670032574
transform 1 0 6624 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1670032574
transform 1 0 10672 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1670032574
transform 1 0 5336 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1670032574
transform -1 0 9844 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1670032574
transform 1 0 5704 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1670032574
transform 1 0 10672 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1670032574
transform 1 0 5704 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref
timestamp 1670032574
transform 1 0 11960 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1670032574
transform -1 0 7728 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1670032574
transform 1 0 12236 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1670032574
transform 1 0 7268 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1670032574
transform 1 0 11960 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1670032574
transform 1 0 7912 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1670032574
transform 1 0 10672 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1670032574
transform 1 0 6624 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1670032574
transform 1 0 10028 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1670032574
transform 1 0 5980 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1670032574
transform 1 0 10028 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1670032574
transform 1 0 7268 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1670032574
transform 1 0 10028 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1670032574
transform 1 0 7268 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1670032574
transform 1 0 12880 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1670032574
transform 1 0 7912 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1670032574
transform 1 0 11592 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1670032574
transform 1 0 6624 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1670032574
transform 1 0 11316 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1670032574
transform 1 0 8740 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  dac.vdac_single.einvp_batch\[0\].pupd_30 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  dac.vdac_single.einvp_batch\[0\].vref_29
timestamp 1670032574
transform -1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  dac.vdac_single.einvp_batch\[0\].vref
timestamp 1670032574
transform -1 0 4508 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__einvp_1  dcdc
timestamp 1670032574
transform 1 0 13340 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1670032574
transform -1 0 9568 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1670032574
transform -1 0 3404 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1670032574
transform 1 0 22448 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1670032574
transform -1 0 20608 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1670032574
transform 1 0 24472 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 17204 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 1670032574
transform -1 0 4048 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1670032574
transform 1 0 11592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1670032574
transform 1 0 18768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  inv1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 13708 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  inv2
timestamp 1670032574
transform -1 0 12880 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1670032574
transform 1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1670032574
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1670032574
transform 1 0 28152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1670032574
transform 1 0 28152 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1670032574
transform 1 0 28152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1670032574
transform 1 0 28152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1670032574
transform 1 0 28152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1670032574
transform 1 0 28152 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1670032574
transform 1 0 28152 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1670032574
transform 1 0 28152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1670032574
transform 1 0 28152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1670032574
transform 1 0 28152 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1670032574
transform 1 0 28152 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1670032574
transform -1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1670032574
transform -1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1670032574
transform -1 0 1840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1670032574
transform -1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1670032574
transform -1 0 1840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1670032574
transform -1 0 1840 0 1 27200
box -38 -48 406 592
<< labels >>
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 conversion_finished_out
port 1 nsew signal tristate
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 rst_n
port 2 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 start_conv_in
port 3 nsew signal input
flabel metal3 s 29200 1368 30000 1488 0 FreeSans 480 0 0 0 tick_result_out[0]
port 4 nsew signal tristate
flabel metal3 s 29200 25848 30000 25968 0 FreeSans 480 0 0 0 tick_result_out[10]
port 5 nsew signal tristate
flabel metal3 s 29200 28296 30000 28416 0 FreeSans 480 0 0 0 tick_result_out[11]
port 6 nsew signal tristate
flabel metal3 s 29200 3816 30000 3936 0 FreeSans 480 0 0 0 tick_result_out[1]
port 7 nsew signal tristate
flabel metal3 s 29200 6264 30000 6384 0 FreeSans 480 0 0 0 tick_result_out[2]
port 8 nsew signal tristate
flabel metal3 s 29200 8712 30000 8832 0 FreeSans 480 0 0 0 tick_result_out[3]
port 9 nsew signal tristate
flabel metal3 s 29200 11160 30000 11280 0 FreeSans 480 0 0 0 tick_result_out[4]
port 10 nsew signal tristate
flabel metal3 s 29200 13608 30000 13728 0 FreeSans 480 0 0 0 tick_result_out[5]
port 11 nsew signal tristate
flabel metal3 s 29200 16056 30000 16176 0 FreeSans 480 0 0 0 tick_result_out[6]
port 12 nsew signal tristate
flabel metal3 s 29200 18504 30000 18624 0 FreeSans 480 0 0 0 tick_result_out[7]
port 13 nsew signal tristate
flabel metal3 s 29200 20952 30000 21072 0 FreeSans 480 0 0 0 tick_result_out[8]
port 14 nsew signal tristate
flabel metal3 s 29200 23400 30000 23520 0 FreeSans 480 0 0 0 tick_result_out[9]
port 15 nsew signal tristate
flabel metal4 s 3344 2128 3664 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 8144 2128 8464 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 12944 2128 13264 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 17744 2128 18064 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 22544 2128 22864 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 27344 2128 27664 27792 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 vdac_result_out[0]
port 17 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 vdac_result_out[1]
port 18 nsew signal tristate
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 vdac_result_out[2]
port 19 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 vdac_result_out[3]
port 20 nsew signal tristate
flabel metal3 s 0 22176 800 22296 0 FreeSans 480 0 0 0 vdac_result_out[4]
port 21 nsew signal tristate
flabel metal3 s 0 27072 800 27192 0 FreeSans 480 0 0 0 vdac_result_out[5]
port 22 nsew signal tristate
flabel metal4 s 5744 2128 6064 27792 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
flabel metal4 s 10544 2128 10864 27792 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
flabel metal4 s 15344 2128 15664 27792 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
flabel metal4 s 20144 2128 20464 27792 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
flabel metal4 s 24944 2128 25264 27792 0 FreeSans 1920 90 0 0 vssd1
port 23 nsew ground bidirectional
rlabel metal1 14996 27744 14996 27744 0 vccd1
rlabel metal1 14996 27200 14996 27200 0 vssd1
rlabel metal1 27002 6630 27002 6630 0 _000_
rlabel metal2 26818 9180 26818 9180 0 _001_
rlabel metal2 26818 11356 26818 11356 0 _002_
rlabel metal2 26910 13532 26910 13532 0 _003_
rlabel metal2 26910 15708 26910 15708 0 _004_
rlabel metal2 26634 17884 26634 17884 0 _005_
rlabel metal2 26450 20060 26450 20060 0 _006_
rlabel metal2 23966 21930 23966 21930 0 _007_
rlabel metal1 25661 22202 25661 22202 0 _008_
rlabel metal2 26634 21148 26634 21148 0 _009_
rlabel metal2 2254 3298 2254 3298 0 _010_
rlabel metal2 1978 8092 1978 8092 0 _011_
rlabel metal2 1794 13022 1794 13022 0 _012_
rlabel metal2 2898 17884 2898 17884 0 _013_
rlabel metal1 2254 20026 2254 20026 0 _014_
rlabel metal1 2254 20570 2254 20570 0 _015_
rlabel metal1 19366 3434 19366 3434 0 _016_
rlabel metal2 9614 13090 9614 13090 0 _017_
rlabel metal1 3910 12614 3910 12614 0 _018_
rlabel metal2 3910 14756 3910 14756 0 _019_
rlabel metal1 3505 15674 3505 15674 0 _020_
rlabel metal2 5290 18258 5290 18258 0 _021_
rlabel metal1 4278 17850 4278 17850 0 _022_
rlabel metal1 11776 14858 11776 14858 0 _023_
rlabel metal1 10810 16456 10810 16456 0 _024_
rlabel metal2 7866 15470 7866 15470 0 _025_
rlabel metal1 7682 17238 7682 17238 0 _026_
rlabel metal2 7406 17374 7406 17374 0 _027_
rlabel metal1 14398 16762 14398 16762 0 _028_
rlabel metal2 16790 9690 16790 9690 0 _029_
rlabel metal2 15134 14042 15134 14042 0 _030_
rlabel metal2 19274 11152 19274 11152 0 _031_
rlabel metal2 25162 3672 25162 3672 0 _032_
rlabel metal1 27048 3706 27048 3706 0 _033_
rlabel metal1 13846 13294 13846 13294 0 _034_
rlabel metal2 16790 13090 16790 13090 0 _035_
rlabel metal2 15410 13702 15410 13702 0 _036_
rlabel metal2 17526 14144 17526 14144 0 _037_
rlabel metal1 20700 20978 20700 20978 0 _038_
rlabel metal1 24886 5746 24886 5746 0 _039_
rlabel metal2 23230 4284 23230 4284 0 _040_
rlabel metal2 22126 4284 22126 4284 0 _041_
rlabel metal2 25714 6324 25714 6324 0 _042_
rlabel metal1 25070 8602 25070 8602 0 _043_
rlabel metal2 23966 11254 23966 11254 0 _044_
rlabel metal2 25438 12852 25438 12852 0 _045_
rlabel metal2 25530 15606 25530 15606 0 _046_
rlabel metal2 24518 17204 24518 17204 0 _047_
rlabel metal1 24334 18734 24334 18734 0 _048_
rlabel metal1 21988 20570 21988 20570 0 _049_
rlabel metal2 20010 21556 20010 21556 0 _050_
rlabel metal2 16882 20468 16882 20468 0 _051_
rlabel metal1 22770 8058 22770 8058 0 _052_
rlabel metal1 21206 17612 21206 17612 0 _053_
rlabel metal1 20608 17578 20608 17578 0 _054_
rlabel metal1 20470 17646 20470 17646 0 _055_
rlabel metal1 19044 17646 19044 17646 0 _056_
rlabel metal1 23506 22508 23506 22508 0 _057_
rlabel metal1 25576 2958 25576 2958 0 _058_
rlabel metal1 16974 13294 16974 13294 0 _059_
rlabel metal1 18998 17034 18998 17034 0 _060_
rlabel metal1 21068 17170 21068 17170 0 _061_
rlabel metal1 19458 5678 19458 5678 0 _062_
rlabel metal2 20838 6562 20838 6562 0 _063_
rlabel metal1 21268 6698 21268 6698 0 _064_
rlabel metal2 21666 6460 21666 6460 0 _065_
rlabel metal1 21574 7514 21574 7514 0 _066_
rlabel metal1 22678 8500 22678 8500 0 _067_
rlabel metal1 20884 10710 20884 10710 0 _068_
rlabel metal1 20562 12648 20562 12648 0 _069_
rlabel metal1 22034 13702 22034 13702 0 _070_
rlabel metal1 21817 12954 21817 12954 0 _071_
rlabel metal1 20792 12614 20792 12614 0 _072_
rlabel metal1 21758 13974 21758 13974 0 _073_
rlabel metal1 20286 17238 20286 17238 0 _074_
rlabel metal2 21942 15232 21942 15232 0 _075_
rlabel metal2 20562 15878 20562 15878 0 _076_
rlabel metal1 18906 15062 18906 15062 0 _077_
rlabel metal1 20884 17170 20884 17170 0 _078_
rlabel metal1 20654 17272 20654 17272 0 _079_
rlabel metal1 19090 17306 19090 17306 0 _080_
rlabel metal2 18814 17850 18814 17850 0 _081_
rlabel metal1 17572 16966 17572 16966 0 _082_
rlabel metal2 16514 17204 16514 17204 0 _083_
rlabel metal2 6302 15946 6302 15946 0 _084_
rlabel metal1 6992 14314 6992 14314 0 _085_
rlabel metal1 5106 15878 5106 15878 0 _086_
rlabel metal1 5612 10642 5612 10642 0 _087_
rlabel metal1 7866 14790 7866 14790 0 _088_
rlabel metal1 9108 11118 9108 11118 0 _089_
rlabel metal1 5014 12818 5014 12818 0 _090_
rlabel metal1 6394 12818 6394 12818 0 _091_
rlabel metal2 12282 12988 12282 12988 0 _092_
rlabel metal1 18492 3434 18492 3434 0 _093_
rlabel metal1 5566 16966 5566 16966 0 _094_
rlabel metal2 6578 14382 6578 14382 0 _095_
rlabel metal2 6762 13260 6762 13260 0 _096_
rlabel metal1 7958 8500 7958 8500 0 _097_
rlabel metal2 15962 10030 15962 10030 0 _098_
rlabel metal2 13938 10880 13938 10880 0 _099_
rlabel metal1 9292 7854 9292 7854 0 _100_
rlabel metal1 6670 9996 6670 9996 0 _101_
rlabel metal1 11362 8942 11362 8942 0 _102_
rlabel metal2 11086 10914 11086 10914 0 _103_
rlabel metal2 12006 10132 12006 10132 0 _104_
rlabel metal1 6440 12614 6440 12614 0 _105_
rlabel metal1 7176 11730 7176 11730 0 _106_
rlabel metal2 12926 11968 12926 11968 0 _107_
rlabel metal1 13248 11730 13248 11730 0 _108_
rlabel metal2 25438 3638 25438 3638 0 _109_
rlabel metal2 27278 3706 27278 3706 0 _110_
rlabel metal2 27278 6596 27278 6596 0 _111_
rlabel metal1 27232 8602 27232 8602 0 _112_
rlabel metal1 27232 10778 27232 10778 0 _113_
rlabel metal2 27278 13430 27278 13430 0 _114_
rlabel metal1 26864 16082 26864 16082 0 _115_
rlabel metal1 26910 18258 26910 18258 0 _116_
rlabel metal1 26910 20434 26910 20434 0 _117_
rlabel metal2 24150 21964 24150 21964 0 _118_
rlabel metal1 25944 21658 25944 21658 0 _119_
rlabel metal2 27278 21692 27278 21692 0 _120_
rlabel metal1 10534 12614 10534 12614 0 _121_
rlabel metal1 15686 17102 15686 17102 0 _122_
rlabel metal2 12466 15436 12466 15436 0 _123_
rlabel metal1 4738 17102 4738 17102 0 _124_
rlabel metal1 2484 3026 2484 3026 0 _125_
rlabel metal1 2484 8466 2484 8466 0 _126_
rlabel metal1 2346 12410 2346 12410 0 _127_
rlabel metal2 2254 17782 2254 17782 0 _128_
rlabel metal2 3910 20298 3910 20298 0 _129_
rlabel metal1 2806 20366 2806 20366 0 _130_
rlabel metal2 18814 3706 18814 3706 0 _131_
rlabel metal1 15034 13158 15034 13158 0 _132_
rlabel metal1 14398 13498 14398 13498 0 _133_
rlabel metal2 12466 13396 12466 13396 0 _134_
rlabel metal2 9706 12716 9706 12716 0 _135_
rlabel metal1 15456 17034 15456 17034 0 _136_
rlabel metal1 15318 13940 15318 13940 0 _137_
rlabel metal1 16376 13158 16376 13158 0 _138_
rlabel metal1 17066 9452 17066 9452 0 _139_
rlabel metal2 16974 10030 16974 10030 0 _140_
rlabel metal1 14030 12818 14030 12818 0 clk
rlabel metal1 20792 15130 20792 15130 0 clknet_0_clk
rlabel metal2 1748 7922 1748 7922 0 clknet_3_0__leaf_clk
rlabel metal2 16238 14144 16238 14144 0 clknet_3_1__leaf_clk
rlabel metal2 1794 21216 1794 21216 0 clknet_3_2__leaf_clk
rlabel metal2 17250 18292 17250 18292 0 clknet_3_3__leaf_clk
rlabel metal1 20378 3570 20378 3570 0 clknet_3_4__leaf_clk
rlabel metal1 22356 6834 22356 6834 0 clknet_3_5__leaf_clk
rlabel metal1 23046 22066 23046 22066 0 clknet_3_6__leaf_clk
rlabel metal1 25760 19890 25760 19890 0 clknet_3_7__leaf_clk
rlabel metal2 26174 1520 26174 1520 0 conversion_finished_out
rlabel metal1 12926 12274 12926 12274 0 dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal2 13386 11356 13386 11356 0 dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal2 12374 12478 12374 12478 0 dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel metal1 12926 13158 12926 13158 0 dac.parallel_cells\[0\].vdac_batch.vout_analog
rlabel metal1 6992 12206 6992 12206 0 dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal2 7590 11356 7590 11356 0 dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal1 7360 12274 7360 12274 0 dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal1 10994 10574 10994 10574 0 dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal1 12742 10030 12742 10030 0 dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel metal2 10442 10812 10442 10812 0 dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal1 4968 9486 4968 9486 0 dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal2 12742 8670 12742 8670 0 dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal2 4646 10880 4646 10880 0 dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal2 7314 8160 7314 8160 0 dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal1 9982 6834 9982 6834 0 dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal1 8280 6766 8280 6766 0 dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal1 8602 9486 8602 9486 0 dac.vdac_single.en_pupd
rlabel metal1 13662 13498 13662 13498 0 dcdc_trig_n_analog_w
rlabel metal1 12926 13906 12926 13906 0 dcdc_trigd_w
rlabel metal1 7774 4182 7774 4182 0 net1
rlabel metal1 28014 10982 28014 10982 0 net10
rlabel metal1 28060 13158 28060 13158 0 net11
rlabel metal2 28198 16116 28198 16116 0 net12
rlabel metal1 28152 17850 28152 17850 0 net13
rlabel metal1 27876 20570 27876 20570 0 net14
rlabel metal1 24196 22202 24196 22202 0 net15
rlabel metal2 1794 3196 1794 3196 0 net16
rlabel metal2 3450 7548 3450 7548 0 net17
rlabel metal1 2254 12206 2254 12206 0 net18
rlabel metal1 1656 17170 1656 17170 0 net19
rlabel metal1 18676 2618 18676 2618 0 net2
rlabel metal1 2484 22610 2484 22610 0 net20
rlabel metal1 2438 27438 2438 27438 0 net21
rlabel metal1 2629 17578 2629 17578 0 net22
rlabel metal1 13195 17238 13195 17238 0 net23
rlabel metal1 23375 3434 23375 3434 0 net24
rlabel metal2 23414 9996 23414 9996 0 net25
rlabel metal1 24978 21930 24978 21930 0 net26
rlabel metal1 17565 19414 17565 19414 0 net27
rlabel metal1 25537 17238 25537 17238 0 net28
rlabel metal1 4600 6222 4600 6222 0 net29
rlabel via1 26174 3349 26174 3349 0 net3
rlabel metal1 9292 9010 9292 9010 0 net30
rlabel metal2 26634 2890 26634 2890 0 net4
rlabel metal1 27370 22066 27370 22066 0 net5
rlabel metal1 27968 21114 27968 21114 0 net6
rlabel metal1 28106 4250 28106 4250 0 net7
rlabel metal1 27738 6188 27738 6188 0 net8
rlabel metal2 28290 8704 28290 8704 0 net9
rlabel metal1 11546 2414 11546 2414 0 rst_n
rlabel metal1 21114 18700 21114 18700 0 sar.compare_end_w
rlabel metal1 23276 4590 23276 4590 0 sar.counter_r\[0\]
rlabel metal2 19550 20128 19550 20128 0 sar.counter_r\[10\]
rlabel metal2 17526 18666 17526 18666 0 sar.counter_r\[11\]
rlabel metal1 22310 7276 22310 7276 0 sar.counter_r\[1\]
rlabel metal2 24150 6154 24150 6154 0 sar.counter_r\[2\]
rlabel metal2 23322 8636 23322 8636 0 sar.counter_r\[3\]
rlabel metal1 21988 12614 21988 12614 0 sar.counter_r\[4\]
rlabel metal2 22310 12546 22310 12546 0 sar.counter_r\[5\]
rlabel metal2 24242 14518 24242 14518 0 sar.counter_r\[6\]
rlabel metal1 24196 16422 24196 16422 0 sar.counter_r\[7\]
rlabel metal2 21298 19618 21298 19618 0 sar.counter_r\[9\]
rlabel metal2 11270 13124 11270 13124 0 sar.current_dac_bit_r\[0\]
rlabel metal2 10626 15776 10626 15776 0 sar.current_dac_bit_r\[1\]
rlabel metal1 8188 14926 8188 14926 0 sar.current_dac_bit_r\[2\]
rlabel metal1 8142 16014 8142 16014 0 sar.current_dac_bit_r\[3\]
rlabel via1 8510 17578 8510 17578 0 sar.current_dac_bit_r\[4\]
rlabel metal1 12995 16966 12995 16966 0 sar.current_dac_bit_r\[5\]
rlabel via1 10994 13498 10994 13498 0 sar.dac_value_r\[0\]
rlabel metal1 2760 11526 2760 11526 0 sar.dac_value_r\[1\]
rlabel metal1 3772 14790 3772 14790 0 sar.dac_value_r\[2\]
rlabel metal1 2208 15674 2208 15674 0 sar.dac_value_r\[3\]
rlabel metal1 5520 20842 5520 20842 0 sar.dac_value_r\[4\]
rlabel metal1 3082 18394 3082 18394 0 sar.dac_value_r\[5\]
rlabel metal1 14030 13362 14030 13362 0 sar.dcdc_dat_out
rlabel metal1 18906 6970 18906 6970 0 sar.next_counter_w\[0\]
rlabel metal1 18216 18938 18216 18938 0 sar.next_counter_w\[10\]
rlabel metal1 15686 16626 15686 16626 0 sar.next_counter_w\[11\]
rlabel metal1 19412 5814 19412 5814 0 sar.next_counter_w\[1\]
rlabel metal1 22540 6426 22540 6426 0 sar.next_counter_w\[2\]
rlabel metal2 21850 8738 21850 8738 0 sar.next_counter_w\[3\]
rlabel metal2 20378 10268 20378 10268 0 sar.next_counter_w\[4\]
rlabel metal1 20608 11866 20608 11866 0 sar.next_counter_w\[5\]
rlabel metal1 22770 14008 22770 14008 0 sar.next_counter_w\[6\]
rlabel metal2 22126 16354 22126 16354 0 sar.next_counter_w\[7\]
rlabel metal2 18446 14382 18446 14382 0 sar.next_counter_w\[8\]
rlabel metal2 20654 17612 20654 17612 0 sar.next_counter_w\[9\]
rlabel metal1 24610 3978 24610 3978 0 sar.next_ticks_w\[0\]
rlabel metal2 19458 21726 19458 21726 0 sar.next_ticks_w\[10\]
rlabel metal2 18262 21080 18262 21080 0 sar.next_ticks_w\[11\]
rlabel metal1 22218 4012 22218 4012 0 sar.next_ticks_w\[1\]
rlabel metal1 26956 6358 26956 6358 0 sar.next_ticks_w\[2\]
rlabel metal2 25990 9180 25990 9180 0 sar.next_ticks_w\[3\]
rlabel metal1 23782 11526 23782 11526 0 sar.next_ticks_w\[4\]
rlabel metal2 25898 13022 25898 13022 0 sar.next_ticks_w\[5\]
rlabel metal2 25990 15810 25990 15810 0 sar.next_ticks_w\[6\]
rlabel metal1 24794 17850 24794 17850 0 sar.next_ticks_w\[7\]
rlabel metal1 24242 19278 24242 19278 0 sar.next_ticks_w\[8\]
rlabel metal1 23460 21590 23460 21590 0 sar.next_ticks_w\[9\]
rlabel metal2 16974 12886 16974 12886 0 sar.state_r\[0\]
rlabel metal1 16928 13362 16928 13362 0 sar.state_r\[1\]
rlabel metal2 17066 13022 17066 13022 0 sar.state_r\[2\]
rlabel metal1 23828 3162 23828 3162 0 sar.ticks_r\[0\]
rlabel metal2 20470 21148 20470 21148 0 sar.ticks_r\[10\]
rlabel metal1 17066 19890 17066 19890 0 sar.ticks_r\[11\]
rlabel metal1 23092 3706 23092 3706 0 sar.ticks_r\[1\]
rlabel metal2 25254 5916 25254 5916 0 sar.ticks_r\[2\]
rlabel metal1 24656 8602 24656 8602 0 sar.ticks_r\[3\]
rlabel metal2 23506 10982 23506 10982 0 sar.ticks_r\[4\]
rlabel metal1 24932 12274 24932 12274 0 sar.ticks_r\[5\]
rlabel metal1 24978 15130 24978 15130 0 sar.ticks_r\[6\]
rlabel metal1 25116 16966 25116 16966 0 sar.ticks_r\[7\]
rlabel metal2 24978 18972 24978 18972 0 sar.ticks_r\[8\]
rlabel metal2 22402 20944 22402 20944 0 sar.ticks_r\[9\]
rlabel metal2 12558 13294 12558 13294 0 sar.time_trigd_n_in
rlabel metal1 18860 2414 18860 2414 0 start_conv_in
rlabel metal2 28382 1853 28382 1853 0 tick_result_out[0]
rlabel metal3 28850 25908 28850 25908 0 tick_result_out[10]
rlabel metal2 28382 27965 28382 27965 0 tick_result_out[11]
rlabel metal2 28382 3791 28382 3791 0 tick_result_out[1]
rlabel metal2 28382 6477 28382 6477 0 tick_result_out[2]
rlabel metal2 28382 9061 28382 9061 0 tick_result_out[3]
rlabel metal2 28382 11373 28382 11373 0 tick_result_out[4]
rlabel via2 28382 13685 28382 13685 0 tick_result_out[5]
rlabel metal2 28382 16269 28382 16269 0 tick_result_out[6]
rlabel via2 28382 18581 28382 18581 0 tick_result_out[7]
rlabel metal2 28382 21165 28382 21165 0 tick_result_out[8]
rlabel via2 28382 23477 28382 23477 0 tick_result_out[9]
rlabel metal3 1142 2652 1142 2652 0 vdac_result_out[0]
rlabel via2 1610 7531 1610 7531 0 vdac_result_out[1]
rlabel metal1 1564 12410 1564 12410 0 vdac_result_out[2]
rlabel via2 1610 17323 1610 17323 0 vdac_result_out[3]
rlabel metal3 1142 22236 1142 22236 0 vdac_result_out[4]
rlabel metal3 1142 27132 1142 27132 0 vdac_result_out[5]
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
