magic
tech sky130A
magscale 1 2
timestamp 1672094039
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 14 2128 59970 57712
<< metal2 >>
rect 1306 59200 1362 60000
rect 3238 59200 3294 60000
rect 5170 59200 5226 60000
rect 7102 59200 7158 60000
rect 8390 59200 8446 60000
rect 10322 59200 10378 60000
rect 12254 59200 12310 60000
rect 14186 59200 14242 60000
rect 16118 59200 16174 60000
rect 18050 59200 18106 60000
rect 19982 59200 20038 60000
rect 21270 59200 21326 60000
rect 23202 59200 23258 60000
rect 25134 59200 25190 60000
rect 27066 59200 27122 60000
rect 28998 59200 29054 60000
rect 30930 59200 30986 60000
rect 32862 59200 32918 60000
rect 34150 59200 34206 60000
rect 36082 59200 36138 60000
rect 38014 59200 38070 60000
rect 39946 59200 40002 60000
rect 41878 59200 41934 60000
rect 43810 59200 43866 60000
rect 45742 59200 45798 60000
rect 47030 59200 47086 60000
rect 48962 59200 49018 60000
rect 50894 59200 50950 60000
rect 52826 59200 52882 60000
rect 54758 59200 54814 60000
rect 56690 59200 56746 60000
rect 58622 59200 58678 60000
rect 59910 59200 59966 60000
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 7102 0 7158 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 16118 0 16174 800
rect 18050 0 18106 800
rect 19982 0 20038 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28998 0 29054 800
rect 30930 0 30986 800
rect 32862 0 32918 800
rect 34794 0 34850 800
rect 36726 0 36782 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 49606 0 49662 800
rect 51538 0 51594 800
rect 52826 0 52882 800
rect 54758 0 54814 800
rect 56690 0 56746 800
rect 58622 0 58678 800
<< obsm2 >>
rect 20 59144 1250 59945
rect 1418 59144 3182 59945
rect 3350 59144 5114 59945
rect 5282 59144 7046 59945
rect 7214 59144 8334 59945
rect 8502 59144 10266 59945
rect 10434 59144 12198 59945
rect 12366 59144 14130 59945
rect 14298 59144 16062 59945
rect 16230 59144 17994 59945
rect 18162 59144 19926 59945
rect 20094 59144 21214 59945
rect 21382 59144 23146 59945
rect 23314 59144 25078 59945
rect 25246 59144 27010 59945
rect 27178 59144 28942 59945
rect 29110 59144 30874 59945
rect 31042 59144 32806 59945
rect 32974 59144 34094 59945
rect 34262 59144 36026 59945
rect 36194 59144 37958 59945
rect 38126 59144 39890 59945
rect 40058 59144 41822 59945
rect 41990 59144 43754 59945
rect 43922 59144 45686 59945
rect 45854 59144 46974 59945
rect 47142 59144 48906 59945
rect 49074 59144 50838 59945
rect 51006 59144 52770 59945
rect 52938 59144 54702 59945
rect 54870 59144 56634 59945
rect 56802 59144 58566 59945
rect 58734 59144 59854 59945
rect 20 856 59964 59144
rect 130 31 1250 856
rect 1418 31 3182 856
rect 3350 31 5114 856
rect 5282 31 7046 856
rect 7214 31 8978 856
rect 9146 31 10910 856
rect 11078 31 12842 856
rect 13010 31 14130 856
rect 14298 31 16062 856
rect 16230 31 17994 856
rect 18162 31 19926 856
rect 20094 31 21858 856
rect 22026 31 23790 856
rect 23958 31 25722 856
rect 25890 31 27010 856
rect 27178 31 28942 856
rect 29110 31 30874 856
rect 31042 31 32806 856
rect 32974 31 34738 856
rect 34906 31 36670 856
rect 36838 31 38602 856
rect 38770 31 39890 856
rect 40058 31 41822 856
rect 41990 31 43754 856
rect 43922 31 45686 856
rect 45854 31 47618 856
rect 47786 31 49550 856
rect 49718 31 51482 856
rect 51650 31 52770 856
rect 52938 31 54702 856
rect 54870 31 56634 856
rect 56802 31 58566 856
rect 58734 31 59964 856
<< metal3 >>
rect 0 59848 800 59968
rect 59200 58488 60000 58608
rect 0 57808 800 57928
rect 59200 56448 60000 56568
rect 0 55768 800 55888
rect 0 54408 800 54528
rect 59200 54408 60000 54528
rect 0 52368 800 52488
rect 59200 52368 60000 52488
rect 0 50328 800 50448
rect 59200 50328 60000 50448
rect 0 48288 800 48408
rect 59200 48288 60000 48408
rect 0 46248 800 46368
rect 59200 46248 60000 46368
rect 59200 44888 60000 45008
rect 0 44208 800 44328
rect 59200 42848 60000 42968
rect 0 42168 800 42288
rect 0 40808 800 40928
rect 59200 40808 60000 40928
rect 0 38768 800 38888
rect 59200 38768 60000 38888
rect 0 36728 800 36848
rect 59200 36728 60000 36848
rect 0 34688 800 34808
rect 59200 34688 60000 34808
rect 0 32648 800 32768
rect 59200 32648 60000 32768
rect 59200 31288 60000 31408
rect 0 30608 800 30728
rect 59200 29248 60000 29368
rect 0 28568 800 28688
rect 0 27208 800 27328
rect 59200 27208 60000 27328
rect 0 25168 800 25288
rect 59200 25168 60000 25288
rect 0 23128 800 23248
rect 59200 23128 60000 23248
rect 0 21088 800 21208
rect 59200 21088 60000 21208
rect 0 19048 800 19168
rect 59200 19048 60000 19168
rect 59200 17688 60000 17808
rect 0 17008 800 17128
rect 59200 15648 60000 15768
rect 0 14968 800 15088
rect 0 13608 800 13728
rect 59200 13608 60000 13728
rect 0 11568 800 11688
rect 59200 11568 60000 11688
rect 0 9528 800 9648
rect 59200 9528 60000 9648
rect 0 7488 800 7608
rect 59200 7488 60000 7608
rect 0 5448 800 5568
rect 59200 5448 60000 5568
rect 59200 4088 60000 4208
rect 0 3408 800 3528
rect 59200 2048 60000 2168
rect 0 1368 800 1488
rect 59200 8 60000 128
<< obsm3 >>
rect 880 59768 59200 59941
rect 800 58688 59200 59768
rect 800 58408 59120 58688
rect 800 58008 59200 58408
rect 880 57728 59200 58008
rect 800 56648 59200 57728
rect 800 56368 59120 56648
rect 800 55968 59200 56368
rect 880 55688 59200 55968
rect 800 54608 59200 55688
rect 880 54328 59120 54608
rect 800 52568 59200 54328
rect 880 52288 59120 52568
rect 800 50528 59200 52288
rect 880 50248 59120 50528
rect 800 48488 59200 50248
rect 880 48208 59120 48488
rect 800 46448 59200 48208
rect 880 46168 59120 46448
rect 800 45088 59200 46168
rect 800 44808 59120 45088
rect 800 44408 59200 44808
rect 880 44128 59200 44408
rect 800 43048 59200 44128
rect 800 42768 59120 43048
rect 800 42368 59200 42768
rect 880 42088 59200 42368
rect 800 41008 59200 42088
rect 880 40728 59120 41008
rect 800 38968 59200 40728
rect 880 38688 59120 38968
rect 800 36928 59200 38688
rect 880 36648 59120 36928
rect 800 34888 59200 36648
rect 880 34608 59120 34888
rect 800 32848 59200 34608
rect 880 32568 59120 32848
rect 800 31488 59200 32568
rect 800 31208 59120 31488
rect 800 30808 59200 31208
rect 880 30528 59200 30808
rect 800 29448 59200 30528
rect 800 29168 59120 29448
rect 800 28768 59200 29168
rect 880 28488 59200 28768
rect 800 27408 59200 28488
rect 880 27128 59120 27408
rect 800 25368 59200 27128
rect 880 25088 59120 25368
rect 800 23328 59200 25088
rect 880 23048 59120 23328
rect 800 21288 59200 23048
rect 880 21008 59120 21288
rect 800 19248 59200 21008
rect 880 18968 59120 19248
rect 800 17888 59200 18968
rect 800 17608 59120 17888
rect 800 17208 59200 17608
rect 880 16928 59200 17208
rect 800 15848 59200 16928
rect 800 15568 59120 15848
rect 800 15168 59200 15568
rect 880 14888 59200 15168
rect 800 13808 59200 14888
rect 880 13528 59120 13808
rect 800 11768 59200 13528
rect 880 11488 59120 11768
rect 800 9728 59200 11488
rect 880 9448 59120 9728
rect 800 7688 59200 9448
rect 880 7408 59120 7688
rect 800 5648 59200 7408
rect 880 5368 59120 5648
rect 800 4288 59200 5368
rect 800 4008 59120 4288
rect 800 3608 59200 4008
rect 880 3328 59200 3608
rect 800 2248 59200 3328
rect 800 1968 59120 2248
rect 800 1568 59200 1968
rect 880 1288 59200 1568
rect 800 208 59200 1288
rect 800 35 59120 208
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< labels >>
rlabel metal3 s 59200 58488 60000 58608 6 tie_hi[0]
port 1 nsew signal output
rlabel metal3 s 59200 21088 60000 21208 6 tie_hi[10]
port 2 nsew signal output
rlabel metal3 s 59200 32648 60000 32768 6 tie_hi[11]
port 3 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 tie_hi[12]
port 4 nsew signal output
rlabel metal2 s 27066 59200 27122 60000 6 tie_hi[13]
port 5 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 tie_hi[14]
port 6 nsew signal output
rlabel metal2 s 28998 59200 29054 60000 6 tie_hi[15]
port 7 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 tie_hi[16]
port 8 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 tie_hi[17]
port 9 nsew signal output
rlabel metal2 s 50894 59200 50950 60000 6 tie_hi[18]
port 10 nsew signal output
rlabel metal2 s 10322 59200 10378 60000 6 tie_hi[19]
port 11 nsew signal output
rlabel metal2 s 52826 59200 52882 60000 6 tie_hi[1]
port 12 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 tie_hi[20]
port 13 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 tie_hi[21]
port 14 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 tie_hi[22]
port 15 nsew signal output
rlabel metal3 s 59200 19048 60000 19168 6 tie_hi[23]
port 16 nsew signal output
rlabel metal2 s 59910 59200 59966 60000 6 tie_hi[24]
port 17 nsew signal output
rlabel metal3 s 59200 13608 60000 13728 6 tie_hi[25]
port 18 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 tie_hi[26]
port 19 nsew signal output
rlabel metal2 s 25134 59200 25190 60000 6 tie_hi[27]
port 20 nsew signal output
rlabel metal3 s 59200 44888 60000 45008 6 tie_hi[28]
port 21 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 tie_hi[29]
port 22 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 tie_hi[2]
port 23 nsew signal output
rlabel metal2 s 14186 59200 14242 60000 6 tie_hi[30]
port 24 nsew signal output
rlabel metal3 s 59200 34688 60000 34808 6 tie_hi[31]
port 25 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 tie_hi[3]
port 26 nsew signal output
rlabel metal2 s 56690 59200 56746 60000 6 tie_hi[4]
port 27 nsew signal output
rlabel metal2 s 32862 59200 32918 60000 6 tie_hi[5]
port 28 nsew signal output
rlabel metal3 s 59200 40808 60000 40928 6 tie_hi[6]
port 29 nsew signal output
rlabel metal2 s 38014 59200 38070 60000 6 tie_hi[7]
port 30 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 tie_hi[8]
port 31 nsew signal output
rlabel metal3 s 59200 29248 60000 29368 6 tie_hi[9]
port 32 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 tie_lo[0]
port 33 nsew signal output
rlabel metal3 s 59200 42848 60000 42968 6 tie_lo[10]
port 34 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 tie_lo[11]
port 35 nsew signal output
rlabel metal2 s 58622 59200 58678 60000 6 tie_lo[12]
port 36 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 tie_lo[13]
port 37 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 tie_lo[14]
port 38 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 tie_lo[15]
port 39 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 tie_lo[16]
port 40 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 tie_lo[17]
port 41 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 tie_lo[18]
port 42 nsew signal output
rlabel metal2 s 34150 59200 34206 60000 6 tie_lo[19]
port 43 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 tie_lo[1]
port 44 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 tie_lo[20]
port 45 nsew signal output
rlabel metal2 s 7102 59200 7158 60000 6 tie_lo[21]
port 46 nsew signal output
rlabel metal2 s 41878 59200 41934 60000 6 tie_lo[22]
port 47 nsew signal output
rlabel metal2 s 18050 59200 18106 60000 6 tie_lo[23]
port 48 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 tie_lo[24]
port 49 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 tie_lo[25]
port 50 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 tie_lo[26]
port 51 nsew signal output
rlabel metal3 s 59200 4088 60000 4208 6 tie_lo[27]
port 52 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 tie_lo[28]
port 53 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 tie_lo[29]
port 54 nsew signal output
rlabel metal3 s 59200 56448 60000 56568 6 tie_lo[2]
port 55 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 tie_lo[30]
port 56 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 tie_lo[31]
port 57 nsew signal output
rlabel metal2 s 16118 59200 16174 60000 6 tie_lo[32]
port 58 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 tie_lo[33]
port 59 nsew signal output
rlabel metal3 s 59200 52368 60000 52488 6 tie_lo[34]
port 60 nsew signal output
rlabel metal3 s 59200 46248 60000 46368 6 tie_lo[35]
port 61 nsew signal output
rlabel metal2 s 5170 59200 5226 60000 6 tie_lo[36]
port 62 nsew signal output
rlabel metal2 s 8390 59200 8446 60000 6 tie_lo[37]
port 63 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 tie_lo[38]
port 64 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 tie_lo[39]
port 65 nsew signal output
rlabel metal2 s 21270 59200 21326 60000 6 tie_lo[3]
port 66 nsew signal output
rlabel metal3 s 59200 23128 60000 23248 6 tie_lo[40]
port 67 nsew signal output
rlabel metal3 s 59200 15648 60000 15768 6 tie_lo[41]
port 68 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 tie_lo[42]
port 69 nsew signal output
rlabel metal2 s 23202 59200 23258 60000 6 tie_lo[43]
port 70 nsew signal output
rlabel metal3 s 59200 8 60000 128 6 tie_lo[44]
port 71 nsew signal output
rlabel metal3 s 59200 17688 60000 17808 6 tie_lo[45]
port 72 nsew signal output
rlabel metal2 s 47030 59200 47086 60000 6 tie_lo[46]
port 73 nsew signal output
rlabel metal3 s 59200 9528 60000 9648 6 tie_lo[47]
port 74 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 tie_lo[48]
port 75 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 tie_lo[49]
port 76 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 tie_lo[4]
port 77 nsew signal output
rlabel metal3 s 59200 54408 60000 54528 6 tie_lo[50]
port 78 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 tie_lo[51]
port 79 nsew signal output
rlabel metal3 s 59200 5448 60000 5568 6 tie_lo[52]
port 80 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 tie_lo[53]
port 81 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 tie_lo[54]
port 82 nsew signal output
rlabel metal2 s 30930 59200 30986 60000 6 tie_lo[55]
port 83 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 tie_lo[56]
port 84 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 tie_lo[57]
port 85 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 tie_lo[58]
port 86 nsew signal output
rlabel metal3 s 59200 2048 60000 2168 6 tie_lo[59]
port 87 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 tie_lo[5]
port 88 nsew signal output
rlabel metal3 s 59200 25168 60000 25288 6 tie_lo[60]
port 89 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 tie_lo[61]
port 90 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 tie_lo[62]
port 91 nsew signal output
rlabel metal3 s 59200 11568 60000 11688 6 tie_lo[63]
port 92 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 tie_lo[64]
port 93 nsew signal output
rlabel metal3 s 59200 31288 60000 31408 6 tie_lo[65]
port 94 nsew signal output
rlabel metal3 s 59200 48288 60000 48408 6 tie_lo[66]
port 95 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 tie_lo[67]
port 96 nsew signal output
rlabel metal3 s 59200 50328 60000 50448 6 tie_lo[68]
port 97 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 tie_lo[69]
port 98 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 tie_lo[6]
port 99 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 tie_lo[70]
port 100 nsew signal output
rlabel metal2 s 18 0 74 800 6 tie_lo[71]
port 101 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 tie_lo[72]
port 102 nsew signal output
rlabel metal2 s 1306 59200 1362 60000 6 tie_lo[73]
port 103 nsew signal output
rlabel metal2 s 19982 59200 20038 60000 6 tie_lo[74]
port 104 nsew signal output
rlabel metal2 s 39946 59200 40002 60000 6 tie_lo[75]
port 105 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 tie_lo[76]
port 106 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 tie_lo[77]
port 107 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 tie_lo[78]
port 108 nsew signal output
rlabel metal2 s 48962 59200 49018 60000 6 tie_lo[79]
port 109 nsew signal output
rlabel metal2 s 36082 59200 36138 60000 6 tie_lo[7]
port 110 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 tie_lo[80]
port 111 nsew signal output
rlabel metal2 s 54758 59200 54814 60000 6 tie_lo[81]
port 112 nsew signal output
rlabel metal3 s 59200 7488 60000 7608 6 tie_lo[82]
port 113 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 tie_lo[83]
port 114 nsew signal output
rlabel metal3 s 59200 36728 60000 36848 6 tie_lo[84]
port 115 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 tie_lo[85]
port 116 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 tie_lo[86]
port 117 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 tie_lo[87]
port 118 nsew signal output
rlabel metal3 s 59200 38768 60000 38888 6 tie_lo[88]
port 119 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 tie_lo[89]
port 120 nsew signal output
rlabel metal2 s 45742 59200 45798 60000 6 tie_lo[8]
port 121 nsew signal output
rlabel metal2 s 43810 59200 43866 60000 6 tie_lo[90]
port 122 nsew signal output
rlabel metal2 s 3238 59200 3294 60000 6 tie_lo[91]
port 123 nsew signal output
rlabel metal2 s 12254 59200 12310 60000 6 tie_lo[92]
port 124 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 tie_lo[93]
port 125 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 tie_lo[94]
port 126 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 tie_lo[95]
port 127 nsew signal output
rlabel metal3 s 59200 27208 60000 27328 6 tie_lo[9]
port 128 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 129 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 130 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 130 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1014404
string GDS_FILE /foss/designs/openlane/const_gen/runs/foo/results/signoff/const_gen.magic.gds
string GDS_START 23752
<< end >>

