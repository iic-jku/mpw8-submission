magic
tech sky130A
magscale 1 2
timestamp 1672093988
<< viali >>
rect 4537 57545 4571 57579
rect 17693 57545 17727 57579
rect 25421 57545 25455 57579
rect 26617 57545 26651 57579
rect 29193 57545 29227 57579
rect 34253 57545 34287 57579
rect 47777 57545 47811 57579
rect 50353 57545 50387 57579
rect 11161 57477 11195 57511
rect 13737 57477 13771 57511
rect 16221 57477 16255 57511
rect 1961 57409 1995 57443
rect 2237 57409 2271 57443
rect 3249 57409 3283 57443
rect 4353 57409 4387 57443
rect 6009 57409 6043 57443
rect 6745 57409 6779 57443
rect 8585 57409 8619 57443
rect 9137 57409 9171 57443
rect 9873 57409 9907 57443
rect 10333 57409 10367 57443
rect 11713 57409 11747 57443
rect 12725 57409 12759 57443
rect 14289 57409 14323 57443
rect 15117 57409 15151 57443
rect 16865 57409 16899 57443
rect 17509 57409 17543 57443
rect 18245 57409 18279 57443
rect 18705 57409 18739 57443
rect 19901 57409 19935 57443
rect 20637 57409 20671 57443
rect 21097 57409 21131 57443
rect 22293 57409 22327 57443
rect 23029 57409 23063 57443
rect 23489 57409 23523 57443
rect 24685 57409 24719 57443
rect 26065 57409 26099 57443
rect 27353 57409 27387 57443
rect 28273 57409 28307 57443
rect 29929 57409 29963 57443
rect 30665 57409 30699 57443
rect 31309 57409 31343 57443
rect 32321 57409 32355 57443
rect 33057 57409 33091 57443
rect 33701 57409 33735 57443
rect 34897 57409 34931 57443
rect 35725 57409 35759 57443
rect 36829 57409 36863 57443
rect 38025 57409 38059 57443
rect 38485 57409 38519 57443
rect 39221 57409 39255 57443
rect 40417 57409 40451 57443
rect 40877 57409 40911 57443
rect 41613 57409 41647 57443
rect 42809 57409 42843 57443
rect 43269 57409 43303 57443
rect 44005 57409 44039 57443
rect 44465 57409 44499 57443
rect 45385 57409 45419 57443
rect 46397 57409 46431 57443
rect 46857 57409 46891 57443
rect 47961 57409 47995 57443
rect 48789 57409 48823 57443
rect 49249 57409 49283 57443
rect 50537 57409 50571 57443
rect 51181 57409 51215 57443
rect 51641 57409 51675 57443
rect 52377 57409 52411 57443
rect 53573 57409 53607 57443
rect 54033 57409 54067 57443
rect 54769 57409 54803 57443
rect 55965 57409 55999 57443
rect 56425 57409 56459 57443
rect 57161 57409 57195 57443
rect 58357 57409 58391 57443
rect 5733 57341 5767 57375
rect 8309 57341 8343 57375
rect 10517 57273 10551 57307
rect 14473 57273 14507 57307
rect 15301 57273 15335 57307
rect 21281 57273 21315 57307
rect 23673 57273 23707 57307
rect 30849 57273 30883 57307
rect 40233 57273 40267 57307
rect 42625 57273 42659 57307
rect 43821 57273 43855 57307
rect 48605 57273 48639 57307
rect 50997 57273 51031 57307
rect 56977 57273 57011 57307
rect 3433 57205 3467 57239
rect 6929 57205 6963 57239
rect 9321 57205 9355 57239
rect 11897 57205 11931 57239
rect 12909 57205 12943 57239
rect 17049 57205 17083 57239
rect 18889 57205 18923 57239
rect 20085 57205 20119 57239
rect 22477 57205 22511 57239
rect 24869 57205 24903 57239
rect 25881 57205 25915 57239
rect 27169 57205 27203 57239
rect 28457 57205 28491 57239
rect 29745 57205 29779 57239
rect 32505 57205 32539 57239
rect 33241 57205 33275 57239
rect 35081 57205 35115 57239
rect 35541 57205 35575 57239
rect 36645 57205 36679 57239
rect 37841 57205 37875 57239
rect 39037 57205 39071 57239
rect 41429 57205 41463 57239
rect 45201 57205 45235 57239
rect 46213 57205 46247 57239
rect 52193 57205 52227 57239
rect 53389 57205 53423 57239
rect 54585 57205 54619 57239
rect 55781 57205 55815 57239
rect 58173 57205 58207 57239
rect 1869 57001 1903 57035
rect 3065 57001 3099 57035
rect 4261 57001 4295 57035
rect 6009 57001 6043 57035
rect 6653 57001 6687 57035
rect 8493 57001 8527 57035
rect 9137 57001 9171 57035
rect 12633 57001 12667 57035
rect 15025 57001 15059 57035
rect 19809 57001 19843 57035
rect 21649 57001 21683 57035
rect 22201 57001 22235 57035
rect 24593 57001 24627 57035
rect 25881 57001 25915 57035
rect 28181 57001 28215 57035
rect 32137 57001 32171 57035
rect 35357 57001 35391 57035
rect 36461 57001 36495 57035
rect 38301 57001 38335 57035
rect 41337 57001 41371 57035
rect 45201 57001 45235 57035
rect 47593 57001 47627 57035
rect 50353 57001 50387 57035
rect 52101 57001 52135 57035
rect 54493 57001 54527 57035
rect 56425 57001 56459 57035
rect 29745 56865 29779 56899
rect 21465 56797 21499 56831
rect 29837 56797 29871 56831
rect 30021 56797 30055 56831
rect 38945 56797 38979 56831
rect 39037 56797 39071 56831
rect 39221 56797 39255 56831
rect 39313 56797 39347 56831
rect 43591 56797 43625 56831
rect 44004 56797 44038 56831
rect 44097 56797 44131 56831
rect 57069 56797 57103 56831
rect 57529 56797 57563 56831
rect 58357 56797 58391 56831
rect 17417 56729 17451 56763
rect 21281 56729 21315 56763
rect 43729 56729 43763 56763
rect 43821 56729 43855 56763
rect 55873 56729 55907 56763
rect 30205 56661 30239 56695
rect 38761 56661 38795 56695
rect 43453 56661 43487 56695
rect 56885 56661 56919 56695
rect 57713 56661 57747 56695
rect 58173 56661 58207 56695
rect 30573 56457 30607 56491
rect 35173 56457 35207 56491
rect 38301 56457 38335 56491
rect 57161 56457 57195 56491
rect 21281 56389 21315 56423
rect 23581 56389 23615 56423
rect 23673 56389 23707 56423
rect 26249 56389 26283 56423
rect 28549 56389 28583 56423
rect 30205 56389 30239 56423
rect 30317 56389 30351 56423
rect 33057 56389 33091 56423
rect 35449 56389 35483 56423
rect 36553 56389 36587 56423
rect 41521 56389 41555 56423
rect 56701 56389 56735 56423
rect 21097 56321 21131 56355
rect 22017 56321 22051 56355
rect 22201 56321 22235 56355
rect 23484 56321 23518 56355
rect 23856 56321 23890 56355
rect 23949 56321 23983 56355
rect 25053 56321 25087 56355
rect 25329 56321 25363 56355
rect 25973 56321 26007 56355
rect 26157 56321 26191 56355
rect 26393 56321 26427 56355
rect 28273 56321 28307 56355
rect 28366 56321 28400 56355
rect 28641 56321 28675 56355
rect 28779 56321 28813 56355
rect 29929 56321 29963 56355
rect 30022 56321 30056 56355
rect 30394 56321 30428 56355
rect 31033 56321 31067 56355
rect 31217 56321 31251 56355
rect 31309 56321 31343 56355
rect 31453 56321 31487 56355
rect 32960 56321 32994 56355
rect 33149 56321 33183 56355
rect 33332 56321 33366 56355
rect 33425 56321 33459 56355
rect 35352 56321 35386 56355
rect 35541 56321 35575 56355
rect 35724 56321 35758 56355
rect 35817 56321 35851 56355
rect 36456 56321 36490 56355
rect 36645 56321 36679 56355
rect 36828 56321 36862 56355
rect 36921 56321 36955 56355
rect 38485 56321 38519 56355
rect 38577 56321 38611 56355
rect 38761 56321 38795 56355
rect 38853 56321 38887 56355
rect 39313 56321 39347 56355
rect 39405 56321 39439 56355
rect 39589 56321 39623 56355
rect 39681 56321 39715 56355
rect 41424 56321 41458 56355
rect 41613 56321 41647 56355
rect 41796 56321 41830 56355
rect 41889 56321 41923 56355
rect 43448 56321 43482 56355
rect 43545 56321 43579 56355
rect 43637 56321 43671 56355
rect 43820 56321 43854 56355
rect 43913 56321 43947 56355
rect 56149 56321 56183 56355
rect 58357 56321 58391 56355
rect 21465 56185 21499 56219
rect 31585 56185 31619 56219
rect 36277 56185 36311 56219
rect 43269 56185 43303 56219
rect 22385 56117 22419 56151
rect 23305 56117 23339 56151
rect 25145 56117 25179 56151
rect 25513 56117 25547 56151
rect 26525 56117 26559 56151
rect 28917 56117 28951 56151
rect 32781 56117 32815 56151
rect 39865 56117 39899 56151
rect 41245 56117 41279 56151
rect 58173 56117 58207 56151
rect 24593 55913 24627 55947
rect 26249 55913 26283 55947
rect 28089 55913 28123 55947
rect 28457 55913 28491 55947
rect 38485 55913 38519 55947
rect 57161 55913 57195 55947
rect 23673 55845 23707 55879
rect 30297 55845 30331 55879
rect 25053 55777 25087 55811
rect 28549 55777 28583 55811
rect 36277 55777 36311 55811
rect 1869 55709 1903 55743
rect 2329 55709 2363 55743
rect 23121 55709 23155 55743
rect 23305 55709 23339 55743
rect 23541 55709 23575 55743
rect 24777 55709 24811 55743
rect 24961 55709 24995 55743
rect 25605 55709 25639 55743
rect 25753 55709 25787 55743
rect 25881 55709 25915 55743
rect 26070 55709 26104 55743
rect 28273 55709 28307 55743
rect 29745 55709 29779 55743
rect 29929 55709 29963 55743
rect 30165 55709 30199 55743
rect 33011 55709 33045 55743
rect 33149 55709 33183 55743
rect 33241 55709 33275 55743
rect 33424 55709 33458 55743
rect 33517 55709 33551 55743
rect 35076 55709 35110 55743
rect 35448 55709 35482 55743
rect 35541 55709 35575 55743
rect 36461 55709 36495 55743
rect 36553 55709 36587 55743
rect 36737 55709 36771 55743
rect 36829 55709 36863 55743
rect 38669 55709 38703 55743
rect 38761 55709 38795 55743
rect 38930 55709 38964 55743
rect 39037 55703 39071 55737
rect 41659 55709 41693 55743
rect 42072 55709 42106 55743
rect 42165 55709 42199 55743
rect 43407 55709 43441 55743
rect 43637 55709 43671 55743
rect 43820 55709 43854 55743
rect 43913 55709 43947 55743
rect 57713 55709 57747 55743
rect 58357 55709 58391 55743
rect 21281 55641 21315 55675
rect 21465 55641 21499 55675
rect 21649 55641 21683 55675
rect 22661 55641 22695 55675
rect 23397 55641 23431 55675
rect 25973 55641 26007 55675
rect 30021 55641 30055 55675
rect 35173 55641 35207 55675
rect 35265 55641 35299 55675
rect 41797 55641 41831 55675
rect 41889 55641 41923 55675
rect 43545 55641 43579 55675
rect 1685 55573 1719 55607
rect 29101 55573 29135 55607
rect 30849 55573 30883 55607
rect 32873 55573 32907 55607
rect 34897 55573 34931 55607
rect 37933 55573 37967 55607
rect 41521 55573 41555 55607
rect 43269 55573 43303 55607
rect 58173 55573 58207 55607
rect 32505 55369 32539 55403
rect 41429 55369 41463 55403
rect 43361 55369 43395 55403
rect 58173 55369 58207 55403
rect 43637 55301 43671 55335
rect 1869 55233 1903 55267
rect 2421 55233 2455 55267
rect 31769 55233 31803 55267
rect 32689 55233 32723 55267
rect 39865 55233 39899 55267
rect 43499 55233 43533 55267
rect 43729 55233 43763 55267
rect 43912 55233 43946 55267
rect 44005 55233 44039 55267
rect 57529 55233 57563 55267
rect 58357 55233 58391 55267
rect 32321 55165 32355 55199
rect 1685 55029 1719 55063
rect 32689 55029 32723 55063
rect 40325 55029 40359 55063
rect 40877 55029 40911 55063
rect 24961 54825 24995 54859
rect 40509 54825 40543 54859
rect 41337 54825 41371 54859
rect 41521 54825 41555 54859
rect 40693 54757 40727 54791
rect 25053 54689 25087 54723
rect 21373 54621 21407 54655
rect 24777 54621 24811 54655
rect 32413 54621 32447 54655
rect 35352 54621 35386 54655
rect 35449 54621 35483 54655
rect 35724 54621 35758 54655
rect 35817 54621 35851 54655
rect 40141 54621 40175 54655
rect 21557 54553 21591 54587
rect 35541 54553 35575 54587
rect 41153 54553 41187 54587
rect 21741 54485 21775 54519
rect 24593 54485 24627 54519
rect 32321 54485 32355 54519
rect 32873 54485 32907 54519
rect 35173 54485 35207 54519
rect 38301 54485 38335 54519
rect 39405 54485 39439 54519
rect 40509 54485 40543 54519
rect 41353 54485 41387 54519
rect 58357 54485 58391 54519
rect 23029 54281 23063 54315
rect 24685 54281 24719 54315
rect 32698 54281 32732 54315
rect 37473 54281 37507 54315
rect 38853 54281 38887 54315
rect 40785 54281 40819 54315
rect 21281 54213 21315 54247
rect 23765 54213 23799 54247
rect 25053 54213 25087 54247
rect 27445 54213 27479 54247
rect 27537 54213 27571 54247
rect 31585 54213 31619 54247
rect 31769 54213 31803 54247
rect 34897 54213 34931 54247
rect 39681 54213 39715 54247
rect 40601 54213 40635 54247
rect 34667 54179 34701 54213
rect 1869 54145 1903 54179
rect 21097 54145 21131 54179
rect 23581 54145 23615 54179
rect 23857 54145 23891 54179
rect 24001 54145 24035 54179
rect 24864 54145 24898 54179
rect 24961 54145 24995 54179
rect 25181 54145 25215 54179
rect 25329 54145 25363 54179
rect 26341 54145 26375 54179
rect 26617 54145 26651 54179
rect 27348 54145 27382 54179
rect 27665 54145 27699 54179
rect 27813 54145 27847 54179
rect 31309 54145 31343 54179
rect 32321 54145 32355 54179
rect 32965 54145 32999 54179
rect 37657 54145 37691 54179
rect 37749 54145 37783 54179
rect 37933 54145 37967 54179
rect 38025 54145 38059 54179
rect 38577 54145 38611 54179
rect 40233 54145 40267 54179
rect 58357 54145 58391 54179
rect 26157 54077 26191 54111
rect 33977 54077 34011 54111
rect 1685 54009 1719 54043
rect 26525 54009 26559 54043
rect 34529 54009 34563 54043
rect 2421 53941 2455 53975
rect 21465 53941 21499 53975
rect 24133 53941 24167 53975
rect 27169 53941 27203 53975
rect 29561 53941 29595 53975
rect 31585 53941 31619 53975
rect 32689 53941 32723 53975
rect 33425 53941 33459 53975
rect 34713 53941 34747 53975
rect 40601 53941 40635 53975
rect 41245 53941 41279 53975
rect 58173 53941 58207 53975
rect 29193 53737 29227 53771
rect 37289 53737 37323 53771
rect 38669 53737 38703 53771
rect 40601 53737 40635 53771
rect 30113 53669 30147 53703
rect 28181 53601 28215 53635
rect 28641 53601 28675 53635
rect 36645 53601 36679 53635
rect 1869 53533 1903 53567
rect 2421 53533 2455 53567
rect 26893 53533 26927 53567
rect 27077 53533 27111 53567
rect 27313 53533 27347 53567
rect 29009 53533 29043 53567
rect 30021 53533 30055 53567
rect 30297 53533 30331 53567
rect 30573 53533 30607 53567
rect 31401 53533 31435 53567
rect 32229 53533 32263 53567
rect 32413 53533 32447 53567
rect 32781 53533 32815 53567
rect 37289 53533 37323 53567
rect 57713 53533 57747 53567
rect 58357 53533 58391 53567
rect 27169 53465 27203 53499
rect 27462 53465 27496 53499
rect 38393 53465 38427 53499
rect 40049 53465 40083 53499
rect 1685 53397 1719 53431
rect 26341 53397 26375 53431
rect 28825 53397 28859 53431
rect 31953 53397 31987 53431
rect 58173 53397 58207 53431
rect 29653 53193 29687 53227
rect 29837 53057 29871 53091
rect 30021 53057 30055 53091
rect 28273 52853 28307 52887
rect 29009 52853 29043 52887
rect 30021 52853 30055 52887
rect 38209 52853 38243 52887
rect 1685 52581 1719 52615
rect 58173 52581 58207 52615
rect 1869 52445 1903 52479
rect 2421 52445 2455 52479
rect 57713 52445 57747 52479
rect 58357 52445 58391 52479
rect 1869 51969 1903 52003
rect 57529 51969 57563 52003
rect 58357 51969 58391 52003
rect 1685 51765 1719 51799
rect 2421 51765 2455 51799
rect 58173 51765 58207 51799
rect 58357 51221 58391 51255
rect 1869 50881 1903 50915
rect 2421 50881 2455 50915
rect 58357 50881 58391 50915
rect 1685 50745 1719 50779
rect 58173 50677 58207 50711
rect 1869 50269 1903 50303
rect 57713 50269 57747 50303
rect 58357 50269 58391 50303
rect 1685 50133 1719 50167
rect 2421 50133 2455 50167
rect 58173 50133 58207 50167
rect 1869 49181 1903 49215
rect 57713 49181 57747 49215
rect 58357 49181 58391 49215
rect 1685 49045 1719 49079
rect 2421 49045 2455 49079
rect 58173 49045 58207 49079
rect 1869 48705 1903 48739
rect 57529 48705 57563 48739
rect 58357 48705 58391 48739
rect 1685 48501 1719 48535
rect 2421 48501 2455 48535
rect 58173 48501 58207 48535
rect 58357 47957 58391 47991
rect 1869 47617 1903 47651
rect 58357 47617 58391 47651
rect 1685 47481 1719 47515
rect 2421 47413 2455 47447
rect 58173 47413 58207 47447
rect 58173 47141 58207 47175
rect 1869 47005 1903 47039
rect 57713 47005 57747 47039
rect 58357 47005 58391 47039
rect 2421 46937 2455 46971
rect 1685 46869 1719 46903
rect 1869 45917 1903 45951
rect 2329 45917 2363 45951
rect 57713 45917 57747 45951
rect 58357 45917 58391 45951
rect 1685 45781 1719 45815
rect 58173 45781 58207 45815
rect 1869 45441 1903 45475
rect 57529 45441 57563 45475
rect 58357 45441 58391 45475
rect 1685 45237 1719 45271
rect 2421 45237 2455 45271
rect 58173 45237 58207 45271
rect 58357 44693 58391 44727
rect 1869 44353 1903 44387
rect 2329 44353 2363 44387
rect 58357 44353 58391 44387
rect 1685 44217 1719 44251
rect 58173 44149 58207 44183
rect 1869 43741 1903 43775
rect 57713 43741 57747 43775
rect 58357 43741 58391 43775
rect 1685 43605 1719 43639
rect 2421 43605 2455 43639
rect 58173 43605 58207 43639
rect 1869 42653 1903 42687
rect 57713 42653 57747 42687
rect 58357 42653 58391 42687
rect 1685 42517 1719 42551
rect 2421 42517 2455 42551
rect 58173 42517 58207 42551
rect 1869 42177 1903 42211
rect 57529 42177 57563 42211
rect 58357 42177 58391 42211
rect 1685 41973 1719 42007
rect 2421 41973 2455 42007
rect 58173 41973 58207 42007
rect 58357 41429 58391 41463
rect 1869 41089 1903 41123
rect 58357 41089 58391 41123
rect 1685 40953 1719 40987
rect 2421 40885 2455 40919
rect 58173 40885 58207 40919
rect 1869 40477 1903 40511
rect 57713 40477 57747 40511
rect 58357 40477 58391 40511
rect 1685 40341 1719 40375
rect 2421 40341 2455 40375
rect 58173 40341 58207 40375
rect 57529 39865 57563 39899
rect 58265 39797 58299 39831
rect 57621 39593 57655 39627
rect 1869 39389 1903 39423
rect 54953 39389 54987 39423
rect 56517 39389 56551 39423
rect 56609 39389 56643 39423
rect 58357 39389 58391 39423
rect 56149 39321 56183 39355
rect 56885 39321 56919 39355
rect 1685 39253 1719 39287
rect 2421 39253 2455 39287
rect 55597 39253 55631 39287
rect 55781 39253 55815 39287
rect 58173 39253 58207 39287
rect 58173 39049 58207 39083
rect 1869 38913 1903 38947
rect 58357 38913 58391 38947
rect 2421 38777 2455 38811
rect 1685 38709 1719 38743
rect 55413 38709 55447 38743
rect 56701 38709 56735 38743
rect 57529 38709 57563 38743
rect 56241 38505 56275 38539
rect 57437 38301 57471 38335
rect 57897 38301 57931 38335
rect 55781 38233 55815 38267
rect 57805 38233 57839 38267
rect 58173 38233 58207 38267
rect 56885 38165 56919 38199
rect 57069 38165 57103 38199
rect 54769 37961 54803 37995
rect 55873 37961 55907 37995
rect 56609 37961 56643 37995
rect 57529 37961 57563 37995
rect 58173 37961 58207 37995
rect 55137 37893 55171 37927
rect 1869 37825 1903 37859
rect 54033 37825 54067 37859
rect 55505 37825 55539 37859
rect 55597 37825 55631 37859
rect 58357 37825 58391 37859
rect 1685 37689 1719 37723
rect 2421 37621 2455 37655
rect 54585 37621 54619 37655
rect 56241 37417 56275 37451
rect 56885 37349 56919 37383
rect 54401 37281 54435 37315
rect 1869 37213 1903 37247
rect 57897 37213 57931 37247
rect 57437 37145 57471 37179
rect 57805 37145 57839 37179
rect 58173 37145 58207 37179
rect 1685 37077 1719 37111
rect 2421 37077 2455 37111
rect 57069 37077 57103 37111
rect 56701 36873 56735 36907
rect 58173 36873 58207 36907
rect 57529 36737 57563 36771
rect 58357 36737 58391 36771
rect 1869 36125 1903 36159
rect 57161 36125 57195 36159
rect 58357 36125 58391 36159
rect 1685 35989 1719 36023
rect 2421 35989 2455 36023
rect 57713 35989 57747 36023
rect 58173 35989 58207 36023
rect 56241 35785 56275 35819
rect 57529 35785 57563 35819
rect 1869 35649 1903 35683
rect 2421 35649 2455 35683
rect 58357 35649 58391 35683
rect 1685 35445 1719 35479
rect 58173 35445 58207 35479
rect 55873 35241 55907 35275
rect 56977 35105 57011 35139
rect 57136 35105 57170 35139
rect 57253 35105 57287 35139
rect 57529 35105 57563 35139
rect 58173 35105 58207 35139
rect 54585 35037 54619 35071
rect 54861 35037 54895 35071
rect 57989 35037 58023 35071
rect 56333 34969 56367 35003
rect 53941 34697 53975 34731
rect 54401 34697 54435 34731
rect 1869 34561 1903 34595
rect 52377 34561 52411 34595
rect 55204 34561 55238 34595
rect 56241 34561 56275 34595
rect 57529 34561 57563 34595
rect 58173 34561 58207 34595
rect 2421 34493 2455 34527
rect 52101 34493 52135 34527
rect 55045 34493 55079 34527
rect 55321 34493 55355 34527
rect 56057 34493 56091 34527
rect 56793 34493 56827 34527
rect 1685 34425 1719 34459
rect 55597 34425 55631 34459
rect 58357 34357 58391 34391
rect 54309 34153 54343 34187
rect 58173 34085 58207 34119
rect 1869 33949 1903 33983
rect 57161 33949 57195 33983
rect 58357 33949 58391 33983
rect 1685 33813 1719 33847
rect 57713 33813 57747 33847
rect 56241 33609 56275 33643
rect 56701 33609 56735 33643
rect 57529 33609 57563 33643
rect 58357 33473 58391 33507
rect 58173 33269 58207 33303
rect 55873 33065 55907 33099
rect 57161 32929 57195 32963
rect 57320 32929 57354 32963
rect 57713 32929 57747 32963
rect 58357 32929 58391 32963
rect 1869 32861 1903 32895
rect 57437 32861 57471 32895
rect 58173 32861 58207 32895
rect 1685 32725 1719 32759
rect 56517 32725 56551 32759
rect 56241 32521 56275 32555
rect 57345 32521 57379 32555
rect 56609 32453 56643 32487
rect 1869 32385 1903 32419
rect 55137 32385 55171 32419
rect 56977 32385 57011 32419
rect 57069 32385 57103 32419
rect 58357 32385 58391 32419
rect 54861 32317 54895 32351
rect 1685 32181 1719 32215
rect 56057 32181 56091 32215
rect 58173 32181 58207 32215
rect 55689 31977 55723 32011
rect 58357 31977 58391 32011
rect 57713 31909 57747 31943
rect 56977 31433 57011 31467
rect 1869 31297 1903 31331
rect 57529 31297 57563 31331
rect 58173 31297 58207 31331
rect 1685 31161 1719 31195
rect 58357 31093 58391 31127
rect 1869 30685 1903 30719
rect 57161 30685 57195 30719
rect 57529 30617 57563 30651
rect 57621 30617 57655 30651
rect 1685 30549 1719 30583
rect 56609 30549 56643 30583
rect 56793 30549 56827 30583
rect 57897 30549 57931 30583
rect 56425 30209 56459 30243
rect 58173 30209 58207 30243
rect 56885 30005 56919 30039
rect 57529 30005 57563 30039
rect 58357 30005 58391 30039
rect 57069 29665 57103 29699
rect 57621 29665 57655 29699
rect 58265 29665 58299 29699
rect 1869 29597 1903 29631
rect 2421 29597 2455 29631
rect 57207 29597 57241 29631
rect 57345 29597 57379 29631
rect 58081 29597 58115 29631
rect 1685 29461 1719 29495
rect 9965 29461 9999 29495
rect 10609 29461 10643 29495
rect 56425 29461 56459 29495
rect 9321 29257 9355 29291
rect 10701 29257 10735 29291
rect 58173 29257 58207 29291
rect 56977 29189 57011 29223
rect 1869 29121 1903 29155
rect 6929 29121 6963 29155
rect 8309 29121 8343 29155
rect 58357 29121 58391 29155
rect 7021 29053 7055 29087
rect 7205 29053 7239 29087
rect 9137 29053 9171 29087
rect 9229 29053 9263 29087
rect 1685 28985 1719 29019
rect 2421 28985 2455 29019
rect 7757 28985 7791 29019
rect 10241 28985 10275 29019
rect 57529 28985 57563 29019
rect 6561 28917 6595 28951
rect 9689 28917 9723 28951
rect 12449 28713 12483 28747
rect 58173 28713 58207 28747
rect 13737 28645 13771 28679
rect 57161 28645 57195 28679
rect 10517 28577 10551 28611
rect 13185 28577 13219 28611
rect 6561 28509 6595 28543
rect 10241 28509 10275 28543
rect 11621 28509 11655 28543
rect 13369 28509 13403 28543
rect 58357 28509 58391 28543
rect 6745 28373 6779 28407
rect 7481 28373 7515 28407
rect 9873 28373 9907 28407
rect 10333 28373 10367 28407
rect 11069 28373 11103 28407
rect 13277 28373 13311 28407
rect 14289 28373 14323 28407
rect 57621 28373 57655 28407
rect 57529 28169 57563 28203
rect 1869 28033 1903 28067
rect 9873 28033 9907 28067
rect 10333 28033 10367 28067
rect 15393 28033 15427 28067
rect 58357 28033 58391 28067
rect 1685 27897 1719 27931
rect 58173 27897 58207 27931
rect 2421 27829 2455 27863
rect 5917 27829 5951 27863
rect 7113 27829 7147 27863
rect 9689 27829 9723 27863
rect 10517 27829 10551 27863
rect 13829 27829 13863 27863
rect 14473 27829 14507 27863
rect 15577 27829 15611 27863
rect 5733 27625 5767 27659
rect 10517 27625 10551 27659
rect 2421 27557 2455 27591
rect 6929 27557 6963 27591
rect 7573 27557 7607 27591
rect 14289 27557 14323 27591
rect 57713 27557 57747 27591
rect 58173 27557 58207 27591
rect 5181 27489 5215 27523
rect 6285 27489 6319 27523
rect 13369 27489 13403 27523
rect 13553 27489 13587 27523
rect 57161 27489 57195 27523
rect 1869 27421 1903 27455
rect 5365 27421 5399 27455
rect 6561 27421 6595 27455
rect 7389 27421 7423 27455
rect 58357 27421 58391 27455
rect 5273 27353 5307 27387
rect 12173 27353 12207 27387
rect 1685 27285 1719 27319
rect 6469 27285 6503 27319
rect 8125 27285 8159 27319
rect 9873 27285 9907 27319
rect 11621 27285 11655 27319
rect 12909 27285 12943 27319
rect 13277 27285 13311 27319
rect 14841 27285 14875 27319
rect 15393 27285 15427 27319
rect 5457 27081 5491 27115
rect 8861 27081 8895 27115
rect 9321 27081 9355 27115
rect 11161 27081 11195 27115
rect 14565 27081 14599 27115
rect 58357 27081 58391 27115
rect 4353 27013 4387 27047
rect 9229 27013 9263 27047
rect 13461 27013 13495 27047
rect 15209 27013 15243 27047
rect 6561 26945 6595 26979
rect 8217 26945 8251 26979
rect 10793 26945 10827 26979
rect 11713 26945 11747 26979
rect 12357 26945 12391 26979
rect 13369 26945 13403 26979
rect 14749 26945 14783 26979
rect 3801 26877 3835 26911
rect 9505 26877 9539 26911
rect 10609 26877 10643 26911
rect 10701 26877 10735 26911
rect 13645 26877 13679 26911
rect 17049 26877 17083 26911
rect 7205 26809 7239 26843
rect 11897 26809 11931 26843
rect 2053 26741 2087 26775
rect 5917 26741 5951 26775
rect 6745 26741 6779 26775
rect 8401 26741 8435 26775
rect 12541 26741 12575 26775
rect 13001 26741 13035 26775
rect 15761 26741 15795 26775
rect 17601 26741 17635 26775
rect 56977 26741 57011 26775
rect 57529 26741 57563 26775
rect 10057 26537 10091 26571
rect 11345 26537 11379 26571
rect 12633 26537 12667 26571
rect 14749 26537 14783 26571
rect 1685 26469 1719 26503
rect 4721 26469 4755 26503
rect 5917 26469 5951 26503
rect 8585 26469 8619 26503
rect 12081 26469 12115 26503
rect 2789 26401 2823 26435
rect 4077 26401 4111 26435
rect 4261 26401 4295 26435
rect 6469 26401 6503 26435
rect 6653 26401 6687 26435
rect 7573 26401 7607 26435
rect 13645 26401 13679 26435
rect 15209 26401 15243 26435
rect 15301 26401 15335 26435
rect 16497 26401 16531 26435
rect 17785 26401 17819 26435
rect 57320 26401 57354 26435
rect 57437 26401 57471 26435
rect 57713 26401 57747 26435
rect 58357 26401 58391 26435
rect 1869 26333 1903 26367
rect 2973 26333 3007 26367
rect 5733 26333 5767 26367
rect 11897 26333 11931 26367
rect 13185 26333 13219 26367
rect 15117 26333 15151 26367
rect 17601 26333 17635 26367
rect 44557 26333 44591 26367
rect 56517 26333 56551 26367
rect 57161 26333 57195 26367
rect 58173 26333 58207 26367
rect 3065 26265 3099 26299
rect 4353 26265 4387 26299
rect 5273 26265 5307 26299
rect 9137 26265 9171 26299
rect 16313 26265 16347 26299
rect 18429 26265 18463 26299
rect 3433 26197 3467 26231
rect 6745 26197 6779 26231
rect 7113 26197 7147 26231
rect 15945 26197 15979 26231
rect 16405 26197 16439 26231
rect 17141 26197 17175 26231
rect 17509 26197 17543 26231
rect 44373 26197 44407 26231
rect 57345 25993 57379 26027
rect 58173 25993 58207 26027
rect 8125 25925 8159 25959
rect 56333 25925 56367 25959
rect 2421 25857 2455 25891
rect 3709 25857 3743 25891
rect 4813 25857 4847 25891
rect 7205 25857 7239 25891
rect 8217 25857 8251 25891
rect 9689 25857 9723 25891
rect 10517 25857 10551 25891
rect 10609 25857 10643 25891
rect 11713 25857 11747 25891
rect 13369 25857 13403 25891
rect 14197 25857 14231 25891
rect 16037 25857 16071 25891
rect 17049 25857 17083 25891
rect 56885 25857 56919 25891
rect 57529 25857 57563 25891
rect 58357 25857 58391 25891
rect 2145 25789 2179 25823
rect 2329 25789 2363 25823
rect 8033 25789 8067 25823
rect 10701 25789 10735 25823
rect 14289 25789 14323 25823
rect 14473 25789 14507 25823
rect 6745 25721 6779 25755
rect 10149 25721 10183 25755
rect 13829 25721 13863 25755
rect 15853 25721 15887 25755
rect 2789 25653 2823 25687
rect 3893 25653 3927 25687
rect 7389 25653 7423 25687
rect 8585 25653 8619 25687
rect 9505 25653 9539 25687
rect 13185 25653 13219 25687
rect 15393 25653 15427 25687
rect 16865 25653 16899 25687
rect 17601 25653 17635 25687
rect 1685 25449 1719 25483
rect 3157 25449 3191 25483
rect 7389 25449 7423 25483
rect 8493 25449 8527 25483
rect 11713 25449 11747 25483
rect 14473 25449 14507 25483
rect 2605 25381 2639 25415
rect 9321 25381 9355 25415
rect 57320 25313 57354 25347
rect 57437 25313 57471 25347
rect 57713 25313 57747 25347
rect 58357 25313 58391 25347
rect 1869 25245 1903 25279
rect 2421 25245 2455 25279
rect 9137 25245 9171 25279
rect 57161 25245 57195 25279
rect 58173 25245 58207 25279
rect 11161 25109 11195 25143
rect 15025 25109 15059 25143
rect 15577 25109 15611 25143
rect 16773 25109 16807 25143
rect 56517 25109 56551 25143
rect 1869 24769 1903 24803
rect 58357 24769 58391 24803
rect 2881 24701 2915 24735
rect 1685 24633 1719 24667
rect 57437 24633 57471 24667
rect 58173 24633 58207 24667
rect 2329 24565 2363 24599
rect 3525 24565 3559 24599
rect 56977 24565 57011 24599
rect 2881 24361 2915 24395
rect 19533 24361 19567 24395
rect 57713 24361 57747 24395
rect 58173 24293 58207 24327
rect 1869 24157 1903 24191
rect 57161 24157 57195 24191
rect 58357 24157 58391 24191
rect 19809 24089 19843 24123
rect 1685 24021 1719 24055
rect 2421 24021 2455 24055
rect 20453 24021 20487 24055
rect 58357 23817 58391 23851
rect 3249 23749 3283 23783
rect 5549 23749 5583 23783
rect 9413 23749 9447 23783
rect 2329 23681 2363 23715
rect 2145 23613 2179 23647
rect 2237 23613 2271 23647
rect 4077 23613 4111 23647
rect 5825 23613 5859 23647
rect 7941 23613 7975 23647
rect 9689 23613 9723 23647
rect 2697 23477 2731 23511
rect 10701 23273 10735 23307
rect 2513 23205 2547 23239
rect 4905 23205 4939 23239
rect 6377 23137 6411 23171
rect 6653 23137 6687 23171
rect 12173 23137 12207 23171
rect 58081 23137 58115 23171
rect 1869 23069 1903 23103
rect 2329 23069 2363 23103
rect 2973 23069 3007 23103
rect 12449 23069 12483 23103
rect 57805 23069 57839 23103
rect 1685 22933 1719 22967
rect 3157 22933 3191 22967
rect 4077 22933 4111 22967
rect 18429 22933 18463 22967
rect 2237 22729 2271 22763
rect 2697 22729 2731 22763
rect 3249 22729 3283 22763
rect 8401 22729 8435 22763
rect 14197 22729 14231 22763
rect 18797 22729 18831 22763
rect 58173 22729 58207 22763
rect 2329 22661 2363 22695
rect 12725 22661 12759 22695
rect 19165 22661 19199 22695
rect 10149 22593 10183 22627
rect 12449 22593 12483 22627
rect 18337 22593 18371 22627
rect 57529 22593 57563 22627
rect 58357 22593 58391 22627
rect 2145 22525 2179 22559
rect 9873 22525 9907 22559
rect 19257 22525 19291 22559
rect 19441 22525 19475 22559
rect 18153 22389 18187 22423
rect 20085 22389 20119 22423
rect 1685 22185 1719 22219
rect 6297 22185 6331 22219
rect 15288 22185 15322 22219
rect 2789 22049 2823 22083
rect 16773 22049 16807 22083
rect 1869 21981 1903 22015
rect 6561 21981 6595 22015
rect 15025 21981 15059 22015
rect 57713 21981 57747 22015
rect 58357 21981 58391 22015
rect 4813 21845 4847 21879
rect 18705 21845 18739 21879
rect 58173 21845 58207 21879
rect 58173 21641 58207 21675
rect 19349 21573 19383 21607
rect 1869 21505 1903 21539
rect 15577 21505 15611 21539
rect 19625 21505 19659 21539
rect 57529 21505 57563 21539
rect 58357 21505 58391 21539
rect 15301 21437 15335 21471
rect 1685 21369 1719 21403
rect 2881 21301 2915 21335
rect 13829 21301 13863 21335
rect 20177 21301 20211 21335
rect 11989 21097 12023 21131
rect 17049 21097 17083 21131
rect 18245 21097 18279 21131
rect 58173 21097 58207 21131
rect 2145 20961 2179 20995
rect 13737 20961 13771 20995
rect 15301 20961 15335 20995
rect 15577 20961 15611 20995
rect 19901 20961 19935 20995
rect 20085 20961 20119 20995
rect 2329 20893 2363 20927
rect 18889 20893 18923 20927
rect 19809 20893 19843 20927
rect 57713 20893 57747 20927
rect 58357 20893 58391 20927
rect 2237 20825 2271 20859
rect 13461 20825 13495 20859
rect 2697 20757 2731 20791
rect 3249 20757 3283 20791
rect 19441 20757 19475 20791
rect 20637 20757 20671 20791
rect 1685 20553 1719 20587
rect 4261 20553 4295 20587
rect 10885 20553 10919 20587
rect 19441 20553 19475 20587
rect 1869 20417 1903 20451
rect 2329 20417 2363 20451
rect 18705 20417 18739 20451
rect 19533 20417 19567 20451
rect 5733 20349 5767 20383
rect 6009 20349 6043 20383
rect 9137 20349 9171 20383
rect 9413 20349 9447 20383
rect 19257 20349 19291 20383
rect 2513 20281 2547 20315
rect 18521 20213 18555 20247
rect 19901 20213 19935 20247
rect 20453 20213 20487 20247
rect 17141 20009 17175 20043
rect 18797 20009 18831 20043
rect 15393 19873 15427 19907
rect 15669 19873 15703 19907
rect 1869 19805 1903 19839
rect 57713 19805 57747 19839
rect 58357 19805 58391 19839
rect 5733 19737 5767 19771
rect 6377 19737 6411 19771
rect 1685 19669 1719 19703
rect 5825 19669 5859 19703
rect 19533 19669 19567 19703
rect 58173 19669 58207 19703
rect 4261 19465 4295 19499
rect 9505 19465 9539 19499
rect 14657 19465 14691 19499
rect 58173 19465 58207 19499
rect 1869 19329 1903 19363
rect 6009 19329 6043 19363
rect 7757 19329 7791 19363
rect 12909 19329 12943 19363
rect 58357 19329 58391 19363
rect 5733 19261 5767 19295
rect 8033 19261 8067 19295
rect 13185 19261 13219 19295
rect 57253 19261 57287 19295
rect 57529 19261 57563 19295
rect 1685 19125 1719 19159
rect 10885 18921 10919 18955
rect 58357 18921 58391 18955
rect 20177 18853 20211 18887
rect 12633 18785 12667 18819
rect 15117 18785 15151 18819
rect 15393 18785 15427 18819
rect 17141 18785 17175 18819
rect 1869 18717 1903 18751
rect 2329 18717 2363 18751
rect 19717 18717 19751 18751
rect 20361 18717 20395 18751
rect 12357 18649 12391 18683
rect 1685 18581 1719 18615
rect 2513 18581 2547 18615
rect 2973 18581 3007 18615
rect 19533 18581 19567 18615
rect 2329 18377 2363 18411
rect 2697 18377 2731 18411
rect 7481 18377 7515 18411
rect 12173 18377 12207 18411
rect 18981 18377 19015 18411
rect 19809 18377 19843 18411
rect 20269 18377 20303 18411
rect 3157 18309 3191 18343
rect 14749 18309 14783 18343
rect 12357 18241 12391 18275
rect 13001 18241 13035 18275
rect 19901 18241 19935 18275
rect 57529 18241 57563 18275
rect 58357 18241 58391 18275
rect 2145 18173 2179 18207
rect 2237 18173 2271 18207
rect 5733 18173 5767 18207
rect 6009 18173 6043 18207
rect 8953 18173 8987 18207
rect 9229 18173 9263 18207
rect 19717 18173 19751 18207
rect 4261 18105 4295 18139
rect 11069 18037 11103 18071
rect 20729 18037 20763 18071
rect 58173 18037 58207 18071
rect 11897 17833 11931 17867
rect 17141 17833 17175 17867
rect 21465 17833 21499 17867
rect 2053 17697 2087 17731
rect 2237 17697 2271 17731
rect 13369 17697 13403 17731
rect 15669 17697 15703 17731
rect 20269 17697 20303 17731
rect 2329 17629 2363 17663
rect 13645 17629 13679 17663
rect 15393 17629 15427 17663
rect 21649 17629 21683 17663
rect 57713 17629 57747 17663
rect 58357 17629 58391 17663
rect 19993 17561 20027 17595
rect 2697 17493 2731 17527
rect 3249 17493 3283 17527
rect 19625 17493 19659 17527
rect 20085 17493 20119 17527
rect 20913 17493 20947 17527
rect 58173 17493 58207 17527
rect 1685 17289 1719 17323
rect 8309 17289 8343 17323
rect 19533 17289 19567 17323
rect 1869 17153 1903 17187
rect 2329 17153 2363 17187
rect 9597 17153 9631 17187
rect 2513 16949 2547 16983
rect 2973 16949 3007 16983
rect 21189 16745 21223 16779
rect 21741 16745 21775 16779
rect 5917 16609 5951 16643
rect 9137 16609 9171 16643
rect 9413 16609 9447 16643
rect 22201 16609 22235 16643
rect 22293 16609 22327 16643
rect 1869 16541 1903 16575
rect 2329 16541 2363 16575
rect 6193 16541 6227 16575
rect 19625 16541 19659 16575
rect 20269 16541 20303 16575
rect 20545 16541 20579 16575
rect 57713 16541 57747 16575
rect 58357 16541 58391 16575
rect 1685 16405 1719 16439
rect 4445 16405 4479 16439
rect 10885 16405 10919 16439
rect 19441 16405 19475 16439
rect 22109 16405 22143 16439
rect 58173 16405 58207 16439
rect 8309 16201 8343 16235
rect 1869 16065 1903 16099
rect 9597 16065 9631 16099
rect 13001 16065 13035 16099
rect 58357 16065 58391 16099
rect 1685 15861 1719 15895
rect 2881 15861 2915 15895
rect 3341 15861 3375 15895
rect 14289 15861 14323 15895
rect 58173 15861 58207 15895
rect 3249 15657 3283 15691
rect 10517 15657 10551 15691
rect 17141 15657 17175 15691
rect 58357 15657 58391 15691
rect 4353 15589 4387 15623
rect 2145 15521 2179 15555
rect 2237 15521 2271 15555
rect 5825 15521 5859 15555
rect 6101 15521 6135 15555
rect 15393 15521 15427 15555
rect 15669 15521 15703 15555
rect 12265 15453 12299 15487
rect 2329 15385 2363 15419
rect 11989 15385 12023 15419
rect 2697 15317 2731 15351
rect 2513 15113 2547 15147
rect 5549 15113 5583 15147
rect 6561 15113 6595 15147
rect 8953 15113 8987 15147
rect 5825 15045 5859 15079
rect 7481 15045 7515 15079
rect 1869 14977 1903 15011
rect 2329 14977 2363 15011
rect 7205 14977 7239 15011
rect 20177 14977 20211 15011
rect 57529 14977 57563 15011
rect 58357 14977 58391 15011
rect 3065 14909 3099 14943
rect 20269 14909 20303 14943
rect 20453 14909 20487 14943
rect 1685 14841 1719 14875
rect 19349 14773 19383 14807
rect 19809 14773 19843 14807
rect 58173 14773 58207 14807
rect 22293 14501 22327 14535
rect 2145 14433 2179 14467
rect 10517 14433 10551 14467
rect 12265 14433 12299 14467
rect 12541 14433 12575 14467
rect 15761 14433 15795 14467
rect 16037 14433 16071 14467
rect 17785 14433 17819 14467
rect 20545 14433 20579 14467
rect 21097 14433 21131 14467
rect 22477 14365 22511 14399
rect 57713 14365 57747 14399
rect 58357 14365 58391 14399
rect 2329 14297 2363 14331
rect 3157 14297 3191 14331
rect 20361 14297 20395 14331
rect 2237 14229 2271 14263
rect 2697 14229 2731 14263
rect 18797 14229 18831 14263
rect 19901 14229 19935 14263
rect 20269 14229 20303 14263
rect 58173 14229 58207 14263
rect 1685 14025 1719 14059
rect 2513 14025 2547 14059
rect 11069 14025 11103 14059
rect 13829 14025 13863 14059
rect 19717 14025 19751 14059
rect 22201 14025 22235 14059
rect 23489 14025 23523 14059
rect 11713 13957 11747 13991
rect 56793 13957 56827 13991
rect 58265 13957 58299 13991
rect 1869 13889 1903 13923
rect 2329 13889 2363 13923
rect 12081 13889 12115 13923
rect 15577 13889 15611 13923
rect 19901 13889 19935 13923
rect 22569 13889 22603 13923
rect 56517 13889 56551 13923
rect 2973 13821 3007 13855
rect 15301 13821 15335 13855
rect 22661 13821 22695 13855
rect 22845 13821 22879 13855
rect 56057 13821 56091 13855
rect 16221 13481 16255 13515
rect 22109 13481 22143 13515
rect 22569 13481 22603 13515
rect 4353 13413 4387 13447
rect 5825 13345 5859 13379
rect 11713 13345 11747 13379
rect 17693 13345 17727 13379
rect 57161 13345 57195 13379
rect 57320 13345 57354 13379
rect 57437 13345 57471 13379
rect 57713 13345 57747 13379
rect 58173 13345 58207 13379
rect 1869 13277 1903 13311
rect 6101 13277 6135 13311
rect 13737 13277 13771 13311
rect 17969 13277 18003 13311
rect 19901 13277 19935 13311
rect 58357 13277 58391 13311
rect 13461 13209 13495 13243
rect 1685 13141 1719 13175
rect 2421 13141 2455 13175
rect 19717 13141 19751 13175
rect 56517 13141 56551 13175
rect 3617 12937 3651 12971
rect 9873 12937 9907 12971
rect 22937 12937 22971 12971
rect 23673 12937 23707 12971
rect 57437 12937 57471 12971
rect 3065 12869 3099 12903
rect 8401 12869 8435 12903
rect 1869 12801 1903 12835
rect 11161 12801 11195 12835
rect 11713 12801 11747 12835
rect 20177 12801 20211 12835
rect 22845 12801 22879 12835
rect 58357 12801 58391 12835
rect 2329 12733 2363 12767
rect 8125 12733 8159 12767
rect 20269 12733 20303 12767
rect 20453 12733 20487 12767
rect 23121 12733 23155 12767
rect 1685 12597 1719 12631
rect 13001 12597 13035 12631
rect 18705 12597 18739 12631
rect 19349 12597 19383 12631
rect 19809 12597 19843 12631
rect 22477 12597 22511 12631
rect 58173 12597 58207 12631
rect 3341 12393 3375 12427
rect 7585 12393 7619 12427
rect 22477 12393 22511 12427
rect 57713 12393 57747 12427
rect 6101 12325 6135 12359
rect 2145 12257 2179 12291
rect 3985 12257 4019 12291
rect 14933 12257 14967 12291
rect 16681 12257 16715 12291
rect 2237 12189 2271 12223
rect 2329 12189 2363 12223
rect 3157 12189 3191 12223
rect 7849 12189 7883 12223
rect 16957 12189 16991 12223
rect 19809 12189 19843 12223
rect 22661 12189 22695 12223
rect 57161 12189 57195 12223
rect 58357 12189 58391 12223
rect 2697 12053 2731 12087
rect 19625 12053 19659 12087
rect 58173 12053 58207 12087
rect 2329 11849 2363 11883
rect 11989 11849 12023 11883
rect 19349 11849 19383 11883
rect 20269 11849 20303 11883
rect 2421 11781 2455 11815
rect 10793 11781 10827 11815
rect 3249 11713 3283 11747
rect 5917 11713 5951 11747
rect 20177 11713 20211 11747
rect 22845 11713 22879 11747
rect 56333 11713 56367 11747
rect 56609 11713 56643 11747
rect 58357 11713 58391 11747
rect 2237 11645 2271 11679
rect 5641 11645 5675 11679
rect 8769 11645 8803 11679
rect 9045 11645 9079 11679
rect 13461 11645 13495 11679
rect 13737 11645 13771 11679
rect 20361 11645 20395 11679
rect 22937 11645 22971 11679
rect 23121 11645 23155 11679
rect 23673 11645 23707 11679
rect 56492 11645 56526 11679
rect 57345 11645 57379 11679
rect 57529 11645 57563 11679
rect 2789 11577 2823 11611
rect 3433 11577 3467 11611
rect 56885 11577 56919 11611
rect 4169 11509 4203 11543
rect 19809 11509 19843 11543
rect 21373 11509 21407 11543
rect 22477 11509 22511 11543
rect 55689 11509 55723 11543
rect 58173 11509 58207 11543
rect 1685 11305 1719 11339
rect 2605 11305 2639 11339
rect 19717 11305 19751 11339
rect 20637 11305 20671 11339
rect 57161 11305 57195 11339
rect 22385 11237 22419 11271
rect 58173 11237 58207 11271
rect 57621 11169 57655 11203
rect 1869 11101 1903 11135
rect 3157 11101 3191 11135
rect 19901 11101 19935 11135
rect 22569 11101 22603 11135
rect 58357 11101 58391 11135
rect 1685 10761 1719 10795
rect 8309 10761 8343 10795
rect 57529 10761 57563 10795
rect 58357 10761 58391 10795
rect 9597 10693 9631 10727
rect 13001 10693 13035 10727
rect 17141 10693 17175 10727
rect 18889 10693 18923 10727
rect 1869 10625 1903 10659
rect 20269 10625 20303 10659
rect 55321 10625 55355 10659
rect 14749 10557 14783 10591
rect 16865 10557 16899 10591
rect 20361 10557 20395 10591
rect 20453 10557 20487 10591
rect 2421 10421 2455 10455
rect 19349 10421 19383 10455
rect 19901 10421 19935 10455
rect 55137 10421 55171 10455
rect 2421 10217 2455 10251
rect 12081 10217 12115 10251
rect 16313 10217 16347 10251
rect 18061 10081 18095 10115
rect 23213 10081 23247 10115
rect 1869 10013 1903 10047
rect 19901 10013 19935 10047
rect 57161 10013 57195 10047
rect 17785 9945 17819 9979
rect 22109 9945 22143 9979
rect 23029 9945 23063 9979
rect 57529 9945 57563 9979
rect 57621 9945 57655 9979
rect 57897 9945 57931 9979
rect 1685 9877 1719 9911
rect 2973 9877 3007 9911
rect 19717 9877 19751 9911
rect 22569 9877 22603 9911
rect 22937 9877 22971 9911
rect 56609 9877 56643 9911
rect 56793 9877 56827 9911
rect 2513 9673 2547 9707
rect 55689 9605 55723 9639
rect 56241 9605 56275 9639
rect 56609 9605 56643 9639
rect 3341 9537 3375 9571
rect 6653 9537 6687 9571
rect 7389 9537 7423 9571
rect 12173 9537 12207 9571
rect 22661 9537 22695 9571
rect 57437 9537 57471 9571
rect 58173 9537 58207 9571
rect 2237 9469 2271 9503
rect 2421 9469 2455 9503
rect 10057 9469 10091 9503
rect 2881 9401 2915 9435
rect 6837 9401 6871 9435
rect 12357 9401 12391 9435
rect 58357 9401 58391 9435
rect 3525 9333 3559 9367
rect 3985 9333 4019 9367
rect 19533 9333 19567 9367
rect 22477 9333 22511 9367
rect 4905 9129 4939 9163
rect 14473 9129 14507 9163
rect 15963 9129 15997 9163
rect 21005 9129 21039 9163
rect 57161 9129 57195 9163
rect 58173 9129 58207 9163
rect 57621 9061 57655 9095
rect 2421 8993 2455 9027
rect 6377 8993 6411 9027
rect 9597 8993 9631 9027
rect 9781 8993 9815 9027
rect 10977 8993 11011 9027
rect 16221 8993 16255 9027
rect 20177 8993 20211 9027
rect 20361 8993 20395 9027
rect 23121 8993 23155 9027
rect 2605 8925 2639 8959
rect 6653 8925 6687 8959
rect 8585 8925 8619 8959
rect 13001 8925 13035 8959
rect 22845 8925 22879 8959
rect 58357 8925 58391 8959
rect 9505 8857 9539 8891
rect 12725 8857 12759 8891
rect 22937 8857 22971 8891
rect 2513 8789 2547 8823
rect 2973 8789 3007 8823
rect 3985 8789 4019 8823
rect 8401 8789 8435 8823
rect 9137 8789 9171 8823
rect 10425 8789 10459 8823
rect 19717 8789 19751 8823
rect 20085 8789 20119 8823
rect 21925 8789 21959 8823
rect 22477 8789 22511 8823
rect 1685 8585 1719 8619
rect 11713 8585 11747 8619
rect 18705 8585 18739 8619
rect 19717 8585 19751 8619
rect 57529 8585 57563 8619
rect 3341 8517 3375 8551
rect 8309 8517 8343 8551
rect 13185 8517 13219 8551
rect 19809 8517 19843 8551
rect 1869 8449 1903 8483
rect 2605 8449 2639 8483
rect 18889 8449 18923 8483
rect 22569 8449 22603 8483
rect 56977 8449 57011 8483
rect 58357 8449 58391 8483
rect 8033 8381 8067 8415
rect 9781 8381 9815 8415
rect 13461 8381 13495 8415
rect 19901 8381 19935 8415
rect 20545 8381 20579 8415
rect 2789 8313 2823 8347
rect 18153 8313 18187 8347
rect 19349 8313 19383 8347
rect 22385 8313 22419 8347
rect 58173 8313 58207 8347
rect 1685 8041 1719 8075
rect 3157 8041 3191 8075
rect 19533 8041 19567 8075
rect 23397 8041 23431 8075
rect 57161 7973 57195 8007
rect 5181 7905 5215 7939
rect 6653 7905 6687 7939
rect 22753 7905 22787 7939
rect 57437 7905 57471 7939
rect 57575 7905 57609 7939
rect 57713 7905 57747 7939
rect 1869 7837 1903 7871
rect 2605 7837 2639 7871
rect 6929 7837 6963 7871
rect 19717 7837 19751 7871
rect 56517 7837 56551 7871
rect 56701 7837 56735 7871
rect 22569 7769 22603 7803
rect 2421 7701 2455 7735
rect 18797 7701 18831 7735
rect 21557 7701 21591 7735
rect 22109 7701 22143 7735
rect 22477 7701 22511 7735
rect 58357 7701 58391 7735
rect 2881 7497 2915 7531
rect 3985 7497 4019 7531
rect 18613 7497 18647 7531
rect 58173 7497 58207 7531
rect 9597 7429 9631 7463
rect 13001 7429 13035 7463
rect 56977 7429 57011 7463
rect 2513 7361 2547 7395
rect 3341 7361 3375 7395
rect 22109 7361 22143 7395
rect 23121 7361 23155 7395
rect 23765 7361 23799 7395
rect 56425 7361 56459 7395
rect 58357 7361 58391 7395
rect 2329 7293 2363 7327
rect 2421 7293 2455 7327
rect 7849 7293 7883 7327
rect 14749 7293 14783 7327
rect 16865 7293 16899 7327
rect 17141 7293 17175 7327
rect 23397 7293 23431 7327
rect 57437 7293 57471 7327
rect 3525 7157 3559 7191
rect 19165 7157 19199 7191
rect 22661 7157 22695 7191
rect 5561 6953 5595 6987
rect 23489 6953 23523 6987
rect 4077 6885 4111 6919
rect 56885 6885 56919 6919
rect 2237 6817 2271 6851
rect 3249 6817 3283 6851
rect 19901 6817 19935 6851
rect 20085 6817 20119 6851
rect 20637 6817 20671 6851
rect 22017 6817 22051 6851
rect 56333 6817 56367 6851
rect 56609 6817 56643 6851
rect 5825 6749 5859 6783
rect 18797 6749 18831 6783
rect 19809 6749 19843 6783
rect 21373 6749 21407 6783
rect 23029 6749 23063 6783
rect 23949 6749 23983 6783
rect 24593 6749 24627 6783
rect 56471 6749 56505 6783
rect 57345 6749 57379 6783
rect 57529 6749 57563 6783
rect 58357 6749 58391 6783
rect 2421 6681 2455 6715
rect 22201 6681 22235 6715
rect 2329 6613 2363 6647
rect 2789 6613 2823 6647
rect 19441 6613 19475 6647
rect 21189 6613 21223 6647
rect 22109 6613 22143 6647
rect 22569 6613 22603 6647
rect 55689 6613 55723 6647
rect 58173 6613 58207 6647
rect 1685 6409 1719 6443
rect 3157 6409 3191 6443
rect 21373 6409 21407 6443
rect 56977 6409 57011 6443
rect 57437 6409 57471 6443
rect 7849 6341 7883 6375
rect 13829 6341 13863 6375
rect 15577 6341 15611 6375
rect 56425 6341 56459 6375
rect 1869 6273 1903 6307
rect 2513 6273 2547 6307
rect 19441 6273 19475 6307
rect 20085 6273 20119 6307
rect 22569 6273 22603 6307
rect 23029 6273 23063 6307
rect 23581 6273 23615 6307
rect 24225 6273 24259 6307
rect 55873 6273 55907 6307
rect 58357 6273 58391 6307
rect 9597 6205 9631 6239
rect 9873 6205 9907 6239
rect 15853 6205 15887 6239
rect 22385 6137 22419 6171
rect 2697 6069 2731 6103
rect 19257 6069 19291 6103
rect 19901 6069 19935 6103
rect 23121 6069 23155 6103
rect 58173 6069 58207 6103
rect 1685 5865 1719 5899
rect 19809 5865 19843 5899
rect 22661 5865 22695 5899
rect 5641 5797 5675 5831
rect 10149 5797 10183 5831
rect 16773 5797 16807 5831
rect 57161 5797 57195 5831
rect 7113 5729 7147 5763
rect 7389 5729 7423 5763
rect 11621 5729 11655 5763
rect 20453 5729 20487 5763
rect 56517 5729 56551 5763
rect 57437 5729 57471 5763
rect 57575 5729 57609 5763
rect 1869 5661 1903 5695
rect 11897 5661 11931 5695
rect 18521 5661 18555 5695
rect 20177 5661 20211 5695
rect 56701 5661 56735 5695
rect 57713 5661 57747 5695
rect 18245 5593 18279 5627
rect 20269 5525 20303 5559
rect 21005 5525 21039 5559
rect 23213 5525 23247 5559
rect 58357 5525 58391 5559
rect 11897 5321 11931 5355
rect 19257 5321 19291 5355
rect 20269 5321 20303 5355
rect 56977 5321 57011 5355
rect 57437 5321 57471 5355
rect 58173 5321 58207 5355
rect 13369 5253 13403 5287
rect 1869 5185 1903 5219
rect 13645 5185 13679 5219
rect 19441 5185 19475 5219
rect 56425 5185 56459 5219
rect 58357 5185 58391 5219
rect 20361 5117 20395 5151
rect 20453 5117 20487 5151
rect 1685 5049 1719 5083
rect 19901 5049 19935 5083
rect 22753 4981 22787 5015
rect 3065 4777 3099 4811
rect 19717 4777 19751 4811
rect 56517 4777 56551 4811
rect 57529 4777 57563 4811
rect 58173 4777 58207 4811
rect 1869 4573 1903 4607
rect 57069 4573 57103 4607
rect 57713 4573 57747 4607
rect 58357 4573 58391 4607
rect 55965 4505 55999 4539
rect 1685 4437 1719 4471
rect 20269 4437 20303 4471
rect 21097 4437 21131 4471
rect 22753 4437 22787 4471
rect 2605 4233 2639 4267
rect 2973 4233 3007 4267
rect 19257 4233 19291 4267
rect 20085 4233 20119 4267
rect 22937 4165 22971 4199
rect 3433 4097 3467 4131
rect 6561 4097 6595 4131
rect 20177 4097 20211 4131
rect 21373 4097 21407 4131
rect 55781 4097 55815 4131
rect 56885 4097 56919 4131
rect 57529 4097 57563 4131
rect 58265 4097 58299 4131
rect 2421 4029 2455 4063
rect 2513 4029 2547 4063
rect 4169 4029 4203 4063
rect 20361 4029 20395 4063
rect 21097 4029 21131 4063
rect 23029 4029 23063 4063
rect 23213 4029 23247 4063
rect 18153 3961 18187 3995
rect 22017 3961 22051 3995
rect 57345 3961 57379 3995
rect 1777 3893 1811 3927
rect 3617 3893 3651 3927
rect 4629 3893 4663 3927
rect 6745 3893 6779 3927
rect 17601 3893 17635 3927
rect 18613 3893 18647 3927
rect 19717 3893 19751 3927
rect 22569 3893 22603 3927
rect 55321 3893 55355 3927
rect 58081 3893 58115 3927
rect 4997 3689 5031 3723
rect 7297 3689 7331 3723
rect 11345 3689 11379 3723
rect 13645 3689 13679 3723
rect 16405 3689 16439 3723
rect 40877 3689 40911 3723
rect 48697 3689 48731 3723
rect 4169 3621 4203 3655
rect 2421 3553 2455 3587
rect 6469 3553 6503 3587
rect 9873 3553 9907 3587
rect 20085 3553 20119 3587
rect 21465 3553 21499 3587
rect 23029 3553 23063 3587
rect 23213 3553 23247 3587
rect 23765 3553 23799 3587
rect 54033 3553 54067 3587
rect 2513 3485 2547 3519
rect 3985 3485 4019 3519
rect 6745 3485 6779 3519
rect 9597 3485 9631 3519
rect 14381 3485 14415 3519
rect 14749 3485 14783 3519
rect 18153 3485 18187 3519
rect 18889 3485 18923 3519
rect 20177 3485 20211 3519
rect 22109 3485 22143 3519
rect 40417 3485 40451 3519
rect 48145 3485 48179 3519
rect 54677 3485 54711 3519
rect 55689 3485 55723 3519
rect 56333 3485 56367 3519
rect 56977 3485 57011 3519
rect 57437 3485 57471 3519
rect 58265 3485 58299 3519
rect 7757 3417 7791 3451
rect 17877 3417 17911 3451
rect 23949 3417 23983 3451
rect 1777 3349 1811 3383
rect 2605 3349 2639 3383
rect 2973 3349 3007 3383
rect 8585 3349 8619 3383
rect 15209 3349 15243 3383
rect 18705 3349 18739 3383
rect 20269 3349 20303 3383
rect 20637 3349 20671 3383
rect 21925 3349 21959 3383
rect 22569 3349 22603 3383
rect 22937 3349 22971 3383
rect 40233 3349 40267 3383
rect 47961 3349 47995 3383
rect 54493 3349 54527 3383
rect 55505 3349 55539 3383
rect 56149 3349 56183 3383
rect 56793 3349 56827 3383
rect 57621 3349 57655 3383
rect 58081 3349 58115 3383
rect 1777 3145 1811 3179
rect 2513 3145 2547 3179
rect 2973 3145 3007 3179
rect 12633 3145 12667 3179
rect 22201 3145 22235 3179
rect 23213 3145 23247 3179
rect 27261 3145 27295 3179
rect 28825 3145 28859 3179
rect 29929 3145 29963 3179
rect 30941 3145 30975 3179
rect 33241 3145 33275 3179
rect 43821 3145 43855 3179
rect 44833 3145 44867 3179
rect 45845 3145 45879 3179
rect 51457 3145 51491 3179
rect 53757 3145 53791 3179
rect 54769 3145 54803 3179
rect 56701 3145 56735 3179
rect 6745 3077 6779 3111
rect 14105 3077 14139 3111
rect 18337 3077 18371 3111
rect 32321 3077 32355 3111
rect 37933 3077 37967 3111
rect 2605 3009 2639 3043
rect 3433 3009 3467 3043
rect 6009 3009 6043 3043
rect 7021 3009 7055 3043
rect 9781 3009 9815 3043
rect 14381 3009 14415 3043
rect 18613 3009 18647 3043
rect 19349 3009 19383 3043
rect 20545 3009 20579 3043
rect 21373 3009 21407 3043
rect 22385 3009 22419 3043
rect 22845 3009 22879 3043
rect 23029 3009 23063 3043
rect 27813 3009 27847 3043
rect 54309 3009 54343 3043
rect 56057 3009 56091 3043
rect 56885 3009 56919 3043
rect 57529 3009 57563 3043
rect 58265 3009 58299 3043
rect 2421 2941 2455 2975
rect 4261 2941 4295 2975
rect 5733 2941 5767 2975
rect 9505 2941 9539 2975
rect 16313 2941 16347 2975
rect 19073 2941 19107 2975
rect 38669 2941 38703 2975
rect 8033 2873 8067 2907
rect 15761 2873 15795 2907
rect 16865 2873 16899 2907
rect 20361 2873 20395 2907
rect 21189 2873 21223 2907
rect 39405 2873 39439 2907
rect 58081 2873 58115 2907
rect 3617 2805 3651 2839
rect 7573 2805 7607 2839
rect 10241 2805 10275 2839
rect 11161 2805 11195 2839
rect 12081 2805 12115 2839
rect 15209 2805 15243 2839
rect 23673 2805 23707 2839
rect 24409 2805 24443 2839
rect 25513 2805 25547 2839
rect 27997 2805 28031 2839
rect 36001 2805 36035 2839
rect 50813 2805 50847 2839
rect 55597 2805 55631 2839
rect 56241 2805 56275 2839
rect 57345 2805 57379 2839
rect 2605 2601 2639 2635
rect 10977 2601 11011 2635
rect 22477 2601 22511 2635
rect 23397 2601 23431 2635
rect 24961 2601 24995 2635
rect 56701 2601 56735 2635
rect 1961 2533 1995 2567
rect 12541 2533 12575 2567
rect 15945 2533 15979 2567
rect 17141 2533 17175 2567
rect 6837 2465 6871 2499
rect 7941 2465 7975 2499
rect 14565 2465 14599 2499
rect 18153 2465 18187 2499
rect 20085 2465 20119 2499
rect 20361 2465 20395 2499
rect 27905 2465 27939 2499
rect 35541 2465 35575 2499
rect 2421 2397 2455 2431
rect 3433 2397 3467 2431
rect 4629 2397 4663 2431
rect 5733 2397 5767 2431
rect 7021 2397 7055 2431
rect 9229 2397 9263 2431
rect 12357 2397 12391 2431
rect 17877 2397 17911 2431
rect 22293 2397 22327 2431
rect 23581 2397 23615 2431
rect 26065 2397 26099 2431
rect 28917 2397 28951 2431
rect 30021 2397 30055 2431
rect 31125 2397 31159 2431
rect 32321 2397 32355 2431
rect 33333 2397 33367 2431
rect 34989 2397 35023 2431
rect 36093 2397 36127 2431
rect 37749 2397 37783 2431
rect 38485 2397 38519 2431
rect 39221 2397 39255 2431
rect 40325 2397 40359 2431
rect 41337 2397 41371 2431
rect 42901 2397 42935 2431
rect 43637 2397 43671 2431
rect 44649 2397 44683 2431
rect 45753 2397 45787 2431
rect 46869 2397 46903 2431
rect 48053 2397 48087 2431
rect 49065 2397 49099 2431
rect 49525 2397 49559 2431
rect 50629 2397 50663 2431
rect 51365 2397 51399 2431
rect 52377 2397 52411 2431
rect 53481 2397 53515 2431
rect 54585 2397 54619 2431
rect 55781 2397 55815 2431
rect 56517 2397 56551 2431
rect 57529 2397 57563 2431
rect 58081 2397 58115 2431
rect 4169 2329 4203 2363
rect 8125 2329 8159 2363
rect 10333 2329 10367 2363
rect 11069 2329 11103 2363
rect 11897 2329 11931 2363
rect 13645 2329 13679 2363
rect 14749 2329 14783 2363
rect 15761 2329 15795 2363
rect 16957 2329 16991 2363
rect 19625 2329 19659 2363
rect 24685 2329 24719 2363
rect 25697 2329 25731 2363
rect 27169 2329 27203 2363
rect 36369 2329 36403 2363
rect 4813 2261 4847 2295
rect 5917 2261 5951 2295
rect 9321 2261 9355 2295
rect 10241 2261 10275 2295
rect 13553 2261 13587 2295
rect 21373 2261 21407 2295
rect 26617 2261 26651 2295
rect 29101 2261 29135 2295
rect 30205 2261 30239 2295
rect 31309 2261 31343 2295
rect 32505 2261 32539 2295
rect 33517 2261 33551 2295
rect 34345 2261 34379 2295
rect 37565 2261 37599 2295
rect 38301 2261 38335 2295
rect 39037 2261 39071 2295
rect 40141 2261 40175 2295
rect 41153 2261 41187 2295
rect 41889 2261 41923 2295
rect 42717 2261 42751 2295
rect 43453 2261 43487 2295
rect 44465 2261 44499 2295
rect 45569 2261 45603 2295
rect 46673 2261 46707 2295
rect 47869 2261 47903 2295
rect 48881 2261 48915 2295
rect 50445 2261 50479 2295
rect 51181 2261 51215 2295
rect 52193 2261 52227 2295
rect 53297 2261 53331 2295
rect 54401 2261 54435 2295
rect 55597 2261 55631 2295
rect 57345 2261 57379 2295
rect 58265 2261 58299 2295
<< metal1 >>
rect 2222 57808 2228 57860
rect 2280 57848 2286 57860
rect 26234 57848 26240 57860
rect 2280 57820 26240 57848
rect 2280 57808 2286 57820
rect 26234 57808 26240 57820
rect 26292 57808 26298 57860
rect 21634 57740 21640 57792
rect 21692 57780 21698 57792
rect 30282 57780 30288 57792
rect 21692 57752 30288 57780
rect 21692 57740 21698 57752
rect 30282 57740 30288 57752
rect 30340 57740 30346 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 4525 57579 4583 57585
rect 4525 57545 4537 57579
rect 4571 57576 4583 57579
rect 17681 57579 17739 57585
rect 4571 57548 17632 57576
rect 4571 57545 4583 57548
rect 4525 57539 4583 57545
rect 11149 57511 11207 57517
rect 11149 57477 11161 57511
rect 11195 57508 11207 57511
rect 11422 57508 11428 57520
rect 11195 57480 11428 57508
rect 11195 57477 11207 57480
rect 11149 57471 11207 57477
rect 11422 57468 11428 57480
rect 11480 57468 11486 57520
rect 13725 57511 13783 57517
rect 13725 57477 13737 57511
rect 13771 57508 13783 57511
rect 13814 57508 13820 57520
rect 13771 57480 13820 57508
rect 13771 57477 13783 57480
rect 13725 57471 13783 57477
rect 13814 57468 13820 57480
rect 13872 57508 13878 57520
rect 16206 57508 16212 57520
rect 13872 57480 14320 57508
rect 16167 57480 16212 57508
rect 13872 57468 13878 57480
rect 1854 57400 1860 57452
rect 1912 57440 1918 57452
rect 1949 57443 2007 57449
rect 1949 57440 1961 57443
rect 1912 57412 1961 57440
rect 1912 57400 1918 57412
rect 1949 57409 1961 57412
rect 1995 57409 2007 57443
rect 2222 57440 2228 57452
rect 2183 57412 2228 57440
rect 1949 57403 2007 57409
rect 2222 57400 2228 57412
rect 2280 57400 2286 57452
rect 3050 57400 3056 57452
rect 3108 57440 3114 57452
rect 3237 57443 3295 57449
rect 3237 57440 3249 57443
rect 3108 57412 3249 57440
rect 3108 57400 3114 57412
rect 3237 57409 3249 57412
rect 3283 57409 3295 57443
rect 3237 57403 3295 57409
rect 4246 57400 4252 57452
rect 4304 57440 4310 57452
rect 4341 57443 4399 57449
rect 4341 57440 4353 57443
rect 4304 57412 4353 57440
rect 4304 57400 4310 57412
rect 4341 57409 4353 57412
rect 4387 57440 4399 57443
rect 4614 57440 4620 57452
rect 4387 57412 4620 57440
rect 4387 57409 4399 57412
rect 4341 57403 4399 57409
rect 4614 57400 4620 57412
rect 4672 57400 4678 57452
rect 5534 57400 5540 57452
rect 5592 57440 5598 57452
rect 5994 57440 6000 57452
rect 5592 57412 6000 57440
rect 5592 57400 5598 57412
rect 5994 57400 6000 57412
rect 6052 57400 6058 57452
rect 6638 57400 6644 57452
rect 6696 57440 6702 57452
rect 6733 57443 6791 57449
rect 6733 57440 6745 57443
rect 6696 57412 6745 57440
rect 6696 57400 6702 57412
rect 6733 57409 6745 57412
rect 6779 57409 6791 57443
rect 6733 57403 6791 57409
rect 7834 57400 7840 57452
rect 7892 57440 7898 57452
rect 8478 57440 8484 57452
rect 7892 57412 8484 57440
rect 7892 57400 7898 57412
rect 8478 57400 8484 57412
rect 8536 57440 8542 57452
rect 8573 57443 8631 57449
rect 8573 57440 8585 57443
rect 8536 57412 8585 57440
rect 8536 57400 8542 57412
rect 8573 57409 8585 57412
rect 8619 57409 8631 57443
rect 8573 57403 8631 57409
rect 9030 57400 9036 57452
rect 9088 57440 9094 57452
rect 9125 57443 9183 57449
rect 9125 57440 9137 57443
rect 9088 57412 9137 57440
rect 9088 57400 9094 57412
rect 9125 57409 9137 57412
rect 9171 57409 9183 57443
rect 9125 57403 9183 57409
rect 9861 57443 9919 57449
rect 9861 57409 9873 57443
rect 9907 57440 9919 57443
rect 10226 57440 10232 57452
rect 9907 57412 10232 57440
rect 9907 57409 9919 57412
rect 9861 57403 9919 57409
rect 10226 57400 10232 57412
rect 10284 57440 10290 57452
rect 10321 57443 10379 57449
rect 10321 57440 10333 57443
rect 10284 57412 10333 57440
rect 10284 57400 10290 57412
rect 10321 57409 10333 57412
rect 10367 57409 10379 57443
rect 11440 57440 11468 57468
rect 11701 57443 11759 57449
rect 11701 57440 11713 57443
rect 11440 57412 11713 57440
rect 10321 57403 10379 57409
rect 11701 57409 11713 57412
rect 11747 57409 11759 57443
rect 11701 57403 11759 57409
rect 12618 57400 12624 57452
rect 12676 57440 12682 57452
rect 14292 57449 14320 57480
rect 16206 57468 16212 57480
rect 16264 57508 16270 57520
rect 17604 57508 17632 57548
rect 17681 57545 17693 57579
rect 17727 57576 17739 57579
rect 22002 57576 22008 57588
rect 17727 57548 22008 57576
rect 17727 57545 17739 57548
rect 17681 57539 17739 57545
rect 22002 57536 22008 57548
rect 22060 57536 22066 57588
rect 25409 57579 25467 57585
rect 25409 57545 25421 57579
rect 25455 57576 25467 57579
rect 25774 57576 25780 57588
rect 25455 57548 25780 57576
rect 25455 57545 25467 57548
rect 25409 57539 25467 57545
rect 25774 57536 25780 57548
rect 25832 57536 25838 57588
rect 26605 57579 26663 57585
rect 26605 57545 26617 57579
rect 26651 57576 26663 57579
rect 26970 57576 26976 57588
rect 26651 57548 26976 57576
rect 26651 57545 26663 57548
rect 26605 57539 26663 57545
rect 26970 57536 26976 57548
rect 27028 57536 27034 57588
rect 29181 57579 29239 57585
rect 29181 57545 29193 57579
rect 29227 57576 29239 57579
rect 29362 57576 29368 57588
rect 29227 57548 29368 57576
rect 29227 57545 29239 57548
rect 29181 57539 29239 57545
rect 29362 57536 29368 57548
rect 29420 57536 29426 57588
rect 34146 57536 34152 57588
rect 34204 57576 34210 57588
rect 34241 57579 34299 57585
rect 34241 57576 34253 57579
rect 34204 57548 34253 57576
rect 34204 57536 34210 57548
rect 34241 57545 34253 57548
rect 34287 57545 34299 57579
rect 34241 57539 34299 57545
rect 21910 57508 21916 57520
rect 16264 57480 16574 57508
rect 17604 57480 21916 57508
rect 16264 57468 16270 57480
rect 12713 57443 12771 57449
rect 12713 57440 12725 57443
rect 12676 57412 12725 57440
rect 12676 57400 12682 57412
rect 12713 57409 12725 57412
rect 12759 57409 12771 57443
rect 12713 57403 12771 57409
rect 14277 57443 14335 57449
rect 14277 57409 14289 57443
rect 14323 57409 14335 57443
rect 14277 57403 14335 57409
rect 15010 57400 15016 57452
rect 15068 57440 15074 57452
rect 15105 57443 15163 57449
rect 15105 57440 15117 57443
rect 15068 57412 15117 57440
rect 15068 57400 15074 57412
rect 15105 57409 15117 57412
rect 15151 57409 15163 57443
rect 16546 57440 16574 57480
rect 21910 57468 21916 57480
rect 21968 57468 21974 57520
rect 16853 57443 16911 57449
rect 16853 57440 16865 57443
rect 16546 57412 16865 57440
rect 15105 57403 15163 57409
rect 16853 57409 16865 57412
rect 16899 57409 16911 57443
rect 16853 57403 16911 57409
rect 17402 57400 17408 57452
rect 17460 57440 17466 57452
rect 17497 57443 17555 57449
rect 17497 57440 17509 57443
rect 17460 57412 17509 57440
rect 17460 57400 17466 57412
rect 17497 57409 17509 57412
rect 17543 57409 17555 57443
rect 17497 57403 17555 57409
rect 18233 57443 18291 57449
rect 18233 57409 18245 57443
rect 18279 57440 18291 57443
rect 18598 57440 18604 57452
rect 18279 57412 18604 57440
rect 18279 57409 18291 57412
rect 18233 57403 18291 57409
rect 18598 57400 18604 57412
rect 18656 57440 18662 57452
rect 18693 57443 18751 57449
rect 18693 57440 18705 57443
rect 18656 57412 18705 57440
rect 18656 57400 18662 57412
rect 18693 57409 18705 57412
rect 18739 57409 18751 57443
rect 18693 57403 18751 57409
rect 19889 57443 19947 57449
rect 19889 57409 19901 57443
rect 19935 57440 19947 57443
rect 19978 57440 19984 57452
rect 19935 57412 19984 57440
rect 19935 57409 19947 57412
rect 19889 57403 19947 57409
rect 19978 57400 19984 57412
rect 20036 57400 20042 57452
rect 20625 57443 20683 57449
rect 20625 57409 20637 57443
rect 20671 57440 20683 57443
rect 20990 57440 20996 57452
rect 20671 57412 20996 57440
rect 20671 57409 20683 57412
rect 20625 57403 20683 57409
rect 20990 57400 20996 57412
rect 21048 57440 21054 57452
rect 21085 57443 21143 57449
rect 21085 57440 21097 57443
rect 21048 57412 21097 57440
rect 21048 57400 21054 57412
rect 21085 57409 21097 57412
rect 21131 57409 21143 57443
rect 21085 57403 21143 57409
rect 22186 57400 22192 57452
rect 22244 57440 22250 57452
rect 22281 57443 22339 57449
rect 22281 57440 22293 57443
rect 22244 57412 22293 57440
rect 22244 57400 22250 57412
rect 22281 57409 22293 57412
rect 22327 57409 22339 57443
rect 22281 57403 22339 57409
rect 23017 57443 23075 57449
rect 23017 57409 23029 57443
rect 23063 57440 23075 57443
rect 23382 57440 23388 57452
rect 23063 57412 23388 57440
rect 23063 57409 23075 57412
rect 23017 57403 23075 57409
rect 23382 57400 23388 57412
rect 23440 57440 23446 57452
rect 23477 57443 23535 57449
rect 23477 57440 23489 57443
rect 23440 57412 23489 57440
rect 23440 57400 23446 57412
rect 23477 57409 23489 57412
rect 23523 57409 23535 57443
rect 23477 57403 23535 57409
rect 24578 57400 24584 57452
rect 24636 57440 24642 57452
rect 24673 57443 24731 57449
rect 24673 57440 24685 57443
rect 24636 57412 24685 57440
rect 24636 57400 24642 57412
rect 24673 57409 24685 57412
rect 24719 57409 24731 57443
rect 25792 57440 25820 57536
rect 26053 57443 26111 57449
rect 26053 57440 26065 57443
rect 25792 57412 26065 57440
rect 24673 57403 24731 57409
rect 26053 57409 26065 57412
rect 26099 57409 26111 57443
rect 26988 57440 27016 57536
rect 27341 57443 27399 57449
rect 27341 57440 27353 57443
rect 26988 57412 27353 57440
rect 26053 57403 26111 57409
rect 27341 57409 27353 57412
rect 27387 57409 27399 57443
rect 27341 57403 27399 57409
rect 28166 57400 28172 57452
rect 28224 57440 28230 57452
rect 28261 57443 28319 57449
rect 28261 57440 28273 57443
rect 28224 57412 28273 57440
rect 28224 57400 28230 57412
rect 28261 57409 28273 57412
rect 28307 57409 28319 57443
rect 29380 57440 29408 57536
rect 29917 57443 29975 57449
rect 29917 57440 29929 57443
rect 29380 57412 29929 57440
rect 28261 57403 28319 57409
rect 29917 57409 29929 57412
rect 29963 57409 29975 57443
rect 29917 57403 29975 57409
rect 30558 57400 30564 57452
rect 30616 57440 30622 57452
rect 30653 57443 30711 57449
rect 30653 57440 30665 57443
rect 30616 57412 30665 57440
rect 30616 57400 30622 57412
rect 30653 57409 30665 57412
rect 30699 57440 30711 57443
rect 31297 57443 31355 57449
rect 31297 57440 31309 57443
rect 30699 57412 31309 57440
rect 30699 57409 30711 57412
rect 30653 57403 30711 57409
rect 31297 57409 31309 57412
rect 31343 57409 31355 57443
rect 31297 57403 31355 57409
rect 31754 57400 31760 57452
rect 31812 57440 31818 57452
rect 32122 57440 32128 57452
rect 31812 57412 32128 57440
rect 31812 57400 31818 57412
rect 32122 57400 32128 57412
rect 32180 57440 32186 57452
rect 32309 57443 32367 57449
rect 32309 57440 32321 57443
rect 32180 57412 32321 57440
rect 32180 57400 32186 57412
rect 32309 57409 32321 57412
rect 32355 57409 32367 57443
rect 32309 57403 32367 57409
rect 32950 57400 32956 57452
rect 33008 57440 33014 57452
rect 33045 57443 33103 57449
rect 33045 57440 33057 57443
rect 33008 57412 33057 57440
rect 33008 57400 33014 57412
rect 33045 57409 33057 57412
rect 33091 57440 33103 57443
rect 33689 57443 33747 57449
rect 33689 57440 33701 57443
rect 33091 57412 33701 57440
rect 33091 57409 33103 57412
rect 33045 57403 33103 57409
rect 33689 57409 33701 57412
rect 33735 57409 33747 57443
rect 34256 57440 34284 57539
rect 45462 57536 45468 57588
rect 45520 57576 45526 57588
rect 47765 57579 47823 57585
rect 47765 57576 47777 57579
rect 45520 57548 47777 57576
rect 45520 57536 45526 57548
rect 47765 57545 47777 57548
rect 47811 57545 47823 57579
rect 47765 57539 47823 57545
rect 50341 57579 50399 57585
rect 50341 57545 50353 57579
rect 50387 57545 50399 57579
rect 50341 57539 50399 57545
rect 42886 57468 42892 57520
rect 42944 57508 42950 57520
rect 50356 57508 50384 57539
rect 50430 57536 50436 57588
rect 50488 57576 50494 57588
rect 50488 57548 55214 57576
rect 50488 57536 50494 57548
rect 42944 57480 50384 57508
rect 42944 57468 42950 57480
rect 34885 57443 34943 57449
rect 34885 57440 34897 57443
rect 34256 57412 34897 57440
rect 33689 57403 33747 57409
rect 34885 57409 34897 57412
rect 34931 57409 34943 57443
rect 34885 57403 34943 57409
rect 35342 57400 35348 57452
rect 35400 57440 35406 57452
rect 35713 57443 35771 57449
rect 35713 57440 35725 57443
rect 35400 57412 35725 57440
rect 35400 57400 35406 57412
rect 35713 57409 35725 57412
rect 35759 57409 35771 57443
rect 35713 57403 35771 57409
rect 36538 57400 36544 57452
rect 36596 57440 36602 57452
rect 36817 57443 36875 57449
rect 36817 57440 36829 57443
rect 36596 57412 36829 57440
rect 36596 57400 36602 57412
rect 36817 57409 36829 57412
rect 36863 57409 36875 57443
rect 36817 57403 36875 57409
rect 37734 57400 37740 57452
rect 37792 57440 37798 57452
rect 38013 57443 38071 57449
rect 38013 57440 38025 57443
rect 37792 57412 38025 57440
rect 37792 57400 37798 57412
rect 38013 57409 38025 57412
rect 38059 57440 38071 57443
rect 38473 57443 38531 57449
rect 38473 57440 38485 57443
rect 38059 57412 38485 57440
rect 38059 57409 38071 57412
rect 38013 57403 38071 57409
rect 38473 57409 38485 57412
rect 38519 57409 38531 57443
rect 38473 57403 38531 57409
rect 38930 57400 38936 57452
rect 38988 57440 38994 57452
rect 39209 57443 39267 57449
rect 39209 57440 39221 57443
rect 38988 57412 39221 57440
rect 38988 57400 38994 57412
rect 39209 57409 39221 57412
rect 39255 57409 39267 57443
rect 39209 57403 39267 57409
rect 40126 57400 40132 57452
rect 40184 57440 40190 57452
rect 40405 57443 40463 57449
rect 40405 57440 40417 57443
rect 40184 57412 40417 57440
rect 40184 57400 40190 57412
rect 40405 57409 40417 57412
rect 40451 57440 40463 57443
rect 40865 57443 40923 57449
rect 40865 57440 40877 57443
rect 40451 57412 40877 57440
rect 40451 57409 40463 57412
rect 40405 57403 40463 57409
rect 40865 57409 40877 57412
rect 40911 57409 40923 57443
rect 40865 57403 40923 57409
rect 41322 57400 41328 57452
rect 41380 57440 41386 57452
rect 41601 57443 41659 57449
rect 41601 57440 41613 57443
rect 41380 57412 41613 57440
rect 41380 57400 41386 57412
rect 41601 57409 41613 57412
rect 41647 57409 41659 57443
rect 42794 57440 42800 57452
rect 42755 57412 42800 57440
rect 41601 57403 41659 57409
rect 42794 57400 42800 57412
rect 42852 57440 42858 57452
rect 43257 57443 43315 57449
rect 43257 57440 43269 57443
rect 42852 57412 43269 57440
rect 42852 57400 42858 57412
rect 43257 57409 43269 57412
rect 43303 57409 43315 57443
rect 43257 57403 43315 57409
rect 43714 57400 43720 57452
rect 43772 57440 43778 57452
rect 43993 57443 44051 57449
rect 43993 57440 44005 57443
rect 43772 57412 44005 57440
rect 43772 57400 43778 57412
rect 43993 57409 44005 57412
rect 44039 57440 44051 57443
rect 44453 57443 44511 57449
rect 44453 57440 44465 57443
rect 44039 57412 44465 57440
rect 44039 57409 44051 57412
rect 43993 57403 44051 57409
rect 44453 57409 44465 57412
rect 44499 57409 44511 57443
rect 44453 57403 44511 57409
rect 44910 57400 44916 57452
rect 44968 57440 44974 57452
rect 45373 57443 45431 57449
rect 45373 57440 45385 57443
rect 44968 57412 45385 57440
rect 44968 57400 44974 57412
rect 45373 57409 45385 57412
rect 45419 57409 45431 57443
rect 45373 57403 45431 57409
rect 46106 57400 46112 57452
rect 46164 57440 46170 57452
rect 46385 57443 46443 57449
rect 46385 57440 46397 57443
rect 46164 57412 46397 57440
rect 46164 57400 46170 57412
rect 46385 57409 46397 57412
rect 46431 57440 46443 57443
rect 46845 57443 46903 57449
rect 46845 57440 46857 57443
rect 46431 57412 46857 57440
rect 46431 57409 46443 57412
rect 46385 57403 46443 57409
rect 46845 57409 46857 57412
rect 46891 57409 46903 57443
rect 46845 57403 46903 57409
rect 47302 57400 47308 57452
rect 47360 57440 47366 57452
rect 47949 57443 48007 57449
rect 47949 57440 47961 57443
rect 47360 57412 47961 57440
rect 47360 57400 47366 57412
rect 47949 57409 47961 57412
rect 47995 57409 48007 57443
rect 47949 57403 48007 57409
rect 48498 57400 48504 57452
rect 48556 57440 48562 57452
rect 48777 57443 48835 57449
rect 48777 57440 48789 57443
rect 48556 57412 48789 57440
rect 48556 57400 48562 57412
rect 48777 57409 48789 57412
rect 48823 57440 48835 57443
rect 49237 57443 49295 57449
rect 49237 57440 49249 57443
rect 48823 57412 49249 57440
rect 48823 57409 48835 57412
rect 48777 57403 48835 57409
rect 49237 57409 49249 57412
rect 49283 57409 49295 57443
rect 49237 57403 49295 57409
rect 49694 57400 49700 57452
rect 49752 57440 49758 57452
rect 50338 57440 50344 57452
rect 49752 57412 50344 57440
rect 49752 57400 49758 57412
rect 50338 57400 50344 57412
rect 50396 57440 50402 57452
rect 50525 57443 50583 57449
rect 50525 57440 50537 57443
rect 50396 57412 50537 57440
rect 50396 57400 50402 57412
rect 50525 57409 50537 57412
rect 50571 57409 50583 57443
rect 50525 57403 50583 57409
rect 51074 57400 51080 57452
rect 51132 57440 51138 57452
rect 51169 57443 51227 57449
rect 51169 57440 51181 57443
rect 51132 57412 51181 57440
rect 51132 57400 51138 57412
rect 51169 57409 51181 57412
rect 51215 57440 51227 57443
rect 51629 57443 51687 57449
rect 51629 57440 51641 57443
rect 51215 57412 51641 57440
rect 51215 57409 51227 57412
rect 51169 57403 51227 57409
rect 51629 57409 51641 57412
rect 51675 57409 51687 57443
rect 51629 57403 51687 57409
rect 52086 57400 52092 57452
rect 52144 57440 52150 57452
rect 52365 57443 52423 57449
rect 52365 57440 52377 57443
rect 52144 57412 52377 57440
rect 52144 57400 52150 57412
rect 52365 57409 52377 57412
rect 52411 57409 52423 57443
rect 52365 57403 52423 57409
rect 53282 57400 53288 57452
rect 53340 57440 53346 57452
rect 53561 57443 53619 57449
rect 53561 57440 53573 57443
rect 53340 57412 53573 57440
rect 53340 57400 53346 57412
rect 53561 57409 53573 57412
rect 53607 57440 53619 57443
rect 54021 57443 54079 57449
rect 54021 57440 54033 57443
rect 53607 57412 54033 57440
rect 53607 57409 53619 57412
rect 53561 57403 53619 57409
rect 54021 57409 54033 57412
rect 54067 57409 54079 57443
rect 54021 57403 54079 57409
rect 54478 57400 54484 57452
rect 54536 57440 54542 57452
rect 54757 57443 54815 57449
rect 54757 57440 54769 57443
rect 54536 57412 54769 57440
rect 54536 57400 54542 57412
rect 54757 57409 54769 57412
rect 54803 57409 54815 57443
rect 54757 57403 54815 57409
rect 5718 57372 5724 57384
rect 5679 57344 5724 57372
rect 5718 57332 5724 57344
rect 5776 57332 5782 57384
rect 8294 57372 8300 57384
rect 8255 57344 8300 57372
rect 8294 57332 8300 57344
rect 8352 57332 8358 57384
rect 18966 57372 18972 57384
rect 14476 57344 18972 57372
rect 14476 57313 14504 57344
rect 18966 57332 18972 57344
rect 19024 57332 19030 57384
rect 28626 57372 28632 57384
rect 21284 57344 28632 57372
rect 10505 57307 10563 57313
rect 10505 57273 10517 57307
rect 10551 57304 10563 57307
rect 14461 57307 14519 57313
rect 10551 57276 14412 57304
rect 10551 57273 10563 57276
rect 10505 57267 10563 57273
rect 3418 57236 3424 57248
rect 3379 57208 3424 57236
rect 3418 57196 3424 57208
rect 3476 57196 3482 57248
rect 6914 57196 6920 57248
rect 6972 57236 6978 57248
rect 9306 57236 9312 57248
rect 6972 57208 7017 57236
rect 9267 57208 9312 57236
rect 6972 57196 6978 57208
rect 9306 57196 9312 57208
rect 9364 57196 9370 57248
rect 11882 57236 11888 57248
rect 11843 57208 11888 57236
rect 11882 57196 11888 57208
rect 11940 57196 11946 57248
rect 12894 57236 12900 57248
rect 12855 57208 12900 57236
rect 12894 57196 12900 57208
rect 12952 57196 12958 57248
rect 14384 57236 14412 57276
rect 14461 57273 14473 57307
rect 14507 57273 14519 57307
rect 14461 57267 14519 57273
rect 15289 57307 15347 57313
rect 15289 57273 15301 57307
rect 15335 57304 15347 57307
rect 20806 57304 20812 57316
rect 15335 57276 20812 57304
rect 15335 57273 15347 57276
rect 15289 57267 15347 57273
rect 20806 57264 20812 57276
rect 20864 57264 20870 57316
rect 21284 57313 21312 57344
rect 28626 57332 28632 57344
rect 28684 57332 28690 57384
rect 40034 57332 40040 57384
rect 40092 57372 40098 57384
rect 40092 57344 43852 57372
rect 40092 57332 40098 57344
rect 21269 57307 21327 57313
rect 21269 57273 21281 57307
rect 21315 57273 21327 57307
rect 21269 57267 21327 57273
rect 23661 57307 23719 57313
rect 23661 57273 23673 57307
rect 23707 57304 23719 57307
rect 25038 57304 25044 57316
rect 23707 57276 25044 57304
rect 23707 57273 23719 57276
rect 23661 57267 23719 57273
rect 25038 57264 25044 57276
rect 25096 57264 25102 57316
rect 30837 57307 30895 57313
rect 30837 57273 30849 57307
rect 30883 57304 30895 57307
rect 33134 57304 33140 57316
rect 30883 57276 33140 57304
rect 30883 57273 30895 57276
rect 30837 57267 30895 57273
rect 33134 57264 33140 57276
rect 33192 57264 33198 57316
rect 37642 57264 37648 57316
rect 37700 57304 37706 57316
rect 40221 57307 40279 57313
rect 40221 57304 40233 57307
rect 37700 57276 40233 57304
rect 37700 57264 37706 57276
rect 40221 57273 40233 57276
rect 40267 57273 40279 57307
rect 40221 57267 40279 57273
rect 40494 57264 40500 57316
rect 40552 57304 40558 57316
rect 43824 57313 43852 57344
rect 44266 57332 44272 57384
rect 44324 57372 44330 57384
rect 44324 57344 51028 57372
rect 44324 57332 44330 57344
rect 42613 57307 42671 57313
rect 42613 57304 42625 57307
rect 40552 57276 42625 57304
rect 40552 57264 40558 57276
rect 42613 57273 42625 57276
rect 42659 57273 42671 57307
rect 42613 57267 42671 57273
rect 43809 57307 43867 57313
rect 43809 57273 43821 57307
rect 43855 57273 43867 57307
rect 43809 57267 43867 57273
rect 44174 57264 44180 57316
rect 44232 57304 44238 57316
rect 51000 57313 51028 57344
rect 48593 57307 48651 57313
rect 48593 57304 48605 57307
rect 44232 57276 48605 57304
rect 44232 57264 44238 57276
rect 48593 57273 48605 57276
rect 48639 57273 48651 57307
rect 48593 57267 48651 57273
rect 50985 57307 51043 57313
rect 50985 57273 50997 57307
rect 51031 57273 51043 57307
rect 55186 57304 55214 57548
rect 55674 57400 55680 57452
rect 55732 57440 55738 57452
rect 55953 57443 56011 57449
rect 55953 57440 55965 57443
rect 55732 57412 55965 57440
rect 55732 57400 55738 57412
rect 55953 57409 55965 57412
rect 55999 57440 56011 57443
rect 56413 57443 56471 57449
rect 56413 57440 56425 57443
rect 55999 57412 56425 57440
rect 55999 57409 56011 57412
rect 55953 57403 56011 57409
rect 56413 57409 56425 57412
rect 56459 57409 56471 57443
rect 56413 57403 56471 57409
rect 56870 57400 56876 57452
rect 56928 57440 56934 57452
rect 57149 57443 57207 57449
rect 57149 57440 57161 57443
rect 56928 57412 57161 57440
rect 56928 57400 56934 57412
rect 57149 57409 57161 57412
rect 57195 57409 57207 57443
rect 57149 57403 57207 57409
rect 58066 57400 58072 57452
rect 58124 57440 58130 57452
rect 58345 57443 58403 57449
rect 58345 57440 58357 57443
rect 58124 57412 58357 57440
rect 58124 57400 58130 57412
rect 58345 57409 58357 57412
rect 58391 57409 58403 57443
rect 58345 57403 58403 57409
rect 56965 57307 57023 57313
rect 56965 57304 56977 57307
rect 55186 57276 56977 57304
rect 50985 57267 51043 57273
rect 56965 57273 56977 57276
rect 57011 57273 57023 57307
rect 56965 57267 57023 57273
rect 16298 57236 16304 57248
rect 14384 57208 16304 57236
rect 16298 57196 16304 57208
rect 16356 57196 16362 57248
rect 17034 57236 17040 57248
rect 16995 57208 17040 57236
rect 17034 57196 17040 57208
rect 17092 57196 17098 57248
rect 18874 57236 18880 57248
rect 18835 57208 18880 57236
rect 18874 57196 18880 57208
rect 18932 57196 18938 57248
rect 20073 57239 20131 57245
rect 20073 57205 20085 57239
rect 20119 57236 20131 57239
rect 22278 57236 22284 57248
rect 20119 57208 22284 57236
rect 20119 57205 20131 57208
rect 20073 57199 20131 57205
rect 22278 57196 22284 57208
rect 22336 57196 22342 57248
rect 22462 57236 22468 57248
rect 22423 57208 22468 57236
rect 22462 57196 22468 57208
rect 22520 57196 22526 57248
rect 24854 57236 24860 57248
rect 24815 57208 24860 57236
rect 24854 57196 24860 57208
rect 24912 57196 24918 57248
rect 25130 57196 25136 57248
rect 25188 57236 25194 57248
rect 25869 57239 25927 57245
rect 25869 57236 25881 57239
rect 25188 57208 25881 57236
rect 25188 57196 25194 57208
rect 25869 57205 25881 57208
rect 25915 57205 25927 57239
rect 27154 57236 27160 57248
rect 27115 57208 27160 57236
rect 25869 57199 25927 57205
rect 27154 57196 27160 57208
rect 27212 57196 27218 57248
rect 28445 57239 28503 57245
rect 28445 57205 28457 57239
rect 28491 57236 28503 57239
rect 28534 57236 28540 57248
rect 28491 57208 28540 57236
rect 28491 57205 28503 57208
rect 28445 57199 28503 57205
rect 28534 57196 28540 57208
rect 28592 57196 28598 57248
rect 29730 57236 29736 57248
rect 29691 57208 29736 57236
rect 29730 57196 29736 57208
rect 29788 57196 29794 57248
rect 32490 57236 32496 57248
rect 32451 57208 32496 57236
rect 32490 57196 32496 57208
rect 32548 57196 32554 57248
rect 33226 57236 33232 57248
rect 33187 57208 33232 57236
rect 33226 57196 33232 57208
rect 33284 57196 33290 57248
rect 34790 57196 34796 57248
rect 34848 57236 34854 57248
rect 35069 57239 35127 57245
rect 35069 57236 35081 57239
rect 34848 57208 35081 57236
rect 34848 57196 34854 57208
rect 35069 57205 35081 57208
rect 35115 57205 35127 57239
rect 35069 57199 35127 57205
rect 35434 57196 35440 57248
rect 35492 57236 35498 57248
rect 35529 57239 35587 57245
rect 35529 57236 35541 57239
rect 35492 57208 35541 57236
rect 35492 57196 35498 57208
rect 35529 57205 35541 57208
rect 35575 57205 35587 57239
rect 35529 57199 35587 57205
rect 36538 57196 36544 57248
rect 36596 57236 36602 57248
rect 36633 57239 36691 57245
rect 36633 57236 36645 57239
rect 36596 57208 36645 57236
rect 36596 57196 36602 57208
rect 36633 57205 36645 57208
rect 36679 57205 36691 57239
rect 36633 57199 36691 57205
rect 37182 57196 37188 57248
rect 37240 57236 37246 57248
rect 37829 57239 37887 57245
rect 37829 57236 37841 57239
rect 37240 57208 37841 57236
rect 37240 57196 37246 57208
rect 37829 57205 37841 57208
rect 37875 57205 37887 57239
rect 39022 57236 39028 57248
rect 38983 57208 39028 57236
rect 37829 57199 37887 57205
rect 39022 57196 39028 57208
rect 39080 57196 39086 57248
rect 41414 57196 41420 57248
rect 41472 57236 41478 57248
rect 41472 57208 41517 57236
rect 41472 57196 41478 57208
rect 42794 57196 42800 57248
rect 42852 57236 42858 57248
rect 45189 57239 45247 57245
rect 45189 57236 45201 57239
rect 42852 57208 45201 57236
rect 42852 57196 42858 57208
rect 45189 57205 45201 57208
rect 45235 57205 45247 57239
rect 46198 57236 46204 57248
rect 46159 57208 46204 57236
rect 45189 57199 45247 57205
rect 46198 57196 46204 57208
rect 46256 57196 46262 57248
rect 52178 57236 52184 57248
rect 52139 57208 52184 57236
rect 52178 57196 52184 57208
rect 52236 57196 52242 57248
rect 53374 57236 53380 57248
rect 53335 57208 53380 57236
rect 53374 57196 53380 57208
rect 53432 57196 53438 57248
rect 54570 57236 54576 57248
rect 54531 57208 54576 57236
rect 54570 57196 54576 57208
rect 54628 57196 54634 57248
rect 54662 57196 54668 57248
rect 54720 57236 54726 57248
rect 55769 57239 55827 57245
rect 55769 57236 55781 57239
rect 54720 57208 55781 57236
rect 54720 57196 54726 57208
rect 55769 57205 55781 57208
rect 55815 57205 55827 57239
rect 58158 57236 58164 57248
rect 58119 57208 58164 57236
rect 55769 57199 55827 57205
rect 58158 57196 58164 57208
rect 58216 57196 58222 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 1854 57032 1860 57044
rect 1815 57004 1860 57032
rect 1854 56992 1860 57004
rect 1912 56992 1918 57044
rect 3050 57032 3056 57044
rect 3011 57004 3056 57032
rect 3050 56992 3056 57004
rect 3108 56992 3114 57044
rect 4249 57035 4307 57041
rect 4249 57001 4261 57035
rect 4295 57032 4307 57035
rect 4614 57032 4620 57044
rect 4295 57004 4620 57032
rect 4295 57001 4307 57004
rect 4249 56995 4307 57001
rect 4614 56992 4620 57004
rect 4672 56992 4678 57044
rect 5994 57032 6000 57044
rect 5955 57004 6000 57032
rect 5994 56992 6000 57004
rect 6052 56992 6058 57044
rect 6638 57032 6644 57044
rect 6599 57004 6644 57032
rect 6638 56992 6644 57004
rect 6696 56992 6702 57044
rect 8478 57032 8484 57044
rect 8439 57004 8484 57032
rect 8478 56992 8484 57004
rect 8536 56992 8542 57044
rect 9030 56992 9036 57044
rect 9088 57032 9094 57044
rect 9125 57035 9183 57041
rect 9125 57032 9137 57035
rect 9088 57004 9137 57032
rect 9088 56992 9094 57004
rect 9125 57001 9137 57004
rect 9171 57001 9183 57035
rect 12618 57032 12624 57044
rect 12579 57004 12624 57032
rect 9125 56995 9183 57001
rect 12618 56992 12624 57004
rect 12676 56992 12682 57044
rect 15010 57032 15016 57044
rect 14971 57004 15016 57032
rect 15010 56992 15016 57004
rect 15068 56992 15074 57044
rect 16298 56992 16304 57044
rect 16356 57032 16362 57044
rect 19797 57035 19855 57041
rect 16356 57004 19380 57032
rect 16356 56992 16362 57004
rect 9306 56924 9312 56976
rect 9364 56964 9370 56976
rect 17862 56964 17868 56976
rect 9364 56936 17868 56964
rect 9364 56924 9370 56936
rect 17862 56924 17868 56936
rect 17920 56924 17926 56976
rect 19352 56964 19380 57004
rect 19797 57001 19809 57035
rect 19843 57032 19855 57035
rect 19978 57032 19984 57044
rect 19843 57004 19984 57032
rect 19843 57001 19855 57004
rect 19797 56995 19855 57001
rect 19978 56992 19984 57004
rect 20036 56992 20042 57044
rect 21634 57032 21640 57044
rect 21595 57004 21640 57032
rect 21634 56992 21640 57004
rect 21692 56992 21698 57044
rect 22186 57032 22192 57044
rect 22147 57004 22192 57032
rect 22186 56992 22192 57004
rect 22244 56992 22250 57044
rect 24578 57032 24584 57044
rect 24539 57004 24584 57032
rect 24578 56992 24584 57004
rect 24636 56992 24642 57044
rect 25869 57035 25927 57041
rect 25869 57001 25881 57035
rect 25915 57032 25927 57035
rect 26234 57032 26240 57044
rect 25915 57004 26240 57032
rect 25915 57001 25927 57004
rect 25869 56995 25927 57001
rect 26234 56992 26240 57004
rect 26292 56992 26298 57044
rect 28166 57032 28172 57044
rect 28127 57004 28172 57032
rect 28166 56992 28172 57004
rect 28224 56992 28230 57044
rect 32122 57032 32128 57044
rect 32083 57004 32128 57032
rect 32122 56992 32128 57004
rect 32180 56992 32186 57044
rect 35342 57032 35348 57044
rect 35303 57004 35348 57032
rect 35342 56992 35348 57004
rect 35400 56992 35406 57044
rect 36446 57032 36452 57044
rect 36407 57004 36452 57032
rect 36446 56992 36452 57004
rect 36504 56992 36510 57044
rect 38289 57035 38347 57041
rect 38289 57001 38301 57035
rect 38335 57032 38347 57035
rect 38930 57032 38936 57044
rect 38335 57004 38936 57032
rect 38335 57001 38347 57004
rect 38289 56995 38347 57001
rect 38930 56992 38936 57004
rect 38988 56992 38994 57044
rect 41322 57032 41328 57044
rect 41283 57004 41328 57032
rect 41322 56992 41328 57004
rect 41380 56992 41386 57044
rect 44910 56992 44916 57044
rect 44968 57032 44974 57044
rect 45189 57035 45247 57041
rect 45189 57032 45201 57035
rect 44968 57004 45201 57032
rect 44968 56992 44974 57004
rect 45189 57001 45201 57004
rect 45235 57001 45247 57035
rect 45189 56995 45247 57001
rect 47302 56992 47308 57044
rect 47360 57032 47366 57044
rect 47581 57035 47639 57041
rect 47581 57032 47593 57035
rect 47360 57004 47593 57032
rect 47360 56992 47366 57004
rect 47581 57001 47593 57004
rect 47627 57001 47639 57035
rect 50338 57032 50344 57044
rect 50299 57004 50344 57032
rect 47581 56995 47639 57001
rect 50338 56992 50344 57004
rect 50396 56992 50402 57044
rect 52086 57032 52092 57044
rect 52047 57004 52092 57032
rect 52086 56992 52092 57004
rect 52144 56992 52150 57044
rect 54478 57032 54484 57044
rect 54439 57004 54484 57032
rect 54478 56992 54484 57004
rect 54536 56992 54542 57044
rect 56413 57035 56471 57041
rect 56413 57001 56425 57035
rect 56459 57032 56471 57035
rect 56870 57032 56876 57044
rect 56459 57004 56876 57032
rect 56459 57001 56471 57004
rect 56413 56995 56471 57001
rect 56870 56992 56876 57004
rect 56928 56992 56934 57044
rect 22094 56964 22100 56976
rect 19352 56936 22100 56964
rect 22094 56924 22100 56936
rect 22152 56924 22158 56976
rect 22462 56924 22468 56976
rect 22520 56964 22526 56976
rect 28902 56964 28908 56976
rect 22520 56936 28908 56964
rect 22520 56924 22526 56936
rect 28902 56924 28908 56936
rect 28960 56924 28966 56976
rect 42702 56924 42708 56976
rect 42760 56964 42766 56976
rect 50430 56964 50436 56976
rect 42760 56936 50436 56964
rect 42760 56924 42766 56936
rect 50430 56924 50436 56936
rect 50488 56924 50494 56976
rect 11882 56856 11888 56908
rect 11940 56896 11946 56908
rect 20438 56896 20444 56908
rect 11940 56868 20444 56896
rect 11940 56856 11946 56868
rect 20438 56856 20444 56868
rect 20496 56856 20502 56908
rect 22278 56856 22284 56908
rect 22336 56896 22342 56908
rect 26418 56896 26424 56908
rect 22336 56868 26424 56896
rect 22336 56856 22342 56868
rect 26418 56856 26424 56868
rect 26476 56856 26482 56908
rect 29730 56896 29736 56908
rect 29691 56868 29736 56896
rect 29730 56856 29736 56868
rect 29788 56856 29794 56908
rect 41414 56896 41420 56908
rect 38948 56868 41420 56896
rect 12894 56788 12900 56840
rect 12952 56828 12958 56840
rect 20714 56828 20720 56840
rect 12952 56800 20720 56828
rect 12952 56788 12958 56800
rect 20714 56788 20720 56800
rect 20772 56788 20778 56840
rect 20806 56788 20812 56840
rect 20864 56828 20870 56840
rect 21453 56831 21511 56837
rect 21453 56828 21465 56831
rect 20864 56800 21465 56828
rect 20864 56788 20870 56800
rect 21453 56797 21465 56800
rect 21499 56797 21511 56831
rect 21453 56791 21511 56797
rect 28442 56788 28448 56840
rect 28500 56828 28506 56840
rect 38948 56837 38976 56868
rect 41414 56856 41420 56868
rect 41472 56856 41478 56908
rect 46198 56896 46204 56908
rect 44008 56868 46204 56896
rect 29825 56831 29883 56837
rect 29825 56828 29837 56831
rect 28500 56800 29837 56828
rect 28500 56788 28506 56800
rect 29825 56797 29837 56800
rect 29871 56797 29883 56831
rect 29825 56791 29883 56797
rect 30009 56831 30067 56837
rect 30009 56797 30021 56831
rect 30055 56797 30067 56831
rect 30009 56791 30067 56797
rect 38933 56831 38991 56837
rect 38933 56797 38945 56831
rect 38979 56797 38991 56831
rect 38933 56791 38991 56797
rect 39025 56831 39083 56837
rect 39025 56797 39037 56831
rect 39071 56797 39083 56831
rect 39206 56828 39212 56840
rect 39167 56800 39212 56828
rect 39025 56791 39083 56797
rect 17402 56760 17408 56772
rect 17363 56732 17408 56760
rect 17402 56720 17408 56732
rect 17460 56720 17466 56772
rect 21269 56763 21327 56769
rect 21269 56729 21281 56763
rect 21315 56760 21327 56763
rect 21358 56760 21364 56772
rect 21315 56732 21364 56760
rect 21315 56729 21327 56732
rect 21269 56723 21327 56729
rect 21358 56720 21364 56732
rect 21416 56720 21422 56772
rect 28258 56720 28264 56772
rect 28316 56760 28322 56772
rect 30024 56760 30052 56791
rect 28316 56732 30052 56760
rect 28316 56720 28322 56732
rect 38654 56720 38660 56772
rect 38712 56760 38718 56772
rect 39040 56760 39068 56791
rect 39206 56788 39212 56800
rect 39264 56788 39270 56840
rect 39298 56788 39304 56840
rect 39356 56828 39362 56840
rect 39356 56800 39401 56828
rect 39356 56788 39362 56800
rect 43530 56788 43536 56840
rect 43588 56837 43594 56840
rect 44008 56837 44036 56868
rect 46198 56856 46204 56868
rect 46256 56856 46262 56908
rect 43588 56831 43637 56837
rect 43588 56797 43591 56831
rect 43625 56797 43637 56831
rect 43588 56791 43637 56797
rect 43992 56831 44050 56837
rect 43992 56797 44004 56831
rect 44038 56797 44050 56831
rect 43992 56791 44050 56797
rect 43588 56788 43594 56791
rect 44082 56788 44088 56840
rect 44140 56828 44146 56840
rect 57054 56828 57060 56840
rect 44140 56800 44185 56828
rect 57015 56800 57060 56828
rect 44140 56788 44146 56800
rect 57054 56788 57060 56800
rect 57112 56788 57118 56840
rect 57514 56828 57520 56840
rect 57475 56800 57520 56828
rect 57514 56788 57520 56800
rect 57572 56788 57578 56840
rect 58342 56828 58348 56840
rect 58303 56800 58348 56828
rect 58342 56788 58348 56800
rect 58400 56788 58406 56840
rect 39574 56760 39580 56772
rect 38712 56732 39580 56760
rect 38712 56720 38718 56732
rect 39574 56720 39580 56732
rect 39632 56720 39638 56772
rect 43717 56763 43775 56769
rect 43717 56729 43729 56763
rect 43763 56729 43775 56763
rect 43717 56723 43775 56729
rect 17034 56652 17040 56704
rect 17092 56692 17098 56704
rect 25958 56692 25964 56704
rect 17092 56664 25964 56692
rect 17092 56652 17098 56664
rect 25958 56652 25964 56664
rect 26016 56652 26022 56704
rect 30098 56652 30104 56704
rect 30156 56692 30162 56704
rect 30193 56695 30251 56701
rect 30193 56692 30205 56695
rect 30156 56664 30205 56692
rect 30156 56652 30162 56664
rect 30193 56661 30205 56664
rect 30239 56661 30251 56695
rect 30193 56655 30251 56661
rect 35894 56652 35900 56704
rect 35952 56692 35958 56704
rect 38749 56695 38807 56701
rect 38749 56692 38761 56695
rect 35952 56664 38761 56692
rect 35952 56652 35958 56664
rect 38749 56661 38761 56664
rect 38795 56661 38807 56695
rect 43438 56692 43444 56704
rect 43399 56664 43444 56692
rect 38749 56655 38807 56661
rect 43438 56652 43444 56664
rect 43496 56652 43502 56704
rect 43732 56692 43760 56723
rect 43806 56720 43812 56772
rect 43864 56760 43870 56772
rect 55861 56763 55919 56769
rect 43864 56732 43909 56760
rect 43864 56720 43870 56732
rect 55861 56729 55873 56763
rect 55907 56760 55919 56763
rect 58360 56760 58388 56788
rect 55907 56732 58388 56760
rect 55907 56729 55919 56732
rect 55861 56723 55919 56729
rect 53374 56692 53380 56704
rect 43732 56664 53380 56692
rect 53374 56652 53380 56664
rect 53432 56652 53438 56704
rect 56778 56652 56784 56704
rect 56836 56692 56842 56704
rect 56873 56695 56931 56701
rect 56873 56692 56885 56695
rect 56836 56664 56885 56692
rect 56836 56652 56842 56664
rect 56873 56661 56885 56664
rect 56919 56661 56931 56695
rect 56873 56655 56931 56661
rect 57701 56695 57759 56701
rect 57701 56661 57713 56695
rect 57747 56692 57759 56695
rect 57882 56692 57888 56704
rect 57747 56664 57888 56692
rect 57747 56661 57759 56664
rect 57701 56655 57759 56661
rect 57882 56652 57888 56664
rect 57940 56652 57946 56704
rect 58066 56652 58072 56704
rect 58124 56692 58130 56704
rect 58161 56695 58219 56701
rect 58161 56692 58173 56695
rect 58124 56664 58173 56692
rect 58124 56652 58130 56664
rect 58161 56661 58173 56664
rect 58207 56661 58219 56695
rect 58161 56655 58219 56661
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 22002 56448 22008 56500
rect 22060 56488 22066 56500
rect 28718 56488 28724 56500
rect 22060 56448 22094 56488
rect 17862 56380 17868 56432
rect 17920 56420 17926 56432
rect 21269 56423 21327 56429
rect 21269 56420 21281 56423
rect 17920 56392 21281 56420
rect 17920 56380 17926 56392
rect 21269 56389 21281 56392
rect 21315 56389 21327 56423
rect 22066 56420 22094 56448
rect 23676 56460 28724 56488
rect 23676 56429 23704 56460
rect 28718 56448 28724 56460
rect 28776 56448 28782 56500
rect 28902 56448 28908 56500
rect 28960 56488 28966 56500
rect 30561 56491 30619 56497
rect 28960 56460 30420 56488
rect 28960 56448 28966 56460
rect 23569 56423 23627 56429
rect 23569 56420 23581 56423
rect 22066 56392 23581 56420
rect 21269 56383 21327 56389
rect 23569 56389 23581 56392
rect 23615 56389 23627 56423
rect 23569 56383 23627 56389
rect 23661 56423 23719 56429
rect 23661 56389 23673 56423
rect 23707 56389 23719 56423
rect 23661 56383 23719 56389
rect 24762 56380 24768 56432
rect 24820 56420 24826 56432
rect 25590 56420 25596 56432
rect 24820 56392 25360 56420
rect 24820 56380 24826 56392
rect 21085 56355 21143 56361
rect 21085 56321 21097 56355
rect 21131 56352 21143 56355
rect 21358 56352 21364 56364
rect 21131 56324 21364 56352
rect 21131 56321 21143 56324
rect 21085 56315 21143 56321
rect 21358 56312 21364 56324
rect 21416 56352 21422 56364
rect 21818 56352 21824 56364
rect 21416 56324 21824 56352
rect 21416 56312 21422 56324
rect 21818 56312 21824 56324
rect 21876 56352 21882 56364
rect 22005 56355 22063 56361
rect 22005 56352 22017 56355
rect 21876 56324 22017 56352
rect 21876 56312 21882 56324
rect 22005 56321 22017 56324
rect 22051 56321 22063 56355
rect 22005 56315 22063 56321
rect 22094 56312 22100 56364
rect 22152 56352 22158 56364
rect 23474 56361 23480 56364
rect 22189 56355 22247 56361
rect 22189 56352 22201 56355
rect 22152 56324 22201 56352
rect 22152 56312 22158 56324
rect 22189 56321 22201 56324
rect 22235 56321 22247 56355
rect 22189 56315 22247 56321
rect 23472 56315 23480 56361
rect 23532 56352 23538 56364
rect 23842 56352 23848 56364
rect 23532 56324 23572 56352
rect 23803 56324 23848 56352
rect 23474 56312 23480 56315
rect 23532 56312 23538 56324
rect 23842 56312 23848 56324
rect 23900 56312 23906 56364
rect 23937 56355 23995 56361
rect 23937 56321 23949 56355
rect 23983 56321 23995 56355
rect 25038 56352 25044 56364
rect 24999 56324 25044 56352
rect 23937 56315 23995 56321
rect 23952 56284 23980 56315
rect 25038 56312 25044 56324
rect 25096 56312 25102 56364
rect 25332 56361 25360 56392
rect 25424 56392 25596 56420
rect 25317 56355 25375 56361
rect 25317 56321 25329 56355
rect 25363 56321 25375 56355
rect 25317 56315 25375 56321
rect 25424 56284 25452 56392
rect 25590 56380 25596 56392
rect 25648 56380 25654 56432
rect 26234 56420 26240 56432
rect 26195 56392 26240 56420
rect 26234 56380 26240 56392
rect 26292 56380 26298 56432
rect 28537 56423 28595 56429
rect 28537 56389 28549 56423
rect 28583 56420 28595 56423
rect 29822 56420 29828 56432
rect 28583 56392 29828 56420
rect 28583 56389 28595 56392
rect 28537 56383 28595 56389
rect 29822 56380 29828 56392
rect 29880 56380 29886 56432
rect 30190 56420 30196 56432
rect 30151 56392 30196 56420
rect 30190 56380 30196 56392
rect 30248 56380 30254 56432
rect 30305 56423 30363 56429
rect 30305 56389 30317 56423
rect 30351 56420 30363 56423
rect 30392 56420 30420 56460
rect 30561 56457 30573 56491
rect 30607 56488 30619 56491
rect 30926 56488 30932 56500
rect 30607 56460 30932 56488
rect 30607 56457 30619 56460
rect 30561 56451 30619 56457
rect 30926 56448 30932 56460
rect 30984 56448 30990 56500
rect 35158 56488 35164 56500
rect 35119 56460 35164 56488
rect 35158 56448 35164 56460
rect 35216 56448 35222 56500
rect 38289 56491 38347 56497
rect 38289 56488 38301 56491
rect 35268 56460 38301 56488
rect 30351 56392 30420 56420
rect 30351 56389 30363 56392
rect 30305 56383 30363 56389
rect 32490 56380 32496 56432
rect 32548 56420 32554 56432
rect 33045 56423 33103 56429
rect 33045 56420 33057 56423
rect 32548 56392 33057 56420
rect 32548 56380 32554 56392
rect 33045 56389 33057 56392
rect 33091 56389 33103 56423
rect 35268 56420 35296 56460
rect 38289 56457 38301 56460
rect 38335 56457 38347 56491
rect 38289 56451 38347 56457
rect 38378 56448 38384 56500
rect 38436 56488 38442 56500
rect 43438 56488 43444 56500
rect 38436 56460 43444 56488
rect 38436 56448 38442 56460
rect 43438 56448 43444 56460
rect 43496 56448 43502 56500
rect 57054 56448 57060 56500
rect 57112 56488 57118 56500
rect 57149 56491 57207 56497
rect 57149 56488 57161 56491
rect 57112 56460 57161 56488
rect 57112 56448 57118 56460
rect 57149 56457 57161 56460
rect 57195 56457 57207 56491
rect 57149 56451 57207 56457
rect 35434 56420 35440 56432
rect 33045 56383 33103 56389
rect 33336 56392 35296 56420
rect 35395 56392 35440 56420
rect 25961 56355 26019 56361
rect 25961 56352 25973 56355
rect 23952 56256 25452 56284
rect 25516 56324 25973 56352
rect 21453 56219 21511 56225
rect 21453 56185 21465 56219
rect 21499 56216 21511 56219
rect 25516 56216 25544 56324
rect 25961 56321 25973 56324
rect 26007 56321 26019 56355
rect 26142 56352 26148 56364
rect 26103 56324 26148 56352
rect 25961 56315 26019 56321
rect 26142 56312 26148 56324
rect 26200 56312 26206 56364
rect 26381 56355 26439 56361
rect 26381 56321 26393 56355
rect 26427 56352 26439 56355
rect 27338 56352 27344 56364
rect 26427 56324 27344 56352
rect 26427 56321 26439 56324
rect 26381 56315 26439 56321
rect 27338 56312 27344 56324
rect 27396 56312 27402 56364
rect 28261 56355 28319 56361
rect 28261 56321 28273 56355
rect 28307 56321 28319 56355
rect 28261 56315 28319 56321
rect 21499 56188 25544 56216
rect 21499 56185 21511 56188
rect 21453 56179 21511 56185
rect 25590 56176 25596 56228
rect 25648 56216 25654 56228
rect 28276 56216 28304 56315
rect 28350 56312 28356 56364
rect 28408 56352 28414 56364
rect 28626 56352 28632 56364
rect 28408 56324 28453 56352
rect 28587 56324 28632 56352
rect 28408 56312 28414 56324
rect 28626 56312 28632 56324
rect 28684 56312 28690 56364
rect 28767 56355 28825 56361
rect 28767 56321 28779 56355
rect 28813 56352 28825 56355
rect 28994 56352 29000 56364
rect 28813 56324 29000 56352
rect 28813 56321 28825 56324
rect 28767 56315 28825 56321
rect 28994 56312 29000 56324
rect 29052 56312 29058 56364
rect 29917 56355 29975 56361
rect 29917 56321 29929 56355
rect 29963 56321 29975 56355
rect 29917 56315 29975 56321
rect 30010 56355 30068 56361
rect 30010 56321 30022 56355
rect 30056 56342 30068 56355
rect 30098 56342 30104 56364
rect 30056 56321 30104 56342
rect 30010 56315 30104 56321
rect 29086 56284 29092 56296
rect 28460 56256 29092 56284
rect 28460 56216 28488 56256
rect 29086 56244 29092 56256
rect 29144 56284 29150 56296
rect 29932 56284 29960 56315
rect 30025 56314 30104 56315
rect 30098 56312 30104 56314
rect 30156 56312 30162 56364
rect 30382 56355 30440 56361
rect 30382 56321 30394 56355
rect 30428 56321 30440 56355
rect 30382 56315 30440 56321
rect 29144 56256 29960 56284
rect 29144 56244 29150 56256
rect 25648 56188 28488 56216
rect 25648 56176 25654 56188
rect 28718 56176 28724 56228
rect 28776 56216 28782 56228
rect 28776 56188 30052 56216
rect 28776 56176 28782 56188
rect 22373 56151 22431 56157
rect 22373 56117 22385 56151
rect 22419 56148 22431 56151
rect 23106 56148 23112 56160
rect 22419 56120 23112 56148
rect 22419 56117 22431 56120
rect 22373 56111 22431 56117
rect 23106 56108 23112 56120
rect 23164 56108 23170 56160
rect 23290 56148 23296 56160
rect 23251 56120 23296 56148
rect 23290 56108 23296 56120
rect 23348 56108 23354 56160
rect 25133 56151 25191 56157
rect 25133 56117 25145 56151
rect 25179 56148 25191 56151
rect 25222 56148 25228 56160
rect 25179 56120 25228 56148
rect 25179 56117 25191 56120
rect 25133 56111 25191 56117
rect 25222 56108 25228 56120
rect 25280 56108 25286 56160
rect 25501 56151 25559 56157
rect 25501 56117 25513 56151
rect 25547 56148 25559 56151
rect 25866 56148 25872 56160
rect 25547 56120 25872 56148
rect 25547 56117 25559 56120
rect 25501 56111 25559 56117
rect 25866 56108 25872 56120
rect 25924 56108 25930 56160
rect 26513 56151 26571 56157
rect 26513 56117 26525 56151
rect 26559 56148 26571 56151
rect 27246 56148 27252 56160
rect 26559 56120 27252 56148
rect 26559 56117 26571 56120
rect 26513 56111 26571 56117
rect 27246 56108 27252 56120
rect 27304 56108 27310 56160
rect 28905 56151 28963 56157
rect 28905 56117 28917 56151
rect 28951 56148 28963 56151
rect 29914 56148 29920 56160
rect 28951 56120 29920 56148
rect 28951 56117 28963 56120
rect 28905 56111 28963 56117
rect 29914 56108 29920 56120
rect 29972 56108 29978 56160
rect 30024 56148 30052 56188
rect 30098 56176 30104 56228
rect 30156 56216 30162 56228
rect 30392 56216 30420 56315
rect 30558 56312 30564 56364
rect 30616 56352 30622 56364
rect 31021 56355 31079 56361
rect 31021 56352 31033 56355
rect 30616 56324 31033 56352
rect 30616 56312 30622 56324
rect 31021 56321 31033 56324
rect 31067 56321 31079 56355
rect 31021 56315 31079 56321
rect 31110 56312 31116 56364
rect 31168 56352 31174 56364
rect 31205 56355 31263 56361
rect 31205 56352 31217 56355
rect 31168 56324 31217 56352
rect 31168 56312 31174 56324
rect 31205 56321 31217 56324
rect 31251 56321 31263 56355
rect 31205 56315 31263 56321
rect 31294 56312 31300 56364
rect 31352 56352 31358 56364
rect 31478 56361 31484 56364
rect 31441 56355 31484 56361
rect 31352 56324 31397 56352
rect 31352 56312 31358 56324
rect 31441 56321 31453 56355
rect 31441 56315 31484 56321
rect 31478 56312 31484 56315
rect 31536 56312 31542 56364
rect 32950 56361 32956 56364
rect 32948 56352 32956 56361
rect 32911 56324 32956 56352
rect 32948 56315 32956 56324
rect 32950 56312 32956 56315
rect 33008 56312 33014 56364
rect 33336 56361 33364 56392
rect 35434 56380 35440 56392
rect 35492 56380 35498 56432
rect 36538 56420 36544 56432
rect 36499 56392 36544 56420
rect 36538 56380 36544 56392
rect 36596 56380 36602 56432
rect 38194 56420 38200 56432
rect 36831 56392 38200 56420
rect 33137 56355 33195 56361
rect 33137 56321 33149 56355
rect 33183 56321 33195 56355
rect 33137 56315 33195 56321
rect 33320 56355 33378 56361
rect 33320 56321 33332 56355
rect 33366 56321 33378 56355
rect 33320 56315 33378 56321
rect 33413 56355 33471 56361
rect 33413 56321 33425 56355
rect 33459 56352 33471 56355
rect 33502 56352 33508 56364
rect 33459 56324 33508 56352
rect 33459 56321 33471 56324
rect 33413 56315 33471 56321
rect 30156 56188 30420 56216
rect 31573 56219 31631 56225
rect 30156 56176 30162 56188
rect 31573 56185 31585 56219
rect 31619 56216 31631 56219
rect 33152 56216 33180 56315
rect 33502 56312 33508 56324
rect 33560 56312 33566 56364
rect 35342 56361 35348 56364
rect 35340 56352 35348 56361
rect 35303 56324 35348 56352
rect 35340 56315 35348 56324
rect 35342 56312 35348 56315
rect 35400 56312 35406 56364
rect 35526 56352 35532 56364
rect 35487 56324 35532 56352
rect 35526 56312 35532 56324
rect 35584 56312 35590 56364
rect 35710 56352 35716 56364
rect 35671 56324 35716 56352
rect 35710 56312 35716 56324
rect 35768 56312 35774 56364
rect 35802 56312 35808 56364
rect 35860 56352 35866 56364
rect 36446 56361 36452 56364
rect 35860 56324 35905 56352
rect 35860 56312 35866 56324
rect 36444 56315 36452 56361
rect 36504 56352 36510 56364
rect 36504 56324 36544 56352
rect 36446 56312 36452 56315
rect 36504 56312 36510 56324
rect 36630 56312 36636 56364
rect 36688 56352 36694 56364
rect 36831 56361 36859 56392
rect 38194 56380 38200 56392
rect 38252 56380 38258 56432
rect 39022 56420 39028 56432
rect 38488 56392 39028 56420
rect 36816 56355 36874 56361
rect 36688 56324 36733 56352
rect 36688 56312 36694 56324
rect 36816 56321 36828 56355
rect 36862 56321 36874 56355
rect 36816 56315 36874 56321
rect 36906 56312 36912 56364
rect 36964 56352 36970 56364
rect 38488 56361 38516 56392
rect 39022 56380 39028 56392
rect 39080 56380 39086 56432
rect 39206 56380 39212 56432
rect 39264 56420 39270 56432
rect 41509 56423 41567 56429
rect 39264 56392 39436 56420
rect 39264 56380 39270 56392
rect 38473 56355 38531 56361
rect 36964 56324 37009 56352
rect 36964 56312 36970 56324
rect 38473 56321 38485 56355
rect 38519 56321 38531 56355
rect 38473 56315 38531 56321
rect 38565 56355 38623 56361
rect 38565 56321 38577 56355
rect 38611 56352 38623 56355
rect 38654 56352 38660 56364
rect 38611 56324 38660 56352
rect 38611 56321 38623 56324
rect 38565 56315 38623 56321
rect 38654 56312 38660 56324
rect 38712 56312 38718 56364
rect 38749 56355 38807 56361
rect 38749 56321 38761 56355
rect 38795 56321 38807 56355
rect 38749 56315 38807 56321
rect 36722 56244 36728 56296
rect 36780 56284 36786 56296
rect 38764 56284 38792 56315
rect 38838 56312 38844 56364
rect 38896 56352 38902 56364
rect 39298 56352 39304 56364
rect 38896 56324 39304 56352
rect 38896 56312 38902 56324
rect 39298 56312 39304 56324
rect 39356 56312 39362 56364
rect 39408 56361 39436 56392
rect 41509 56389 41521 56423
rect 41555 56420 41567 56423
rect 52178 56420 52184 56432
rect 41555 56392 52184 56420
rect 41555 56389 41567 56392
rect 41509 56383 41567 56389
rect 52178 56380 52184 56392
rect 52236 56380 52242 56432
rect 56689 56423 56747 56429
rect 56689 56389 56701 56423
rect 56735 56420 56747 56423
rect 57514 56420 57520 56432
rect 56735 56392 57520 56420
rect 56735 56389 56747 56392
rect 56689 56383 56747 56389
rect 57514 56380 57520 56392
rect 57572 56380 57578 56432
rect 39393 56355 39451 56361
rect 39393 56321 39405 56355
rect 39439 56321 39451 56355
rect 39574 56352 39580 56364
rect 39535 56324 39580 56352
rect 39393 56315 39451 56321
rect 38930 56284 38936 56296
rect 36780 56256 38936 56284
rect 36780 56244 36786 56256
rect 38930 56244 38936 56256
rect 38988 56284 38994 56296
rect 39408 56284 39436 56315
rect 39574 56312 39580 56324
rect 39632 56312 39638 56364
rect 39669 56355 39727 56361
rect 39669 56321 39681 56355
rect 39715 56352 39727 56355
rect 40494 56352 40500 56364
rect 39715 56324 40500 56352
rect 39715 56321 39727 56324
rect 39669 56315 39727 56321
rect 40494 56312 40500 56324
rect 40552 56312 40558 56364
rect 41412 56355 41470 56361
rect 41412 56321 41424 56355
rect 41458 56352 41470 56355
rect 41601 56355 41659 56361
rect 41458 56324 41552 56352
rect 41458 56321 41470 56324
rect 41412 56315 41470 56321
rect 41524 56296 41552 56324
rect 41601 56321 41613 56355
rect 41647 56352 41659 56355
rect 41690 56352 41696 56364
rect 41647 56324 41696 56352
rect 41647 56321 41659 56324
rect 41601 56315 41659 56321
rect 41690 56312 41696 56324
rect 41748 56312 41754 56364
rect 41784 56355 41842 56361
rect 41784 56321 41796 56355
rect 41830 56321 41842 56355
rect 41784 56315 41842 56321
rect 41877 56355 41935 56361
rect 41877 56321 41889 56355
rect 41923 56352 41935 56355
rect 42150 56352 42156 56364
rect 41923 56324 42156 56352
rect 41923 56321 41935 56324
rect 41877 56315 41935 56321
rect 38988 56256 39436 56284
rect 38988 56244 38994 56256
rect 41506 56244 41512 56296
rect 41564 56244 41570 56296
rect 41800 56284 41828 56315
rect 42150 56312 42156 56324
rect 42208 56312 42214 56364
rect 43438 56361 43444 56364
rect 43436 56352 43444 56361
rect 43399 56324 43444 56352
rect 43436 56315 43444 56324
rect 43438 56312 43444 56315
rect 43496 56312 43502 56364
rect 43533 56355 43591 56361
rect 43533 56321 43545 56355
rect 43579 56321 43591 56355
rect 43533 56315 43591 56321
rect 42794 56284 42800 56296
rect 41800 56256 42800 56284
rect 42794 56244 42800 56256
rect 42852 56244 42858 56296
rect 33410 56216 33416 56228
rect 31619 56188 32904 56216
rect 33152 56188 33416 56216
rect 31619 56185 31631 56188
rect 31573 56179 31631 56185
rect 32769 56151 32827 56157
rect 32769 56148 32781 56151
rect 30024 56120 32781 56148
rect 32769 56117 32781 56120
rect 32815 56117 32827 56151
rect 32876 56148 32904 56188
rect 33410 56176 33416 56188
rect 33468 56176 33474 56228
rect 36262 56216 36268 56228
rect 36223 56188 36268 56216
rect 36262 56176 36268 56188
rect 36320 56176 36326 56228
rect 36630 56176 36636 56228
rect 36688 56216 36694 56228
rect 43257 56219 43315 56225
rect 43257 56216 43269 56219
rect 36688 56188 43269 56216
rect 36688 56176 36694 56188
rect 43257 56185 43269 56188
rect 43303 56185 43315 56219
rect 43257 56179 43315 56185
rect 33318 56148 33324 56160
rect 32876 56120 33324 56148
rect 32769 56111 32827 56117
rect 33318 56108 33324 56120
rect 33376 56108 33382 56160
rect 35710 56108 35716 56160
rect 35768 56148 35774 56160
rect 39853 56151 39911 56157
rect 39853 56148 39865 56151
rect 35768 56120 39865 56148
rect 35768 56108 35774 56120
rect 39853 56117 39865 56120
rect 39899 56117 39911 56151
rect 41230 56148 41236 56160
rect 41191 56120 41236 56148
rect 39853 56111 39911 56117
rect 41230 56108 41236 56120
rect 41288 56108 41294 56160
rect 43548 56148 43576 56315
rect 43622 56312 43628 56364
rect 43680 56352 43686 56364
rect 43808 56355 43866 56361
rect 43680 56324 43725 56352
rect 43680 56312 43686 56324
rect 43808 56321 43820 56355
rect 43854 56321 43866 56355
rect 43808 56315 43866 56321
rect 43824 56216 43852 56315
rect 43898 56312 43904 56364
rect 43956 56352 43962 56364
rect 44082 56352 44088 56364
rect 43956 56324 44088 56352
rect 43956 56312 43962 56324
rect 44082 56312 44088 56324
rect 44140 56312 44146 56364
rect 56137 56355 56195 56361
rect 56137 56321 56149 56355
rect 56183 56352 56195 56355
rect 57974 56352 57980 56364
rect 56183 56324 57980 56352
rect 56183 56321 56195 56324
rect 56137 56315 56195 56321
rect 57974 56312 57980 56324
rect 58032 56312 58038 56364
rect 58345 56355 58403 56361
rect 58345 56321 58357 56355
rect 58391 56352 58403 56355
rect 58434 56352 58440 56364
rect 58391 56324 58440 56352
rect 58391 56321 58403 56324
rect 58345 56315 58403 56321
rect 58434 56312 58440 56324
rect 58492 56312 58498 56364
rect 58158 56284 58164 56296
rect 51046 56256 58164 56284
rect 44266 56216 44272 56228
rect 43824 56188 44272 56216
rect 44266 56176 44272 56188
rect 44324 56176 44330 56228
rect 51046 56148 51074 56256
rect 58158 56244 58164 56256
rect 58216 56244 58222 56296
rect 58158 56148 58164 56160
rect 43548 56120 51074 56148
rect 58119 56120 58164 56148
rect 58158 56108 58164 56120
rect 58216 56108 58222 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 6914 55904 6920 55956
rect 6972 55944 6978 55956
rect 6972 55916 22094 55944
rect 6972 55904 6978 55916
rect 22066 55808 22094 55916
rect 23842 55904 23848 55956
rect 23900 55944 23906 55956
rect 24581 55947 24639 55953
rect 24581 55944 24593 55947
rect 23900 55916 24593 55944
rect 23900 55904 23906 55916
rect 24581 55913 24593 55916
rect 24627 55913 24639 55947
rect 24581 55907 24639 55913
rect 26142 55904 26148 55956
rect 26200 55944 26206 55956
rect 26237 55947 26295 55953
rect 26237 55944 26249 55947
rect 26200 55916 26249 55944
rect 26200 55904 26206 55916
rect 26237 55913 26249 55916
rect 26283 55913 26295 55947
rect 26237 55907 26295 55913
rect 28077 55947 28135 55953
rect 28077 55913 28089 55947
rect 28123 55944 28135 55947
rect 28350 55944 28356 55956
rect 28123 55916 28356 55944
rect 28123 55913 28135 55916
rect 28077 55907 28135 55913
rect 28350 55904 28356 55916
rect 28408 55904 28414 55956
rect 28442 55904 28448 55956
rect 28500 55944 28506 55956
rect 28500 55916 28545 55944
rect 28500 55904 28506 55916
rect 28994 55904 29000 55956
rect 29052 55944 29058 55956
rect 30098 55944 30104 55956
rect 29052 55916 30104 55944
rect 29052 55904 29058 55916
rect 30098 55904 30104 55916
rect 30156 55904 30162 55956
rect 32950 55904 32956 55956
rect 33008 55944 33014 55956
rect 35066 55944 35072 55956
rect 33008 55916 35072 55944
rect 33008 55904 33014 55916
rect 35066 55904 35072 55916
rect 35124 55944 35130 55956
rect 36446 55944 36452 55956
rect 35124 55916 36452 55944
rect 35124 55904 35130 55916
rect 36446 55904 36452 55916
rect 36504 55904 36510 55956
rect 38194 55904 38200 55956
rect 38252 55944 38258 55956
rect 38473 55947 38531 55953
rect 38473 55944 38485 55947
rect 38252 55916 38485 55944
rect 38252 55904 38258 55916
rect 38473 55913 38485 55916
rect 38519 55913 38531 55947
rect 38473 55907 38531 55913
rect 42150 55904 42156 55956
rect 42208 55944 42214 55956
rect 43898 55944 43904 55956
rect 42208 55916 43904 55944
rect 42208 55904 42214 55916
rect 43898 55904 43904 55916
rect 43956 55904 43962 55956
rect 57149 55947 57207 55953
rect 57149 55913 57161 55947
rect 57195 55944 57207 55947
rect 58434 55944 58440 55956
rect 57195 55916 58440 55944
rect 57195 55913 57207 55916
rect 57149 55907 57207 55913
rect 58434 55904 58440 55916
rect 58492 55904 58498 55956
rect 23661 55879 23719 55885
rect 23661 55845 23673 55879
rect 23707 55876 23719 55879
rect 23750 55876 23756 55888
rect 23707 55848 23756 55876
rect 23707 55845 23719 55848
rect 23661 55839 23719 55845
rect 23750 55836 23756 55848
rect 23808 55836 23814 55888
rect 24780 55848 25728 55876
rect 24780 55808 24808 55848
rect 22066 55780 24808 55808
rect 24854 55768 24860 55820
rect 24912 55808 24918 55820
rect 25041 55811 25099 55817
rect 25041 55808 25053 55811
rect 24912 55780 25053 55808
rect 24912 55768 24918 55780
rect 25041 55777 25053 55780
rect 25087 55777 25099 55811
rect 25700 55808 25728 55848
rect 25774 55836 25780 55888
rect 25832 55876 25838 55888
rect 30282 55876 30288 55888
rect 25832 55848 30144 55876
rect 30243 55848 30288 55876
rect 25832 55836 25838 55848
rect 27062 55808 27068 55820
rect 25700 55780 27068 55808
rect 25041 55771 25099 55777
rect 27062 55768 27068 55780
rect 27120 55768 27126 55820
rect 27338 55768 27344 55820
rect 27396 55808 27402 55820
rect 28534 55808 28540 55820
rect 27396 55780 28396 55808
rect 28495 55780 28540 55808
rect 27396 55768 27402 55780
rect 1762 55700 1768 55752
rect 1820 55740 1826 55752
rect 1857 55743 1915 55749
rect 1857 55740 1869 55743
rect 1820 55712 1869 55740
rect 1820 55700 1826 55712
rect 1857 55709 1869 55712
rect 1903 55740 1915 55743
rect 2317 55743 2375 55749
rect 2317 55740 2329 55743
rect 1903 55712 2329 55740
rect 1903 55709 1915 55712
rect 1857 55703 1915 55709
rect 2317 55709 2329 55712
rect 2363 55709 2375 55743
rect 2317 55703 2375 55709
rect 3418 55700 3424 55752
rect 3476 55740 3482 55752
rect 23106 55740 23112 55752
rect 3476 55712 22692 55740
rect 23067 55712 23112 55740
rect 3476 55700 3482 55712
rect 21269 55675 21327 55681
rect 21269 55641 21281 55675
rect 21315 55672 21327 55675
rect 21358 55672 21364 55684
rect 21315 55644 21364 55672
rect 21315 55641 21327 55644
rect 21269 55635 21327 55641
rect 21358 55632 21364 55644
rect 21416 55632 21422 55684
rect 22664 55681 22692 55712
rect 23106 55700 23112 55712
rect 23164 55700 23170 55752
rect 23290 55740 23296 55752
rect 23251 55712 23296 55740
rect 23290 55700 23296 55712
rect 23348 55700 23354 55752
rect 23529 55743 23587 55749
rect 23529 55709 23541 55743
rect 23575 55740 23587 55743
rect 23934 55740 23940 55752
rect 23575 55712 23940 55740
rect 23575 55709 23587 55712
rect 23529 55703 23587 55709
rect 23934 55700 23940 55712
rect 23992 55700 23998 55752
rect 24762 55740 24768 55752
rect 24723 55712 24768 55740
rect 24762 55700 24768 55712
rect 24820 55700 24826 55752
rect 24949 55743 25007 55749
rect 24949 55709 24961 55743
rect 24995 55740 25007 55743
rect 25222 55740 25228 55752
rect 24995 55712 25228 55740
rect 24995 55709 25007 55712
rect 24949 55703 25007 55709
rect 25222 55700 25228 55712
rect 25280 55700 25286 55752
rect 25590 55740 25596 55752
rect 25551 55712 25596 55740
rect 25590 55700 25596 55712
rect 25648 55700 25654 55752
rect 25774 55749 25780 55752
rect 25741 55743 25780 55749
rect 25741 55709 25753 55743
rect 25741 55703 25780 55709
rect 25774 55700 25780 55703
rect 25832 55700 25838 55752
rect 25866 55700 25872 55752
rect 25924 55740 25930 55752
rect 25924 55712 25969 55740
rect 25924 55700 25930 55712
rect 26050 55700 26056 55752
rect 26108 55749 26114 55752
rect 26108 55740 26116 55749
rect 28258 55740 28264 55752
rect 26108 55712 26153 55740
rect 28219 55712 28264 55740
rect 26108 55703 26116 55712
rect 26108 55700 26114 55703
rect 28258 55700 28264 55712
rect 28316 55700 28322 55752
rect 28368 55740 28396 55780
rect 28534 55768 28540 55780
rect 28592 55768 28598 55820
rect 30116 55808 30144 55848
rect 30282 55836 30288 55848
rect 30340 55836 30346 55888
rect 41230 55876 41236 55888
rect 33428 55848 41236 55876
rect 28644 55780 30052 55808
rect 30116 55780 31754 55808
rect 28644 55740 28672 55780
rect 28368 55712 28672 55740
rect 29733 55743 29791 55749
rect 29733 55709 29745 55743
rect 29779 55709 29791 55743
rect 29914 55740 29920 55752
rect 29875 55712 29920 55740
rect 29733 55703 29791 55709
rect 21453 55675 21511 55681
rect 21453 55641 21465 55675
rect 21499 55641 21511 55675
rect 21453 55635 21511 55641
rect 21637 55675 21695 55681
rect 21637 55641 21649 55675
rect 21683 55672 21695 55675
rect 22649 55675 22707 55681
rect 21683 55644 22094 55672
rect 21683 55641 21695 55644
rect 21637 55635 21695 55641
rect 1670 55604 1676 55616
rect 1631 55576 1676 55604
rect 1670 55564 1676 55576
rect 1728 55564 1734 55616
rect 18966 55564 18972 55616
rect 19024 55604 19030 55616
rect 21468 55604 21496 55635
rect 19024 55576 21496 55604
rect 22066 55604 22094 55644
rect 22649 55641 22661 55675
rect 22695 55672 22707 55675
rect 23385 55675 23443 55681
rect 23385 55672 23397 55675
rect 22695 55644 23397 55672
rect 22695 55641 22707 55644
rect 22649 55635 22707 55641
rect 23385 55641 23397 55644
rect 23431 55641 23443 55675
rect 25958 55672 25964 55684
rect 25919 55644 25964 55672
rect 23385 55635 23443 55641
rect 25958 55632 25964 55644
rect 26016 55632 26022 55684
rect 29748 55672 29776 55703
rect 29914 55700 29920 55712
rect 29972 55700 29978 55752
rect 30024 55740 30052 55780
rect 30190 55749 30196 55752
rect 30153 55743 30196 55749
rect 30153 55740 30165 55743
rect 30024 55712 30165 55740
rect 30153 55709 30165 55712
rect 30248 55740 30254 55752
rect 31478 55740 31484 55752
rect 30248 55712 31484 55740
rect 30153 55703 30196 55709
rect 30190 55700 30196 55703
rect 30248 55700 30254 55712
rect 31478 55700 31484 55712
rect 31536 55700 31542 55752
rect 26068 55644 29776 55672
rect 30009 55675 30067 55681
rect 26068 55604 26096 55644
rect 30009 55641 30021 55675
rect 30055 55641 30067 55675
rect 30009 55635 30067 55641
rect 22066 55576 26096 55604
rect 19024 55564 19030 55576
rect 27062 55564 27068 55616
rect 27120 55604 27126 55616
rect 29089 55607 29147 55613
rect 29089 55604 29101 55607
rect 27120 55576 29101 55604
rect 27120 55564 27126 55576
rect 29089 55573 29101 55576
rect 29135 55604 29147 55607
rect 30024 55604 30052 55635
rect 30834 55604 30840 55616
rect 29135 55576 30052 55604
rect 30795 55576 30840 55604
rect 29135 55573 29147 55576
rect 29089 55567 29147 55573
rect 30834 55564 30840 55576
rect 30892 55604 30898 55616
rect 31294 55604 31300 55616
rect 30892 55576 31300 55604
rect 30892 55564 30898 55576
rect 31294 55564 31300 55576
rect 31352 55564 31358 55616
rect 31726 55604 31754 55780
rect 32950 55700 32956 55752
rect 33008 55749 33014 55752
rect 33008 55743 33057 55749
rect 33008 55709 33011 55743
rect 33045 55709 33057 55743
rect 33134 55740 33140 55752
rect 33095 55712 33140 55740
rect 33008 55703 33057 55709
rect 33008 55700 33014 55703
rect 33134 55700 33140 55712
rect 33192 55700 33198 55752
rect 33428 55749 33456 55848
rect 41230 55836 41236 55848
rect 41288 55836 41294 55888
rect 41874 55836 41880 55888
rect 41932 55876 41938 55888
rect 43622 55876 43628 55888
rect 41932 55848 43628 55876
rect 41932 55836 41938 55848
rect 43622 55836 43628 55848
rect 43680 55836 43686 55888
rect 36265 55811 36323 55817
rect 36265 55808 36277 55811
rect 34716 55780 36277 55808
rect 33229 55743 33287 55749
rect 33229 55709 33241 55743
rect 33275 55709 33287 55743
rect 33229 55703 33287 55709
rect 33412 55743 33470 55749
rect 33412 55709 33424 55743
rect 33458 55709 33470 55743
rect 33412 55703 33470 55709
rect 33244 55672 33272 55703
rect 33502 55700 33508 55752
rect 33560 55740 33566 55752
rect 34606 55740 34612 55752
rect 33560 55712 34612 55740
rect 33560 55700 33566 55712
rect 34606 55700 34612 55712
rect 34664 55700 34670 55752
rect 34716 55672 34744 55780
rect 36265 55777 36277 55780
rect 36311 55777 36323 55811
rect 37182 55808 37188 55820
rect 36265 55771 36323 55777
rect 36464 55780 37188 55808
rect 35066 55749 35072 55752
rect 35064 55740 35072 55749
rect 35027 55712 35072 55740
rect 35064 55703 35072 55712
rect 35124 55740 35130 55752
rect 35342 55740 35348 55752
rect 35124 55712 35348 55740
rect 35066 55700 35072 55703
rect 35124 55700 35130 55712
rect 35342 55700 35348 55712
rect 35400 55700 35406 55752
rect 35436 55743 35494 55749
rect 35436 55709 35448 55743
rect 35482 55709 35494 55743
rect 35436 55703 35494 55709
rect 35529 55743 35587 55749
rect 35529 55709 35541 55743
rect 35575 55740 35587 55743
rect 35802 55740 35808 55752
rect 35575 55712 35808 55740
rect 35575 55709 35587 55712
rect 35529 55703 35587 55709
rect 33244 55644 34744 55672
rect 34790 55632 34796 55684
rect 34848 55672 34854 55684
rect 35161 55675 35219 55681
rect 35161 55672 35173 55675
rect 34848 55644 35173 55672
rect 34848 55632 34854 55644
rect 35161 55641 35173 55644
rect 35207 55641 35219 55675
rect 35161 55635 35219 55641
rect 35250 55632 35256 55684
rect 35308 55672 35314 55684
rect 35452 55672 35480 55703
rect 35802 55700 35808 55712
rect 35860 55700 35866 55752
rect 36464 55749 36492 55780
rect 37182 55768 37188 55780
rect 37240 55768 37246 55820
rect 40034 55808 40040 55820
rect 38672 55780 40040 55808
rect 36449 55743 36507 55749
rect 36449 55709 36461 55743
rect 36495 55709 36507 55743
rect 36449 55703 36507 55709
rect 36538 55700 36544 55752
rect 36596 55740 36602 55752
rect 36722 55740 36728 55752
rect 36596 55712 36641 55740
rect 36683 55712 36728 55740
rect 36596 55700 36602 55712
rect 36722 55700 36728 55712
rect 36780 55700 36786 55752
rect 36814 55700 36820 55752
rect 36872 55740 36878 55752
rect 38672 55749 38700 55780
rect 40034 55768 40040 55780
rect 40092 55768 40098 55820
rect 41892 55780 42656 55808
rect 38657 55743 38715 55749
rect 36872 55712 36917 55740
rect 36872 55700 36878 55712
rect 38657 55709 38669 55743
rect 38703 55709 38715 55743
rect 38657 55703 38715 55709
rect 38746 55700 38752 55752
rect 38804 55740 38810 55752
rect 38918 55743 38976 55749
rect 38804 55712 38849 55740
rect 38804 55700 38810 55712
rect 38918 55709 38930 55743
rect 38964 55730 38976 55743
rect 38918 55703 38936 55709
rect 35894 55672 35900 55684
rect 35308 55644 35353 55672
rect 35452 55644 35900 55672
rect 35308 55632 35314 55644
rect 35894 55632 35900 55644
rect 35952 55632 35958 55684
rect 38930 55678 38936 55703
rect 38988 55678 38994 55730
rect 39022 55700 39028 55752
rect 39080 55734 39086 55752
rect 39080 55706 39119 55734
rect 39080 55700 39086 55706
rect 41506 55700 41512 55752
rect 41564 55740 41570 55752
rect 41647 55743 41705 55749
rect 41647 55740 41659 55743
rect 41564 55712 41659 55740
rect 41564 55700 41570 55712
rect 41647 55709 41659 55712
rect 41693 55740 41705 55743
rect 41892 55740 41920 55780
rect 41693 55712 41920 55740
rect 42060 55743 42118 55749
rect 41693 55709 41705 55712
rect 41647 55703 41705 55709
rect 42060 55709 42072 55743
rect 42106 55709 42118 55743
rect 42060 55703 42118 55709
rect 39025 55697 39083 55700
rect 41785 55675 41843 55681
rect 37844 55644 38884 55672
rect 32861 55607 32919 55613
rect 32861 55604 32873 55607
rect 31726 55576 32873 55604
rect 32861 55573 32873 55576
rect 32907 55573 32919 55607
rect 32861 55567 32919 55573
rect 34514 55564 34520 55616
rect 34572 55604 34578 55616
rect 34885 55607 34943 55613
rect 34885 55604 34897 55607
rect 34572 55576 34897 55604
rect 34572 55564 34578 55576
rect 34885 55573 34897 55576
rect 34931 55573 34943 55607
rect 34885 55567 34943 55573
rect 35526 55564 35532 55616
rect 35584 55604 35590 55616
rect 37844 55604 37872 55644
rect 35584 55576 37872 55604
rect 35584 55564 35590 55576
rect 37918 55564 37924 55616
rect 37976 55604 37982 55616
rect 38746 55604 38752 55616
rect 37976 55576 38752 55604
rect 37976 55564 37982 55576
rect 38746 55564 38752 55576
rect 38804 55564 38810 55616
rect 38856 55604 38884 55644
rect 41785 55641 41797 55675
rect 41831 55641 41843 55675
rect 41785 55635 41843 55641
rect 41509 55607 41567 55613
rect 41509 55604 41521 55607
rect 38856 55576 41521 55604
rect 41509 55573 41521 55576
rect 41555 55573 41567 55607
rect 41800 55604 41828 55635
rect 41874 55632 41880 55684
rect 41932 55672 41938 55684
rect 42076 55672 42104 55703
rect 42150 55700 42156 55752
rect 42208 55740 42214 55752
rect 42628 55740 42656 55780
rect 43438 55749 43444 55752
rect 43395 55743 43444 55749
rect 43395 55740 43407 55743
rect 42208 55712 42253 55740
rect 42628 55712 43407 55740
rect 42208 55700 42214 55712
rect 43395 55709 43407 55712
rect 43441 55709 43444 55743
rect 43395 55703 43444 55709
rect 43438 55700 43444 55703
rect 43496 55740 43502 55752
rect 43640 55749 43668 55836
rect 45462 55808 45468 55820
rect 43824 55780 45468 55808
rect 43824 55749 43852 55780
rect 45462 55768 45468 55780
rect 45520 55768 45526 55820
rect 43625 55743 43683 55749
rect 43496 55712 43543 55740
rect 43496 55700 43502 55712
rect 43625 55709 43637 55743
rect 43671 55709 43683 55743
rect 43625 55703 43683 55709
rect 43808 55743 43866 55749
rect 43808 55709 43820 55743
rect 43854 55709 43866 55743
rect 43808 55703 43866 55709
rect 43898 55700 43904 55752
rect 43956 55740 43962 55752
rect 57701 55743 57759 55749
rect 43956 55712 44001 55740
rect 43956 55700 43962 55712
rect 57701 55709 57713 55743
rect 57747 55740 57759 55743
rect 58342 55740 58348 55752
rect 57747 55712 58348 55740
rect 57747 55709 57759 55712
rect 57701 55703 57759 55709
rect 58342 55700 58348 55712
rect 58400 55700 58406 55752
rect 42886 55672 42892 55684
rect 41932 55644 41977 55672
rect 42076 55644 42892 55672
rect 41932 55632 41938 55644
rect 42886 55632 42892 55644
rect 42944 55632 42950 55684
rect 43533 55675 43591 55681
rect 43533 55641 43545 55675
rect 43579 55641 43591 55675
rect 43533 55635 43591 55641
rect 42702 55604 42708 55616
rect 41800 55576 42708 55604
rect 41509 55567 41567 55573
rect 42702 55564 42708 55576
rect 42760 55564 42766 55616
rect 43254 55604 43260 55616
rect 43215 55576 43260 55604
rect 43254 55564 43260 55576
rect 43312 55564 43318 55616
rect 43548 55604 43576 55635
rect 54570 55604 54576 55616
rect 43548 55576 54576 55604
rect 54570 55564 54576 55576
rect 54628 55564 54634 55616
rect 58161 55607 58219 55613
rect 58161 55573 58173 55607
rect 58207 55604 58219 55607
rect 58526 55604 58532 55616
rect 58207 55576 58532 55604
rect 58207 55573 58219 55576
rect 58161 55567 58219 55573
rect 58526 55564 58532 55576
rect 58584 55564 58590 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 30834 55400 30840 55412
rect 22066 55372 30840 55400
rect 8294 55292 8300 55344
rect 8352 55332 8358 55344
rect 22066 55332 22094 55372
rect 30834 55360 30840 55372
rect 30892 55360 30898 55412
rect 32493 55403 32551 55409
rect 32493 55400 32505 55403
rect 31726 55372 32505 55400
rect 31726 55332 31754 55372
rect 32493 55369 32505 55372
rect 32539 55369 32551 55403
rect 32493 55363 32551 55369
rect 41046 55360 41052 55412
rect 41104 55400 41110 55412
rect 41417 55403 41475 55409
rect 41417 55400 41429 55403
rect 41104 55372 41429 55400
rect 41104 55360 41110 55372
rect 41417 55369 41429 55372
rect 41463 55369 41475 55403
rect 41417 55363 41475 55369
rect 43349 55403 43407 55409
rect 43349 55369 43361 55403
rect 43395 55369 43407 55403
rect 43349 55363 43407 55369
rect 58161 55403 58219 55409
rect 58161 55369 58173 55403
rect 58207 55400 58219 55403
rect 58342 55400 58348 55412
rect 58207 55372 58348 55400
rect 58207 55369 58219 55372
rect 58161 55363 58219 55369
rect 8352 55304 22094 55332
rect 26896 55304 31754 55332
rect 8352 55292 8358 55304
rect 1857 55267 1915 55273
rect 1857 55233 1869 55267
rect 1903 55264 1915 55267
rect 2409 55267 2467 55273
rect 2409 55264 2421 55267
rect 1903 55236 2421 55264
rect 1903 55233 1915 55236
rect 1857 55227 1915 55233
rect 2409 55233 2421 55236
rect 2455 55264 2467 55267
rect 3510 55264 3516 55276
rect 2455 55236 3516 55264
rect 2455 55233 2467 55236
rect 2409 55227 2467 55233
rect 3510 55224 3516 55236
rect 3568 55224 3574 55276
rect 21358 55224 21364 55276
rect 21416 55264 21422 55276
rect 21818 55264 21824 55276
rect 21416 55236 21824 55264
rect 21416 55224 21422 55236
rect 21818 55224 21824 55236
rect 21876 55264 21882 55276
rect 26896 55264 26924 55304
rect 35250 55292 35256 55344
rect 35308 55332 35314 55344
rect 43364 55332 43392 55363
rect 58342 55360 58348 55372
rect 58400 55360 58406 55412
rect 35308 55304 43392 55332
rect 43625 55335 43683 55341
rect 35308 55292 35314 55304
rect 43625 55301 43637 55335
rect 43671 55332 43683 55335
rect 54662 55332 54668 55344
rect 43671 55304 54668 55332
rect 43671 55301 43683 55304
rect 43625 55295 43683 55301
rect 54662 55292 54668 55304
rect 54720 55292 54726 55344
rect 21876 55236 26924 55264
rect 21876 55224 21882 55236
rect 27338 55224 27344 55276
rect 27396 55264 27402 55276
rect 28994 55264 29000 55276
rect 27396 55236 29000 55264
rect 27396 55224 27402 55236
rect 28994 55224 29000 55236
rect 29052 55224 29058 55276
rect 31757 55267 31815 55273
rect 31757 55233 31769 55267
rect 31803 55264 31815 55267
rect 32674 55264 32680 55276
rect 31803 55236 32680 55264
rect 31803 55233 31815 55236
rect 31757 55227 31815 55233
rect 32674 55224 32680 55236
rect 32732 55224 32738 55276
rect 36538 55264 36544 55276
rect 32876 55236 36544 55264
rect 31846 55156 31852 55208
rect 31904 55196 31910 55208
rect 32309 55199 32367 55205
rect 32309 55196 32321 55199
rect 31904 55168 32321 55196
rect 31904 55156 31910 55168
rect 32309 55165 32321 55168
rect 32355 55196 32367 55199
rect 32876 55196 32904 55236
rect 36538 55224 36544 55236
rect 36596 55264 36602 55276
rect 37734 55264 37740 55276
rect 36596 55236 37740 55264
rect 36596 55224 36602 55236
rect 37734 55224 37740 55236
rect 37792 55264 37798 55276
rect 38654 55264 38660 55276
rect 37792 55236 38660 55264
rect 37792 55224 37798 55236
rect 38654 55224 38660 55236
rect 38712 55224 38718 55276
rect 39853 55267 39911 55273
rect 39853 55233 39865 55267
rect 39899 55264 39911 55267
rect 40034 55264 40040 55276
rect 39899 55236 40040 55264
rect 39899 55233 39911 55236
rect 39853 55227 39911 55233
rect 40034 55224 40040 55236
rect 40092 55224 40098 55276
rect 43438 55224 43444 55276
rect 43496 55273 43502 55276
rect 43496 55267 43545 55273
rect 43496 55233 43499 55267
rect 43533 55233 43545 55267
rect 43714 55264 43720 55276
rect 43675 55236 43720 55264
rect 43496 55227 43545 55233
rect 43496 55224 43502 55227
rect 43714 55224 43720 55236
rect 43772 55224 43778 55276
rect 43900 55267 43958 55273
rect 43900 55233 43912 55267
rect 43946 55233 43958 55267
rect 43900 55227 43958 55233
rect 32355 55168 32904 55196
rect 43916 55196 43944 55227
rect 43990 55224 43996 55276
rect 44048 55264 44054 55276
rect 44048 55236 44093 55264
rect 44048 55224 44054 55236
rect 44174 55224 44180 55276
rect 44232 55224 44238 55276
rect 57517 55267 57575 55273
rect 57517 55233 57529 55267
rect 57563 55264 57575 55267
rect 57974 55264 57980 55276
rect 57563 55236 57980 55264
rect 57563 55233 57575 55236
rect 57517 55227 57575 55233
rect 57974 55224 57980 55236
rect 58032 55264 58038 55276
rect 58345 55267 58403 55273
rect 58345 55264 58357 55267
rect 58032 55236 58357 55264
rect 58032 55224 58038 55236
rect 58345 55233 58357 55236
rect 58391 55233 58403 55267
rect 58345 55227 58403 55233
rect 44192 55196 44220 55224
rect 43916 55168 44220 55196
rect 32355 55165 32367 55168
rect 32309 55159 32367 55165
rect 1670 55060 1676 55072
rect 1631 55032 1676 55060
rect 1670 55020 1676 55032
rect 1728 55020 1734 55072
rect 32398 55020 32404 55072
rect 32456 55060 32462 55072
rect 32677 55063 32735 55069
rect 32677 55060 32689 55063
rect 32456 55032 32689 55060
rect 32456 55020 32462 55032
rect 32677 55029 32689 55032
rect 32723 55060 32735 55063
rect 36814 55060 36820 55072
rect 32723 55032 36820 55060
rect 32723 55029 32735 55032
rect 32677 55023 32735 55029
rect 36814 55020 36820 55032
rect 36872 55020 36878 55072
rect 40310 55060 40316 55072
rect 40271 55032 40316 55060
rect 40310 55020 40316 55032
rect 40368 55020 40374 55072
rect 40862 55060 40868 55072
rect 40823 55032 40868 55060
rect 40862 55020 40868 55032
rect 40920 55020 40926 55072
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 24949 54859 25007 54865
rect 24949 54825 24961 54859
rect 24995 54856 25007 54859
rect 25222 54856 25228 54868
rect 24995 54828 25228 54856
rect 24995 54825 25007 54828
rect 24949 54819 25007 54825
rect 25222 54816 25228 54828
rect 25280 54816 25286 54868
rect 40310 54816 40316 54868
rect 40368 54856 40374 54868
rect 40497 54859 40555 54865
rect 40497 54856 40509 54859
rect 40368 54828 40509 54856
rect 40368 54816 40374 54828
rect 40497 54825 40509 54828
rect 40543 54856 40555 54859
rect 41046 54856 41052 54868
rect 40543 54828 41052 54856
rect 40543 54825 40555 54828
rect 40497 54819 40555 54825
rect 41046 54816 41052 54828
rect 41104 54816 41110 54868
rect 41322 54856 41328 54868
rect 41283 54828 41328 54856
rect 41322 54816 41328 54828
rect 41380 54816 41386 54868
rect 41506 54856 41512 54868
rect 41467 54828 41512 54856
rect 41506 54816 41512 54828
rect 41564 54816 41570 54868
rect 33226 54748 33232 54800
rect 33284 54788 33290 54800
rect 40681 54791 40739 54797
rect 33284 54760 35480 54788
rect 33284 54748 33290 54760
rect 25041 54723 25099 54729
rect 25041 54689 25053 54723
rect 25087 54720 25099 54723
rect 25130 54720 25136 54732
rect 25087 54692 25136 54720
rect 25087 54689 25099 54692
rect 25041 54683 25099 54689
rect 25130 54680 25136 54692
rect 25188 54680 25194 54732
rect 27890 54680 27896 54732
rect 27948 54720 27954 54732
rect 34514 54720 34520 54732
rect 27948 54692 34520 54720
rect 27948 54680 27954 54692
rect 34514 54680 34520 54692
rect 34572 54680 34578 54732
rect 21358 54652 21364 54664
rect 21319 54624 21364 54652
rect 21358 54612 21364 54624
rect 21416 54612 21422 54664
rect 24762 54652 24768 54664
rect 24723 54624 24768 54652
rect 24762 54612 24768 54624
rect 24820 54612 24826 54664
rect 32398 54652 32404 54664
rect 32359 54624 32404 54652
rect 32398 54612 32404 54624
rect 32456 54612 32462 54664
rect 35342 54661 35348 54664
rect 35340 54652 35348 54661
rect 35303 54624 35348 54652
rect 35340 54615 35348 54624
rect 35342 54612 35348 54615
rect 35400 54612 35406 54664
rect 35452 54661 35480 54760
rect 40681 54757 40693 54791
rect 40727 54788 40739 54791
rect 42150 54788 42156 54800
rect 40727 54760 42156 54788
rect 40727 54757 40739 54760
rect 40681 54751 40739 54757
rect 42150 54748 42156 54760
rect 42208 54748 42214 54800
rect 35437 54655 35495 54661
rect 35437 54621 35449 54655
rect 35483 54621 35495 54655
rect 35710 54652 35716 54664
rect 35671 54624 35716 54652
rect 35437 54615 35495 54621
rect 35710 54612 35716 54624
rect 35768 54612 35774 54664
rect 35802 54612 35808 54664
rect 35860 54652 35866 54664
rect 35860 54624 35905 54652
rect 35860 54612 35866 54624
rect 40034 54612 40040 54664
rect 40092 54652 40098 54664
rect 40129 54655 40187 54661
rect 40129 54652 40141 54655
rect 40092 54624 40141 54652
rect 40092 54612 40098 54624
rect 40129 54621 40141 54624
rect 40175 54621 40187 54655
rect 43254 54652 43260 54664
rect 40129 54615 40187 54621
rect 40236 54624 43260 54652
rect 20438 54544 20444 54596
rect 20496 54584 20502 54596
rect 21545 54587 21603 54593
rect 21545 54584 21557 54587
rect 20496 54556 21557 54584
rect 20496 54544 20502 54556
rect 21545 54553 21557 54556
rect 21591 54553 21603 54587
rect 21545 54547 21603 54553
rect 25038 54544 25044 54596
rect 25096 54584 25102 54596
rect 35529 54587 35587 54593
rect 25096 54556 35204 54584
rect 25096 54544 25102 54556
rect 21729 54519 21787 54525
rect 21729 54485 21741 54519
rect 21775 54516 21787 54519
rect 23566 54516 23572 54528
rect 21775 54488 23572 54516
rect 21775 54485 21787 54488
rect 21729 54479 21787 54485
rect 23566 54476 23572 54488
rect 23624 54476 23630 54528
rect 24581 54519 24639 54525
rect 24581 54485 24593 54519
rect 24627 54516 24639 54519
rect 25130 54516 25136 54528
rect 24627 54488 25136 54516
rect 24627 54485 24639 54488
rect 24581 54479 24639 54485
rect 25130 54476 25136 54488
rect 25188 54476 25194 54528
rect 32306 54516 32312 54528
rect 32267 54488 32312 54516
rect 32306 54476 32312 54488
rect 32364 54476 32370 54528
rect 32766 54476 32772 54528
rect 32824 54516 32830 54528
rect 35176 54525 35204 54556
rect 35529 54553 35541 54587
rect 35575 54584 35587 54587
rect 40236 54584 40264 54624
rect 43254 54612 43260 54624
rect 43312 54612 43318 54664
rect 40862 54584 40868 54596
rect 35575 54556 40264 54584
rect 40512 54556 40868 54584
rect 35575 54553 35587 54556
rect 35529 54547 35587 54553
rect 32861 54519 32919 54525
rect 32861 54516 32873 54519
rect 32824 54488 32873 54516
rect 32824 54476 32830 54488
rect 32861 54485 32873 54488
rect 32907 54485 32919 54519
rect 32861 54479 32919 54485
rect 35161 54519 35219 54525
rect 35161 54485 35173 54519
rect 35207 54485 35219 54519
rect 35161 54479 35219 54485
rect 36446 54476 36452 54528
rect 36504 54516 36510 54528
rect 37918 54516 37924 54528
rect 36504 54488 37924 54516
rect 36504 54476 36510 54488
rect 37918 54476 37924 54488
rect 37976 54516 37982 54528
rect 38289 54519 38347 54525
rect 38289 54516 38301 54519
rect 37976 54488 38301 54516
rect 37976 54476 37982 54488
rect 38289 54485 38301 54488
rect 38335 54516 38347 54519
rect 38562 54516 38568 54528
rect 38335 54488 38568 54516
rect 38335 54485 38347 54488
rect 38289 54479 38347 54485
rect 38562 54476 38568 54488
rect 38620 54476 38626 54528
rect 39390 54516 39396 54528
rect 39351 54488 39396 54516
rect 39390 54476 39396 54488
rect 39448 54516 39454 54528
rect 40512 54525 40540 54556
rect 40862 54544 40868 54556
rect 40920 54584 40926 54596
rect 41141 54587 41199 54593
rect 41141 54584 41153 54587
rect 40920 54556 41153 54584
rect 40920 54544 40926 54556
rect 41141 54553 41153 54556
rect 41187 54553 41199 54587
rect 41141 54547 41199 54553
rect 40497 54519 40555 54525
rect 40497 54516 40509 54519
rect 39448 54488 40509 54516
rect 39448 54476 39454 54488
rect 40497 54485 40509 54488
rect 40543 54485 40555 54519
rect 40497 54479 40555 54485
rect 41046 54476 41052 54528
rect 41104 54516 41110 54528
rect 41341 54519 41399 54525
rect 41341 54516 41353 54519
rect 41104 54488 41353 54516
rect 41104 54476 41110 54488
rect 41341 54485 41353 54488
rect 41387 54485 41399 54519
rect 58342 54516 58348 54528
rect 58303 54488 58348 54516
rect 41341 54479 41399 54485
rect 58342 54476 58348 54488
rect 58400 54476 58406 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 21910 54272 21916 54324
rect 21968 54312 21974 54324
rect 23017 54315 23075 54321
rect 23017 54312 23029 54315
rect 21968 54284 23029 54312
rect 21968 54272 21974 54284
rect 23017 54281 23029 54284
rect 23063 54281 23075 54315
rect 24673 54315 24731 54321
rect 24673 54312 24685 54315
rect 23017 54275 23075 54281
rect 23768 54284 24685 54312
rect 20714 54204 20720 54256
rect 20772 54244 20778 54256
rect 21269 54247 21327 54253
rect 21269 54244 21281 54247
rect 20772 54216 21281 54244
rect 20772 54204 20778 54216
rect 21269 54213 21281 54216
rect 21315 54213 21327 54247
rect 23032 54244 23060 54275
rect 23768 54253 23796 54284
rect 24673 54281 24685 54284
rect 24719 54281 24731 54315
rect 24673 54275 24731 54281
rect 24762 54272 24768 54324
rect 24820 54312 24826 54324
rect 28258 54312 28264 54324
rect 24820 54284 28264 54312
rect 24820 54272 24826 54284
rect 23753 54247 23811 54253
rect 23032 54216 23704 54244
rect 21269 54207 21327 54213
rect 1857 54179 1915 54185
rect 1857 54145 1869 54179
rect 1903 54176 1915 54179
rect 21085 54179 21143 54185
rect 1903 54148 2452 54176
rect 1903 54145 1915 54148
rect 1857 54139 1915 54145
rect 1670 54040 1676 54052
rect 1631 54012 1676 54040
rect 1670 54000 1676 54012
rect 1728 54000 1734 54052
rect 2424 53981 2452 54148
rect 21085 54145 21097 54179
rect 21131 54176 21143 54179
rect 21358 54176 21364 54188
rect 21131 54148 21364 54176
rect 21131 54145 21143 54148
rect 21085 54139 21143 54145
rect 21358 54136 21364 54148
rect 21416 54136 21422 54188
rect 23566 54176 23572 54188
rect 23527 54148 23572 54176
rect 23566 54136 23572 54148
rect 23624 54136 23630 54188
rect 23676 54176 23704 54216
rect 23753 54213 23765 54247
rect 23799 54213 23811 54247
rect 25038 54244 25044 54256
rect 24999 54216 25044 54244
rect 23753 54207 23811 54213
rect 25038 54204 25044 54216
rect 25096 54204 25102 54256
rect 23845 54179 23903 54185
rect 23845 54176 23857 54179
rect 23676 54148 23857 54176
rect 23845 54145 23857 54148
rect 23891 54145 23903 54179
rect 23845 54139 23903 54145
rect 23934 54136 23940 54188
rect 23992 54185 23998 54188
rect 23992 54179 24047 54185
rect 23992 54145 24001 54179
rect 24035 54176 24047 54179
rect 24670 54176 24676 54188
rect 24035 54148 24676 54176
rect 24035 54145 24047 54148
rect 23992 54139 24047 54145
rect 23992 54136 23998 54139
rect 24670 54136 24676 54148
rect 24728 54136 24734 54188
rect 24854 54185 24860 54188
rect 24852 54176 24860 54185
rect 24815 54148 24860 54176
rect 24852 54139 24860 54148
rect 24854 54136 24860 54139
rect 24912 54136 24918 54188
rect 24949 54179 25007 54185
rect 24949 54145 24961 54179
rect 24995 54145 25007 54179
rect 24949 54139 25007 54145
rect 18874 54068 18880 54120
rect 18932 54108 18938 54120
rect 24964 54108 24992 54139
rect 25130 54136 25136 54188
rect 25188 54185 25194 54188
rect 25188 54179 25227 54185
rect 25215 54145 25227 54179
rect 25188 54139 25227 54145
rect 25317 54179 25375 54185
rect 25317 54145 25329 54179
rect 25363 54176 25375 54179
rect 25590 54176 25596 54188
rect 25363 54148 25596 54176
rect 25363 54145 25375 54148
rect 25317 54139 25375 54145
rect 25188 54136 25194 54139
rect 25590 54136 25596 54148
rect 25648 54136 25654 54188
rect 25976 54176 26004 54284
rect 28258 54272 28264 54284
rect 28316 54272 28322 54324
rect 32306 54272 32312 54324
rect 32364 54312 32370 54324
rect 32686 54315 32744 54321
rect 32686 54312 32698 54315
rect 32364 54284 32698 54312
rect 32364 54272 32370 54284
rect 32686 54281 32698 54284
rect 32732 54281 32744 54315
rect 32686 54275 32744 54281
rect 34532 54284 34928 54312
rect 26418 54204 26424 54256
rect 26476 54244 26482 54256
rect 27433 54247 27491 54253
rect 27433 54244 27445 54247
rect 26476 54216 27445 54244
rect 26476 54204 26482 54216
rect 27433 54213 27445 54216
rect 27479 54213 27491 54247
rect 27433 54207 27491 54213
rect 27525 54247 27583 54253
rect 27525 54213 27537 54247
rect 27571 54244 27583 54247
rect 27890 54244 27896 54256
rect 27571 54216 27896 54244
rect 27571 54213 27583 54216
rect 27525 54207 27583 54213
rect 27890 54204 27896 54216
rect 27948 54204 27954 54256
rect 31573 54247 31631 54253
rect 31573 54213 31585 54247
rect 31619 54213 31631 54247
rect 31573 54207 31631 54213
rect 31757 54247 31815 54253
rect 31757 54213 31769 54247
rect 31803 54244 31815 54247
rect 34532 54244 34560 54284
rect 34900 54253 34928 54284
rect 35710 54272 35716 54324
rect 35768 54312 35774 54324
rect 37461 54315 37519 54321
rect 37461 54312 37473 54315
rect 35768 54284 37473 54312
rect 35768 54272 35774 54284
rect 37461 54281 37473 54284
rect 37507 54281 37519 54315
rect 37461 54275 37519 54281
rect 37734 54272 37740 54324
rect 37792 54312 37798 54324
rect 38841 54315 38899 54321
rect 38841 54312 38853 54315
rect 37792 54284 38853 54312
rect 37792 54272 37798 54284
rect 38841 54281 38853 54284
rect 38887 54281 38899 54315
rect 38841 54275 38899 54281
rect 40773 54315 40831 54321
rect 40773 54281 40785 54315
rect 40819 54312 40831 54315
rect 41874 54312 41880 54324
rect 40819 54284 41880 54312
rect 40819 54281 40831 54284
rect 40773 54275 40831 54281
rect 41874 54272 41880 54284
rect 41932 54272 41938 54324
rect 31803 54216 34560 54244
rect 34885 54247 34943 54253
rect 31803 54213 31815 54216
rect 31757 54207 31815 54213
rect 34655 54213 34713 54219
rect 26329 54179 26387 54185
rect 26329 54176 26341 54179
rect 25976 54148 26341 54176
rect 26329 54145 26341 54148
rect 26375 54145 26387 54179
rect 26329 54139 26387 54145
rect 26605 54179 26663 54185
rect 26605 54145 26617 54179
rect 26651 54176 26663 54179
rect 27154 54176 27160 54188
rect 26651 54148 27160 54176
rect 26651 54145 26663 54148
rect 26605 54139 26663 54145
rect 27154 54136 27160 54148
rect 27212 54136 27218 54188
rect 27338 54185 27344 54188
rect 27336 54176 27344 54185
rect 27299 54148 27344 54176
rect 27336 54139 27344 54148
rect 27338 54136 27344 54139
rect 27396 54136 27402 54188
rect 27653 54179 27711 54185
rect 27653 54176 27665 54179
rect 27448 54148 27665 54176
rect 18932 54080 24992 54108
rect 26145 54111 26203 54117
rect 18932 54068 18938 54080
rect 26145 54077 26157 54111
rect 26191 54108 26203 54111
rect 27448 54108 27476 54148
rect 27653 54145 27665 54148
rect 27699 54145 27711 54179
rect 27653 54139 27711 54145
rect 27801 54179 27859 54185
rect 27801 54145 27813 54179
rect 27847 54176 27859 54179
rect 29086 54176 29092 54188
rect 27847 54148 29092 54176
rect 27847 54145 27859 54148
rect 27801 54139 27859 54145
rect 29086 54136 29092 54148
rect 29144 54176 29150 54188
rect 31297 54179 31355 54185
rect 31297 54176 31309 54179
rect 29144 54148 31309 54176
rect 29144 54136 29150 54148
rect 31297 54145 31309 54148
rect 31343 54145 31355 54179
rect 31588 54176 31616 54207
rect 31846 54176 31852 54188
rect 31588 54148 31852 54176
rect 31297 54139 31355 54145
rect 31846 54136 31852 54148
rect 31904 54136 31910 54188
rect 32309 54179 32367 54185
rect 32309 54145 32321 54179
rect 32355 54176 32367 54179
rect 32766 54176 32772 54188
rect 32355 54148 32772 54176
rect 32355 54145 32367 54148
rect 32309 54139 32367 54145
rect 26191 54080 27476 54108
rect 26191 54077 26203 54080
rect 26145 54071 26203 54077
rect 28626 54068 28632 54120
rect 28684 54108 28690 54120
rect 32324 54108 32352 54139
rect 32766 54136 32772 54148
rect 32824 54136 32830 54188
rect 32950 54176 32956 54188
rect 32911 54148 32956 54176
rect 32950 54136 32956 54148
rect 33008 54136 33014 54188
rect 34655 54179 34667 54213
rect 34701 54179 34713 54213
rect 34885 54213 34897 54247
rect 34931 54244 34943 54247
rect 36722 54244 36728 54256
rect 34931 54216 36728 54244
rect 34931 54213 34943 54216
rect 34885 54207 34943 54213
rect 36722 54204 36728 54216
rect 36780 54204 36786 54256
rect 36814 54204 36820 54256
rect 36872 54244 36878 54256
rect 38654 54244 38660 54256
rect 36872 54216 38660 54244
rect 36872 54204 36878 54216
rect 34655 54176 34713 54179
rect 36446 54176 36452 54188
rect 33980 54148 36452 54176
rect 28684 54080 32352 54108
rect 32784 54108 32812 54136
rect 33980 54117 34008 54148
rect 36446 54136 36452 54148
rect 36504 54136 36510 54188
rect 37642 54176 37648 54188
rect 37603 54148 37648 54176
rect 37642 54136 37648 54148
rect 37700 54136 37706 54188
rect 37734 54136 37740 54188
rect 37792 54176 37798 54188
rect 38028 54185 38056 54216
rect 38654 54204 38660 54216
rect 38712 54204 38718 54256
rect 39390 54204 39396 54256
rect 39448 54244 39454 54256
rect 39669 54247 39727 54253
rect 39669 54244 39681 54247
rect 39448 54216 39681 54244
rect 39448 54204 39454 54216
rect 39669 54213 39681 54216
rect 39715 54244 39727 54247
rect 40589 54247 40647 54253
rect 40589 54244 40601 54247
rect 39715 54216 40601 54244
rect 39715 54213 39727 54216
rect 39669 54207 39727 54213
rect 40589 54213 40601 54216
rect 40635 54213 40647 54247
rect 40589 54207 40647 54213
rect 37921 54179 37979 54185
rect 37792 54148 37837 54176
rect 37792 54136 37798 54148
rect 37921 54145 37933 54179
rect 37967 54145 37979 54179
rect 37921 54139 37979 54145
rect 38013 54179 38071 54185
rect 38013 54145 38025 54179
rect 38059 54145 38071 54179
rect 38562 54176 38568 54188
rect 38523 54148 38568 54176
rect 38013 54139 38071 54145
rect 33965 54111 34023 54117
rect 33965 54108 33977 54111
rect 32784 54080 33977 54108
rect 28684 54068 28690 54080
rect 33965 54077 33977 54080
rect 34011 54077 34023 54111
rect 33965 54071 34023 54077
rect 36722 54068 36728 54120
rect 36780 54108 36786 54120
rect 37936 54108 37964 54139
rect 38562 54136 38568 54148
rect 38620 54176 38626 54188
rect 40221 54179 40279 54185
rect 40221 54176 40233 54179
rect 38620 54148 40233 54176
rect 38620 54136 38626 54148
rect 40221 54145 40233 54148
rect 40267 54176 40279 54179
rect 40310 54176 40316 54188
rect 40267 54148 40316 54176
rect 40267 54145 40279 54148
rect 40221 54139 40279 54145
rect 40310 54136 40316 54148
rect 40368 54136 40374 54188
rect 58342 54176 58348 54188
rect 58303 54148 58348 54176
rect 58342 54136 58348 54148
rect 58400 54136 58406 54188
rect 36780 54080 37964 54108
rect 36780 54068 36786 54080
rect 25222 54000 25228 54052
rect 25280 54040 25286 54052
rect 26513 54043 26571 54049
rect 26513 54040 26525 54043
rect 25280 54012 26525 54040
rect 25280 54000 25286 54012
rect 26513 54009 26525 54012
rect 26559 54040 26571 54043
rect 27338 54040 27344 54052
rect 26559 54012 27344 54040
rect 26559 54009 26571 54012
rect 26513 54003 26571 54009
rect 27338 54000 27344 54012
rect 27396 54000 27402 54052
rect 30466 54000 30472 54052
rect 30524 54040 30530 54052
rect 32306 54040 32312 54052
rect 30524 54012 32312 54040
rect 30524 54000 30530 54012
rect 2409 53975 2467 53981
rect 2409 53941 2421 53975
rect 2455 53972 2467 53975
rect 4798 53972 4804 53984
rect 2455 53944 4804 53972
rect 2455 53941 2467 53944
rect 2409 53935 2467 53941
rect 4798 53932 4804 53944
rect 4856 53932 4862 53984
rect 21453 53975 21511 53981
rect 21453 53941 21465 53975
rect 21499 53972 21511 53975
rect 23382 53972 23388 53984
rect 21499 53944 23388 53972
rect 21499 53941 21511 53944
rect 21453 53935 21511 53941
rect 23382 53932 23388 53944
rect 23440 53932 23446 53984
rect 24118 53972 24124 53984
rect 24079 53944 24124 53972
rect 24118 53932 24124 53944
rect 24176 53932 24182 53984
rect 27062 53932 27068 53984
rect 27120 53972 27126 53984
rect 27157 53975 27215 53981
rect 27157 53972 27169 53975
rect 27120 53944 27169 53972
rect 27120 53932 27126 53944
rect 27157 53941 27169 53944
rect 27203 53941 27215 53975
rect 27157 53935 27215 53941
rect 28994 53932 29000 53984
rect 29052 53972 29058 53984
rect 31588 53981 31616 54012
rect 32306 54000 32312 54012
rect 32364 54000 32370 54052
rect 32398 54000 32404 54052
rect 32456 54040 32462 54052
rect 34517 54043 34575 54049
rect 32456 54012 34468 54040
rect 32456 54000 32462 54012
rect 29549 53975 29607 53981
rect 29549 53972 29561 53975
rect 29052 53944 29561 53972
rect 29052 53932 29058 53944
rect 29549 53941 29561 53944
rect 29595 53941 29607 53975
rect 29549 53935 29607 53941
rect 31573 53975 31631 53981
rect 31573 53941 31585 53975
rect 31619 53941 31631 53975
rect 32674 53972 32680 53984
rect 32635 53944 32680 53972
rect 31573 53935 31631 53941
rect 32674 53932 32680 53944
rect 32732 53972 32738 53984
rect 33413 53975 33471 53981
rect 33413 53972 33425 53975
rect 32732 53944 33425 53972
rect 32732 53932 32738 53944
rect 33413 53941 33425 53944
rect 33459 53941 33471 53975
rect 34440 53972 34468 54012
rect 34517 54009 34529 54043
rect 34563 54040 34575 54043
rect 34606 54040 34612 54052
rect 34563 54012 34612 54040
rect 34563 54009 34575 54012
rect 34517 54003 34575 54009
rect 34606 54000 34612 54012
rect 34664 54040 34670 54052
rect 35802 54040 35808 54052
rect 34664 54012 35808 54040
rect 34664 54000 34670 54012
rect 35802 54000 35808 54012
rect 35860 54000 35866 54052
rect 34701 53975 34759 53981
rect 34701 53972 34713 53975
rect 34440 53944 34713 53972
rect 33413 53935 33471 53941
rect 34701 53941 34713 53944
rect 34747 53941 34759 53975
rect 34701 53935 34759 53941
rect 40034 53932 40040 53984
rect 40092 53972 40098 53984
rect 40589 53975 40647 53981
rect 40589 53972 40601 53975
rect 40092 53944 40601 53972
rect 40092 53932 40098 53944
rect 40589 53941 40601 53944
rect 40635 53972 40647 53975
rect 41233 53975 41291 53981
rect 41233 53972 41245 53975
rect 40635 53944 41245 53972
rect 40635 53941 40647 53944
rect 40589 53935 40647 53941
rect 41233 53941 41245 53944
rect 41279 53972 41291 53975
rect 41322 53972 41328 53984
rect 41279 53944 41328 53972
rect 41279 53941 41291 53944
rect 41233 53935 41291 53941
rect 41322 53932 41328 53944
rect 41380 53932 41386 53984
rect 58161 53975 58219 53981
rect 58161 53941 58173 53975
rect 58207 53972 58219 53975
rect 59170 53972 59176 53984
rect 58207 53944 59176 53972
rect 58207 53941 58219 53944
rect 58161 53935 58219 53941
rect 59170 53932 59176 53944
rect 59228 53932 59234 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 27338 53728 27344 53780
rect 27396 53768 27402 53780
rect 28442 53768 28448 53780
rect 27396 53740 28448 53768
rect 27396 53728 27402 53740
rect 28442 53728 28448 53740
rect 28500 53728 28506 53780
rect 29181 53771 29239 53777
rect 29181 53737 29193 53771
rect 29227 53768 29239 53771
rect 29227 53740 29776 53768
rect 29227 53737 29239 53740
rect 29181 53731 29239 53737
rect 24670 53592 24676 53644
rect 24728 53632 24734 53644
rect 28169 53635 28227 53641
rect 24728 53604 27200 53632
rect 24728 53592 24734 53604
rect 1857 53567 1915 53573
rect 1857 53533 1869 53567
rect 1903 53564 1915 53567
rect 2409 53567 2467 53573
rect 2409 53564 2421 53567
rect 1903 53536 2421 53564
rect 1903 53533 1915 53536
rect 1857 53527 1915 53533
rect 2409 53533 2421 53536
rect 2455 53564 2467 53567
rect 11698 53564 11704 53576
rect 2455 53536 11704 53564
rect 2455 53533 2467 53536
rect 2409 53527 2467 53533
rect 11698 53524 11704 53536
rect 11756 53524 11762 53576
rect 23382 53524 23388 53576
rect 23440 53564 23446 53576
rect 26881 53567 26939 53573
rect 26881 53564 26893 53567
rect 23440 53536 26893 53564
rect 23440 53524 23446 53536
rect 26881 53533 26893 53536
rect 26927 53533 26939 53567
rect 27062 53564 27068 53576
rect 27023 53536 27068 53564
rect 26881 53527 26939 53533
rect 27062 53524 27068 53536
rect 27120 53524 27126 53576
rect 27172 53564 27200 53604
rect 28169 53601 28181 53635
rect 28215 53632 28227 53635
rect 28626 53632 28632 53644
rect 28215 53604 28632 53632
rect 28215 53601 28227 53604
rect 28169 53595 28227 53601
rect 28626 53592 28632 53604
rect 28684 53592 28690 53644
rect 29748 53632 29776 53740
rect 36722 53728 36728 53780
rect 36780 53768 36786 53780
rect 37277 53771 37335 53777
rect 37277 53768 37289 53771
rect 36780 53740 37289 53768
rect 36780 53728 36786 53740
rect 37277 53737 37289 53740
rect 37323 53737 37335 53771
rect 37277 53731 37335 53737
rect 38654 53728 38660 53780
rect 38712 53768 38718 53780
rect 38712 53740 38757 53768
rect 38712 53728 38718 53740
rect 40310 53728 40316 53780
rect 40368 53768 40374 53780
rect 40589 53771 40647 53777
rect 40589 53768 40601 53771
rect 40368 53740 40601 53768
rect 40368 53728 40374 53740
rect 40589 53737 40601 53740
rect 40635 53737 40647 53771
rect 40589 53731 40647 53737
rect 30098 53700 30104 53712
rect 30059 53672 30104 53700
rect 30098 53660 30104 53672
rect 30156 53660 30162 53712
rect 32674 53632 32680 53644
rect 28736 53604 29132 53632
rect 29748 53604 30328 53632
rect 27301 53567 27359 53573
rect 27301 53564 27313 53567
rect 27172 53536 27313 53564
rect 27301 53533 27313 53536
rect 27347 53564 27359 53567
rect 28736 53564 28764 53604
rect 27347 53536 28764 53564
rect 27347 53533 27359 53536
rect 27301 53527 27359 53533
rect 28902 53524 28908 53576
rect 28960 53564 28966 53576
rect 28997 53567 29055 53573
rect 28997 53564 29009 53567
rect 28960 53536 29009 53564
rect 28960 53524 28966 53536
rect 28997 53533 29009 53536
rect 29043 53533 29055 53567
rect 29104 53564 29132 53604
rect 29730 53564 29736 53576
rect 29104 53536 29736 53564
rect 28997 53527 29055 53533
rect 29730 53524 29736 53536
rect 29788 53524 29794 53576
rect 30006 53564 30012 53576
rect 29967 53536 30012 53564
rect 30006 53524 30012 53536
rect 30064 53524 30070 53576
rect 30300 53573 30328 53604
rect 31726 53604 32680 53632
rect 30285 53567 30343 53573
rect 30285 53533 30297 53567
rect 30331 53564 30343 53567
rect 30466 53564 30472 53576
rect 30331 53536 30472 53564
rect 30331 53533 30343 53536
rect 30285 53527 30343 53533
rect 30466 53524 30472 53536
rect 30524 53524 30530 53576
rect 30558 53524 30564 53576
rect 30616 53564 30622 53576
rect 31389 53567 31447 53573
rect 31389 53564 31401 53567
rect 30616 53536 31401 53564
rect 30616 53524 30622 53536
rect 31389 53533 31401 53536
rect 31435 53564 31447 53567
rect 31726 53564 31754 53604
rect 32674 53592 32680 53604
rect 32732 53632 32738 53644
rect 36633 53635 36691 53641
rect 36633 53632 36645 53635
rect 32732 53604 36645 53632
rect 32732 53592 32738 53604
rect 31435 53536 31754 53564
rect 31435 53533 31447 53536
rect 31389 53527 31447 53533
rect 31846 53524 31852 53576
rect 31904 53564 31910 53576
rect 32217 53567 32275 53573
rect 32217 53564 32229 53567
rect 31904 53536 32229 53564
rect 31904 53524 31910 53536
rect 32217 53533 32229 53536
rect 32263 53533 32275 53567
rect 32398 53564 32404 53576
rect 32359 53536 32404 53564
rect 32217 53527 32275 53533
rect 32398 53524 32404 53536
rect 32456 53524 32462 53576
rect 32784 53573 32812 53604
rect 36633 53601 36645 53604
rect 36679 53601 36691 53635
rect 36633 53595 36691 53601
rect 32769 53567 32827 53573
rect 32769 53533 32781 53567
rect 32815 53533 32827 53567
rect 36648 53564 36676 53595
rect 37277 53567 37335 53573
rect 37277 53564 37289 53567
rect 36648 53536 37289 53564
rect 32769 53527 32827 53533
rect 37277 53533 37289 53536
rect 37323 53564 37335 53567
rect 39390 53564 39396 53576
rect 37323 53536 39396 53564
rect 37323 53533 37335 53536
rect 37277 53527 37335 53533
rect 39390 53524 39396 53536
rect 39448 53524 39454 53576
rect 57701 53567 57759 53573
rect 57701 53533 57713 53567
rect 57747 53564 57759 53567
rect 58342 53564 58348 53576
rect 57747 53536 58348 53564
rect 57747 53533 57759 53536
rect 57701 53527 57759 53533
rect 58342 53524 58348 53536
rect 58400 53524 58406 53576
rect 27157 53499 27215 53505
rect 27157 53465 27169 53499
rect 27203 53465 27215 53499
rect 27157 53459 27215 53465
rect 27450 53499 27508 53505
rect 27450 53465 27462 53499
rect 27496 53496 27508 53499
rect 30926 53496 30932 53508
rect 27496 53468 30932 53496
rect 27496 53465 27508 53468
rect 27450 53459 27508 53465
rect 1670 53428 1676 53440
rect 1631 53400 1676 53428
rect 1670 53388 1676 53400
rect 1728 53388 1734 53440
rect 5718 53388 5724 53440
rect 5776 53428 5782 53440
rect 26329 53431 26387 53437
rect 26329 53428 26341 53431
rect 5776 53400 26341 53428
rect 5776 53388 5782 53400
rect 26329 53397 26341 53400
rect 26375 53428 26387 53431
rect 27172 53428 27200 53459
rect 30926 53456 30932 53468
rect 30984 53456 30990 53508
rect 38378 53496 38384 53508
rect 38339 53468 38384 53496
rect 38378 53456 38384 53468
rect 38436 53496 38442 53508
rect 40034 53496 40040 53508
rect 38436 53468 40040 53496
rect 38436 53456 38442 53468
rect 40034 53456 40040 53468
rect 40092 53456 40098 53508
rect 26375 53400 27200 53428
rect 26375 53397 26387 53400
rect 26329 53391 26387 53397
rect 28442 53388 28448 53440
rect 28500 53428 28506 53440
rect 28813 53431 28871 53437
rect 28813 53428 28825 53431
rect 28500 53400 28825 53428
rect 28500 53388 28506 53400
rect 28813 53397 28825 53400
rect 28859 53397 28871 53431
rect 31938 53428 31944 53440
rect 31899 53400 31944 53428
rect 28813 53391 28871 53397
rect 31938 53388 31944 53400
rect 31996 53388 32002 53440
rect 58161 53431 58219 53437
rect 58161 53397 58173 53431
rect 58207 53428 58219 53431
rect 59630 53428 59636 53440
rect 58207 53400 59636 53428
rect 58207 53397 58219 53400
rect 58161 53391 58219 53397
rect 59630 53388 59636 53400
rect 59688 53388 59694 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 28258 53184 28264 53236
rect 28316 53224 28322 53236
rect 29641 53227 29699 53233
rect 29641 53224 29653 53227
rect 28316 53196 29653 53224
rect 28316 53184 28322 53196
rect 29641 53193 29653 53196
rect 29687 53193 29699 53227
rect 29641 53187 29699 53193
rect 29730 53184 29736 53236
rect 29788 53224 29794 53236
rect 30190 53224 30196 53236
rect 29788 53196 30196 53224
rect 29788 53184 29794 53196
rect 30190 53184 30196 53196
rect 30248 53224 30254 53236
rect 31938 53224 31944 53236
rect 30248 53196 31944 53224
rect 30248 53184 30254 53196
rect 31938 53184 31944 53196
rect 31996 53184 32002 53236
rect 30558 53156 30564 53168
rect 29840 53128 30564 53156
rect 28902 53048 28908 53100
rect 28960 53088 28966 53100
rect 29840 53097 29868 53128
rect 30558 53116 30564 53128
rect 30616 53116 30622 53168
rect 29825 53091 29883 53097
rect 29825 53088 29837 53091
rect 28960 53060 29837 53088
rect 28960 53048 28966 53060
rect 29825 53057 29837 53060
rect 29871 53057 29883 53091
rect 30006 53088 30012 53100
rect 29919 53060 30012 53088
rect 29825 53051 29883 53057
rect 30006 53048 30012 53060
rect 30064 53088 30070 53100
rect 31846 53088 31852 53100
rect 30064 53060 31852 53088
rect 30064 53048 30070 53060
rect 31846 53048 31852 53060
rect 31904 53048 31910 53100
rect 27890 52844 27896 52896
rect 27948 52884 27954 52896
rect 28261 52887 28319 52893
rect 28261 52884 28273 52887
rect 27948 52856 28273 52884
rect 27948 52844 27954 52856
rect 28261 52853 28273 52856
rect 28307 52884 28319 52887
rect 28902 52884 28908 52896
rect 28307 52856 28908 52884
rect 28307 52853 28319 52856
rect 28261 52847 28319 52853
rect 28902 52844 28908 52856
rect 28960 52884 28966 52896
rect 28997 52887 29055 52893
rect 28997 52884 29009 52887
rect 28960 52856 29009 52884
rect 28960 52844 28966 52856
rect 28997 52853 29009 52856
rect 29043 52853 29055 52887
rect 28997 52847 29055 52853
rect 30009 52887 30067 52893
rect 30009 52853 30021 52887
rect 30055 52884 30067 52887
rect 30466 52884 30472 52896
rect 30055 52856 30472 52884
rect 30055 52853 30067 52856
rect 30009 52847 30067 52853
rect 30466 52844 30472 52856
rect 30524 52844 30530 52896
rect 38197 52887 38255 52893
rect 38197 52853 38209 52887
rect 38243 52884 38255 52887
rect 38378 52884 38384 52896
rect 38243 52856 38384 52884
rect 38243 52853 38255 52856
rect 38197 52847 38255 52853
rect 38378 52844 38384 52856
rect 38436 52844 38442 52896
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1670 52612 1676 52624
rect 1631 52584 1676 52612
rect 1670 52572 1676 52584
rect 1728 52572 1734 52624
rect 58161 52615 58219 52621
rect 58161 52581 58173 52615
rect 58207 52612 58219 52615
rect 59262 52612 59268 52624
rect 58207 52584 59268 52612
rect 58207 52581 58219 52584
rect 58161 52575 58219 52581
rect 59262 52572 59268 52584
rect 59320 52572 59326 52624
rect 1857 52479 1915 52485
rect 1857 52445 1869 52479
rect 1903 52476 1915 52479
rect 2409 52479 2467 52485
rect 2409 52476 2421 52479
rect 1903 52448 2421 52476
rect 1903 52445 1915 52448
rect 1857 52439 1915 52445
rect 2409 52445 2421 52448
rect 2455 52476 2467 52479
rect 5534 52476 5540 52488
rect 2455 52448 5540 52476
rect 2455 52445 2467 52448
rect 2409 52439 2467 52445
rect 5534 52436 5540 52448
rect 5592 52436 5598 52488
rect 57701 52479 57759 52485
rect 57701 52445 57713 52479
rect 57747 52476 57759 52479
rect 58342 52476 58348 52488
rect 57747 52448 58348 52476
rect 57747 52445 57759 52448
rect 57701 52439 57759 52445
rect 58342 52436 58348 52448
rect 58400 52436 58406 52488
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1857 52003 1915 52009
rect 1857 51969 1869 52003
rect 1903 52000 1915 52003
rect 57517 52003 57575 52009
rect 1903 51972 2452 52000
rect 1903 51969 1915 51972
rect 1857 51963 1915 51969
rect 1670 51796 1676 51808
rect 1631 51768 1676 51796
rect 1670 51756 1676 51768
rect 1728 51756 1734 51808
rect 2424 51805 2452 51972
rect 57517 51969 57529 52003
rect 57563 52000 57575 52003
rect 58342 52000 58348 52012
rect 57563 51972 58348 52000
rect 57563 51969 57575 51972
rect 57517 51963 57575 51969
rect 58342 51960 58348 51972
rect 58400 51960 58406 52012
rect 2409 51799 2467 51805
rect 2409 51765 2421 51799
rect 2455 51796 2467 51799
rect 4890 51796 4896 51808
rect 2455 51768 4896 51796
rect 2455 51765 2467 51768
rect 2409 51759 2467 51765
rect 4890 51756 4896 51768
rect 4948 51756 4954 51808
rect 58161 51799 58219 51805
rect 58161 51765 58173 51799
rect 58207 51796 58219 51799
rect 58986 51796 58992 51808
rect 58207 51768 58992 51796
rect 58207 51765 58219 51768
rect 58161 51759 58219 51765
rect 58986 51756 58992 51768
rect 59044 51756 59050 51808
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 58342 51252 58348 51264
rect 58303 51224 58348 51252
rect 58342 51212 58348 51224
rect 58400 51212 58406 51264
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1857 50915 1915 50921
rect 1857 50881 1869 50915
rect 1903 50912 1915 50915
rect 2409 50915 2467 50921
rect 2409 50912 2421 50915
rect 1903 50884 2421 50912
rect 1903 50881 1915 50884
rect 1857 50875 1915 50881
rect 2409 50881 2421 50884
rect 2455 50912 2467 50915
rect 16574 50912 16580 50924
rect 2455 50884 16580 50912
rect 2455 50881 2467 50884
rect 2409 50875 2467 50881
rect 16574 50872 16580 50884
rect 16632 50872 16638 50924
rect 58342 50912 58348 50924
rect 58303 50884 58348 50912
rect 58342 50872 58348 50884
rect 58400 50872 58406 50924
rect 1670 50776 1676 50788
rect 1631 50748 1676 50776
rect 1670 50736 1676 50748
rect 1728 50736 1734 50788
rect 58161 50711 58219 50717
rect 58161 50677 58173 50711
rect 58207 50708 58219 50711
rect 58894 50708 58900 50720
rect 58207 50680 58900 50708
rect 58207 50677 58219 50680
rect 58161 50671 58219 50677
rect 58894 50668 58900 50680
rect 58952 50668 58958 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 58158 50328 58164 50380
rect 58216 50368 58222 50380
rect 58618 50368 58624 50380
rect 58216 50340 58624 50368
rect 58216 50328 58222 50340
rect 58618 50328 58624 50340
rect 58676 50328 58682 50380
rect 1857 50303 1915 50309
rect 1857 50269 1869 50303
rect 1903 50300 1915 50303
rect 57701 50303 57759 50309
rect 1903 50272 2452 50300
rect 1903 50269 1915 50272
rect 1857 50263 1915 50269
rect 2424 50176 2452 50272
rect 57701 50269 57713 50303
rect 57747 50300 57759 50303
rect 58342 50300 58348 50312
rect 57747 50272 58348 50300
rect 57747 50269 57759 50272
rect 57701 50263 57759 50269
rect 58342 50260 58348 50272
rect 58400 50260 58406 50312
rect 1670 50164 1676 50176
rect 1631 50136 1676 50164
rect 1670 50124 1676 50136
rect 1728 50124 1734 50176
rect 2406 50164 2412 50176
rect 2367 50136 2412 50164
rect 2406 50124 2412 50136
rect 2464 50124 2470 50176
rect 58161 50167 58219 50173
rect 58161 50133 58173 50167
rect 58207 50164 58219 50167
rect 59078 50164 59084 50176
rect 58207 50136 59084 50164
rect 58207 50133 58219 50136
rect 58161 50127 58219 50133
rect 59078 50124 59084 50136
rect 59136 50124 59142 50176
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 2406 49920 2412 49972
rect 2464 49960 2470 49972
rect 13446 49960 13452 49972
rect 2464 49932 13452 49960
rect 2464 49920 2470 49932
rect 13446 49920 13452 49932
rect 13504 49920 13510 49972
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1857 49215 1915 49221
rect 1857 49181 1869 49215
rect 1903 49212 1915 49215
rect 57701 49215 57759 49221
rect 1903 49184 2452 49212
rect 1903 49181 1915 49184
rect 1857 49175 1915 49181
rect 2424 49088 2452 49184
rect 57701 49181 57713 49215
rect 57747 49212 57759 49215
rect 58342 49212 58348 49224
rect 57747 49184 58348 49212
rect 57747 49181 57759 49184
rect 57701 49175 57759 49181
rect 58342 49172 58348 49184
rect 58400 49172 58406 49224
rect 1670 49076 1676 49088
rect 1631 49048 1676 49076
rect 1670 49036 1676 49048
rect 1728 49036 1734 49088
rect 2406 49076 2412 49088
rect 2367 49048 2412 49076
rect 2406 49036 2412 49048
rect 2464 49036 2470 49088
rect 58161 49079 58219 49085
rect 58161 49045 58173 49079
rect 58207 49076 58219 49079
rect 58802 49076 58808 49088
rect 58207 49048 58808 49076
rect 58207 49045 58219 49048
rect 58161 49039 58219 49045
rect 58802 49036 58808 49048
rect 58860 49036 58866 49088
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 2406 48832 2412 48884
rect 2464 48872 2470 48884
rect 13354 48872 13360 48884
rect 2464 48844 13360 48872
rect 2464 48832 2470 48844
rect 13354 48832 13360 48844
rect 13412 48832 13418 48884
rect 1857 48739 1915 48745
rect 1857 48705 1869 48739
rect 1903 48736 1915 48739
rect 2406 48736 2412 48748
rect 1903 48708 2412 48736
rect 1903 48705 1915 48708
rect 1857 48699 1915 48705
rect 2406 48696 2412 48708
rect 2464 48696 2470 48748
rect 57517 48739 57575 48745
rect 57517 48705 57529 48739
rect 57563 48736 57575 48739
rect 58342 48736 58348 48748
rect 57563 48708 58348 48736
rect 57563 48705 57575 48708
rect 57517 48699 57575 48705
rect 58342 48696 58348 48708
rect 58400 48696 58406 48748
rect 1670 48532 1676 48544
rect 1631 48504 1676 48532
rect 1670 48492 1676 48504
rect 1728 48492 1734 48544
rect 2406 48532 2412 48544
rect 2367 48504 2412 48532
rect 2406 48492 2412 48504
rect 2464 48492 2470 48544
rect 58161 48535 58219 48541
rect 58161 48501 58173 48535
rect 58207 48532 58219 48535
rect 59814 48532 59820 48544
rect 58207 48504 59820 48532
rect 58207 48501 58219 48504
rect 58161 48495 58219 48501
rect 59814 48492 59820 48504
rect 59872 48492 59878 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 58342 47988 58348 48000
rect 58303 47960 58348 47988
rect 58342 47948 58348 47960
rect 58400 47948 58406 48000
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1857 47651 1915 47657
rect 1857 47617 1869 47651
rect 1903 47648 1915 47651
rect 58342 47648 58348 47660
rect 1903 47620 2452 47648
rect 58303 47620 58348 47648
rect 1903 47617 1915 47620
rect 1857 47611 1915 47617
rect 1670 47512 1676 47524
rect 1631 47484 1676 47512
rect 1670 47472 1676 47484
rect 1728 47472 1734 47524
rect 2424 47453 2452 47620
rect 58342 47608 58348 47620
rect 58400 47608 58406 47660
rect 5534 47540 5540 47592
rect 5592 47580 5598 47592
rect 17126 47580 17132 47592
rect 5592 47552 17132 47580
rect 5592 47540 5598 47552
rect 17126 47540 17132 47552
rect 17184 47540 17190 47592
rect 2409 47447 2467 47453
rect 2409 47413 2421 47447
rect 2455 47444 2467 47447
rect 9214 47444 9220 47456
rect 2455 47416 9220 47444
rect 2455 47413 2467 47416
rect 2409 47407 2467 47413
rect 9214 47404 9220 47416
rect 9272 47404 9278 47456
rect 55950 47404 55956 47456
rect 56008 47444 56014 47456
rect 58161 47447 58219 47453
rect 58161 47444 58173 47447
rect 56008 47416 58173 47444
rect 56008 47404 56014 47416
rect 58161 47413 58173 47416
rect 58207 47413 58219 47447
rect 58161 47407 58219 47413
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 58161 47175 58219 47181
rect 58161 47141 58173 47175
rect 58207 47172 58219 47175
rect 59538 47172 59544 47184
rect 58207 47144 59544 47172
rect 58207 47141 58219 47144
rect 58161 47135 58219 47141
rect 59538 47132 59544 47144
rect 59596 47132 59602 47184
rect 1857 47039 1915 47045
rect 1857 47005 1869 47039
rect 1903 47036 1915 47039
rect 57701 47039 57759 47045
rect 1903 47008 2452 47036
rect 1903 47005 1915 47008
rect 1857 46999 1915 47005
rect 2424 46977 2452 47008
rect 57701 47005 57713 47039
rect 57747 47036 57759 47039
rect 58342 47036 58348 47048
rect 57747 47008 58348 47036
rect 57747 47005 57759 47008
rect 57701 46999 57759 47005
rect 58342 46996 58348 47008
rect 58400 46996 58406 47048
rect 2409 46971 2467 46977
rect 2409 46937 2421 46971
rect 2455 46968 2467 46971
rect 6638 46968 6644 46980
rect 2455 46940 6644 46968
rect 2455 46937 2467 46940
rect 2409 46931 2467 46937
rect 6638 46928 6644 46940
rect 6696 46928 6702 46980
rect 1670 46900 1676 46912
rect 1631 46872 1676 46900
rect 1670 46860 1676 46872
rect 1728 46860 1734 46912
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 1854 45948 1860 45960
rect 1767 45920 1860 45948
rect 1854 45908 1860 45920
rect 1912 45948 1918 45960
rect 2317 45951 2375 45957
rect 2317 45948 2329 45951
rect 1912 45920 2329 45948
rect 1912 45908 1918 45920
rect 2317 45917 2329 45920
rect 2363 45917 2375 45951
rect 2317 45911 2375 45917
rect 57701 45951 57759 45957
rect 57701 45917 57713 45951
rect 57747 45948 57759 45951
rect 58342 45948 58348 45960
rect 57747 45920 58348 45948
rect 57747 45917 57759 45920
rect 57701 45911 57759 45917
rect 58342 45908 58348 45920
rect 58400 45908 58406 45960
rect 1670 45812 1676 45824
rect 1631 45784 1676 45812
rect 1670 45772 1676 45784
rect 1728 45772 1734 45824
rect 58161 45815 58219 45821
rect 58161 45781 58173 45815
rect 58207 45812 58219 45815
rect 58710 45812 58716 45824
rect 58207 45784 58716 45812
rect 58207 45781 58219 45784
rect 58161 45775 58219 45781
rect 58710 45772 58716 45784
rect 58768 45772 58774 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 3510 45568 3516 45620
rect 3568 45608 3574 45620
rect 7466 45608 7472 45620
rect 3568 45580 7472 45608
rect 3568 45568 3574 45580
rect 7466 45568 7472 45580
rect 7524 45568 7530 45620
rect 1857 45475 1915 45481
rect 1857 45441 1869 45475
rect 1903 45472 1915 45475
rect 57517 45475 57575 45481
rect 1903 45444 2452 45472
rect 1903 45441 1915 45444
rect 1857 45435 1915 45441
rect 1670 45268 1676 45280
rect 1631 45240 1676 45268
rect 1670 45228 1676 45240
rect 1728 45228 1734 45280
rect 2424 45277 2452 45444
rect 57517 45441 57529 45475
rect 57563 45472 57575 45475
rect 58342 45472 58348 45484
rect 57563 45444 58348 45472
rect 57563 45441 57575 45444
rect 57517 45435 57575 45441
rect 58342 45432 58348 45444
rect 58400 45432 58406 45484
rect 2409 45271 2467 45277
rect 2409 45237 2421 45271
rect 2455 45268 2467 45271
rect 9306 45268 9312 45280
rect 2455 45240 9312 45268
rect 2455 45237 2467 45240
rect 2409 45231 2467 45237
rect 9306 45228 9312 45240
rect 9364 45228 9370 45280
rect 57238 45228 57244 45280
rect 57296 45268 57302 45280
rect 58161 45271 58219 45277
rect 58161 45268 58173 45271
rect 57296 45240 58173 45268
rect 57296 45228 57302 45240
rect 58161 45237 58173 45240
rect 58207 45237 58219 45271
rect 58161 45231 58219 45237
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 4890 44820 4896 44872
rect 4948 44860 4954 44872
rect 18782 44860 18788 44872
rect 4948 44832 18788 44860
rect 4948 44820 4954 44832
rect 18782 44820 18788 44832
rect 18840 44820 18846 44872
rect 58342 44724 58348 44736
rect 58303 44696 58348 44724
rect 58342 44684 58348 44696
rect 58400 44684 58406 44736
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1857 44387 1915 44393
rect 1857 44353 1869 44387
rect 1903 44384 1915 44387
rect 1946 44384 1952 44396
rect 1903 44356 1952 44384
rect 1903 44353 1915 44356
rect 1857 44347 1915 44353
rect 1946 44344 1952 44356
rect 2004 44384 2010 44396
rect 2317 44387 2375 44393
rect 2317 44384 2329 44387
rect 2004 44356 2329 44384
rect 2004 44344 2010 44356
rect 2317 44353 2329 44356
rect 2363 44353 2375 44387
rect 58342 44384 58348 44396
rect 58303 44356 58348 44384
rect 2317 44347 2375 44353
rect 58342 44344 58348 44356
rect 58400 44344 58406 44396
rect 57974 44276 57980 44328
rect 58032 44316 58038 44328
rect 58618 44316 58624 44328
rect 58032 44288 58624 44316
rect 58032 44276 58038 44288
rect 58618 44276 58624 44288
rect 58676 44276 58682 44328
rect 1670 44248 1676 44260
rect 1631 44220 1676 44248
rect 1670 44208 1676 44220
rect 1728 44208 1734 44260
rect 58161 44183 58219 44189
rect 58161 44149 58173 44183
rect 58207 44180 58219 44183
rect 58618 44180 58624 44192
rect 58207 44152 58624 44180
rect 58207 44149 58219 44152
rect 58161 44143 58219 44149
rect 58618 44140 58624 44152
rect 58676 44140 58682 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1857 43775 1915 43781
rect 1857 43741 1869 43775
rect 1903 43772 1915 43775
rect 57701 43775 57759 43781
rect 1903 43744 2452 43772
rect 1903 43741 1915 43744
rect 1857 43735 1915 43741
rect 1670 43636 1676 43648
rect 1631 43608 1676 43636
rect 1670 43596 1676 43608
rect 1728 43596 1734 43648
rect 2424 43645 2452 43744
rect 57701 43741 57713 43775
rect 57747 43772 57759 43775
rect 58342 43772 58348 43784
rect 57747 43744 58348 43772
rect 57747 43741 57759 43744
rect 57701 43735 57759 43741
rect 58342 43732 58348 43744
rect 58400 43732 58406 43784
rect 2409 43639 2467 43645
rect 2409 43605 2421 43639
rect 2455 43636 2467 43639
rect 5258 43636 5264 43648
rect 2455 43608 5264 43636
rect 2455 43605 2467 43608
rect 2409 43599 2467 43605
rect 5258 43596 5264 43608
rect 5316 43596 5322 43648
rect 58161 43639 58219 43645
rect 58161 43605 58173 43639
rect 58207 43636 58219 43639
rect 59722 43636 59728 43648
rect 58207 43608 59728 43636
rect 58207 43605 58219 43608
rect 58161 43599 58219 43605
rect 59722 43596 59728 43608
rect 59780 43596 59786 43648
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 1857 42687 1915 42693
rect 1857 42653 1869 42687
rect 1903 42684 1915 42687
rect 57701 42687 57759 42693
rect 1903 42656 2452 42684
rect 1903 42653 1915 42656
rect 1857 42647 1915 42653
rect 1670 42548 1676 42560
rect 1631 42520 1676 42548
rect 1670 42508 1676 42520
rect 1728 42508 1734 42560
rect 2424 42557 2452 42656
rect 57701 42653 57713 42687
rect 57747 42684 57759 42687
rect 58342 42684 58348 42696
rect 57747 42656 58348 42684
rect 57747 42653 57759 42656
rect 57701 42647 57759 42653
rect 58342 42644 58348 42656
rect 58400 42644 58406 42696
rect 2409 42551 2467 42557
rect 2409 42517 2421 42551
rect 2455 42548 2467 42551
rect 6270 42548 6276 42560
rect 2455 42520 6276 42548
rect 2455 42517 2467 42520
rect 2409 42511 2467 42517
rect 6270 42508 6276 42520
rect 6328 42508 6334 42560
rect 56962 42508 56968 42560
rect 57020 42548 57026 42560
rect 58161 42551 58219 42557
rect 58161 42548 58173 42551
rect 57020 42520 58173 42548
rect 57020 42508 57026 42520
rect 58161 42517 58173 42520
rect 58207 42517 58219 42551
rect 58161 42511 58219 42517
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 1857 42211 1915 42217
rect 1857 42177 1869 42211
rect 1903 42208 1915 42211
rect 57517 42211 57575 42217
rect 1903 42180 2452 42208
rect 1903 42177 1915 42180
rect 1857 42171 1915 42177
rect 1670 42004 1676 42016
rect 1631 41976 1676 42004
rect 1670 41964 1676 41976
rect 1728 41964 1734 42016
rect 2424 42013 2452 42180
rect 57517 42177 57529 42211
rect 57563 42208 57575 42211
rect 58342 42208 58348 42220
rect 57563 42180 58348 42208
rect 57563 42177 57575 42180
rect 57517 42171 57575 42177
rect 58342 42168 58348 42180
rect 58400 42168 58406 42220
rect 2409 42007 2467 42013
rect 2409 41973 2421 42007
rect 2455 42004 2467 42007
rect 2498 42004 2504 42016
rect 2455 41976 2504 42004
rect 2455 41973 2467 41976
rect 2409 41967 2467 41973
rect 2498 41964 2504 41976
rect 2556 41964 2562 42016
rect 58161 42007 58219 42013
rect 58161 41973 58173 42007
rect 58207 42004 58219 42007
rect 59446 42004 59452 42016
rect 58207 41976 59452 42004
rect 58207 41973 58219 41976
rect 58161 41967 58219 41973
rect 59446 41964 59452 41976
rect 59504 41964 59510 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 2498 41760 2504 41812
rect 2556 41800 2562 41812
rect 13906 41800 13912 41812
rect 2556 41772 13912 41800
rect 2556 41760 2562 41772
rect 13906 41760 13912 41772
rect 13964 41760 13970 41812
rect 58342 41460 58348 41472
rect 58303 41432 58348 41460
rect 58342 41420 58348 41432
rect 58400 41420 58406 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1857 41123 1915 41129
rect 1857 41089 1869 41123
rect 1903 41120 1915 41123
rect 58342 41120 58348 41132
rect 1903 41092 2452 41120
rect 58303 41092 58348 41120
rect 1903 41089 1915 41092
rect 1857 41083 1915 41089
rect 1670 40984 1676 40996
rect 1631 40956 1676 40984
rect 1670 40944 1676 40956
rect 1728 40944 1734 40996
rect 2424 40925 2452 41092
rect 58342 41080 58348 41092
rect 58400 41080 58406 41132
rect 2409 40919 2467 40925
rect 2409 40885 2421 40919
rect 2455 40916 2467 40919
rect 3510 40916 3516 40928
rect 2455 40888 3516 40916
rect 2455 40885 2467 40888
rect 2409 40879 2467 40885
rect 3510 40876 3516 40888
rect 3568 40876 3574 40928
rect 58158 40916 58164 40928
rect 58119 40888 58164 40916
rect 58158 40876 58164 40888
rect 58216 40876 58222 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 1857 40511 1915 40517
rect 1857 40477 1869 40511
rect 1903 40508 1915 40511
rect 57701 40511 57759 40517
rect 1903 40480 2452 40508
rect 1903 40477 1915 40480
rect 1857 40471 1915 40477
rect 1670 40372 1676 40384
rect 1631 40344 1676 40372
rect 1670 40332 1676 40344
rect 1728 40332 1734 40384
rect 2424 40381 2452 40480
rect 57701 40477 57713 40511
rect 57747 40508 57759 40511
rect 58342 40508 58348 40520
rect 57747 40480 58348 40508
rect 57747 40477 57759 40480
rect 57701 40471 57759 40477
rect 58342 40468 58348 40480
rect 58400 40468 58406 40520
rect 2409 40375 2467 40381
rect 2409 40341 2421 40375
rect 2455 40372 2467 40375
rect 3694 40372 3700 40384
rect 2455 40344 3700 40372
rect 2455 40341 2467 40344
rect 2409 40335 2467 40341
rect 3694 40332 3700 40344
rect 3752 40332 3758 40384
rect 57330 40332 57336 40384
rect 57388 40372 57394 40384
rect 58161 40375 58219 40381
rect 58161 40372 58173 40375
rect 57388 40344 58173 40372
rect 57388 40332 57394 40344
rect 58161 40341 58173 40344
rect 58207 40341 58219 40375
rect 58161 40335 58219 40341
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 3694 40128 3700 40180
rect 3752 40168 3758 40180
rect 11790 40168 11796 40180
rect 3752 40140 11796 40168
rect 3752 40128 3758 40140
rect 11790 40128 11796 40140
rect 11848 40128 11854 40180
rect 57517 39899 57575 39905
rect 57517 39865 57529 39899
rect 57563 39896 57575 39899
rect 58342 39896 58348 39908
rect 57563 39868 58348 39896
rect 57563 39865 57575 39868
rect 57517 39859 57575 39865
rect 58342 39856 58348 39868
rect 58400 39856 58406 39908
rect 57882 39788 57888 39840
rect 57940 39828 57946 39840
rect 58253 39831 58311 39837
rect 58253 39828 58265 39831
rect 57940 39800 58265 39828
rect 57940 39788 57946 39800
rect 58253 39797 58265 39800
rect 58299 39797 58311 39831
rect 58253 39791 58311 39797
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 57609 39627 57667 39633
rect 57609 39593 57621 39627
rect 57655 39624 57667 39627
rect 57974 39624 57980 39636
rect 57655 39596 57980 39624
rect 57655 39593 57667 39596
rect 57609 39587 57667 39593
rect 56686 39448 56692 39500
rect 56744 39448 56750 39500
rect 1857 39423 1915 39429
rect 1857 39389 1869 39423
rect 1903 39420 1915 39423
rect 54941 39423 54999 39429
rect 1903 39392 2452 39420
rect 1903 39389 1915 39392
rect 1857 39383 1915 39389
rect 1670 39284 1676 39296
rect 1631 39256 1676 39284
rect 1670 39244 1676 39256
rect 1728 39244 1734 39296
rect 2424 39293 2452 39392
rect 54941 39389 54953 39423
rect 54987 39420 54999 39423
rect 56226 39420 56232 39432
rect 54987 39392 56232 39420
rect 54987 39389 54999 39392
rect 54941 39383 54999 39389
rect 56226 39380 56232 39392
rect 56284 39420 56290 39432
rect 56505 39423 56563 39429
rect 56505 39420 56517 39423
rect 56284 39392 56517 39420
rect 56284 39380 56290 39392
rect 56505 39389 56517 39392
rect 56551 39389 56563 39423
rect 56505 39383 56563 39389
rect 56597 39423 56655 39429
rect 56597 39389 56609 39423
rect 56643 39420 56655 39423
rect 57624 39420 57652 39587
rect 57974 39584 57980 39596
rect 58032 39584 58038 39636
rect 58342 39420 58348 39432
rect 56643 39392 57652 39420
rect 58303 39392 58348 39420
rect 56643 39389 56655 39392
rect 56597 39383 56655 39389
rect 58342 39380 58348 39392
rect 58400 39380 58406 39432
rect 56134 39352 56140 39364
rect 56095 39324 56140 39352
rect 56134 39312 56140 39324
rect 56192 39312 56198 39364
rect 56873 39355 56931 39361
rect 56873 39321 56885 39355
rect 56919 39352 56931 39355
rect 59814 39352 59820 39364
rect 56919 39324 59820 39352
rect 56919 39321 56931 39324
rect 56873 39315 56931 39321
rect 59814 39312 59820 39324
rect 59872 39312 59878 39364
rect 2409 39287 2467 39293
rect 2409 39253 2421 39287
rect 2455 39284 2467 39287
rect 3418 39284 3424 39296
rect 2455 39256 3424 39284
rect 2455 39253 2467 39256
rect 2409 39247 2467 39253
rect 3418 39244 3424 39256
rect 3476 39244 3482 39296
rect 55585 39287 55643 39293
rect 55585 39253 55597 39287
rect 55631 39284 55643 39287
rect 55674 39284 55680 39296
rect 55631 39256 55680 39284
rect 55631 39253 55643 39256
rect 55585 39247 55643 39253
rect 55674 39244 55680 39256
rect 55732 39244 55738 39296
rect 55769 39287 55827 39293
rect 55769 39253 55781 39287
rect 55815 39284 55827 39287
rect 57422 39284 57428 39296
rect 55815 39256 57428 39284
rect 55815 39253 55827 39256
rect 55769 39247 55827 39253
rect 57422 39244 57428 39256
rect 57480 39244 57486 39296
rect 57606 39244 57612 39296
rect 57664 39284 57670 39296
rect 58161 39287 58219 39293
rect 58161 39284 58173 39287
rect 57664 39256 58173 39284
rect 57664 39244 57670 39256
rect 58161 39253 58173 39256
rect 58207 39253 58219 39287
rect 58161 39247 58219 39253
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 56134 39040 56140 39092
rect 56192 39080 56198 39092
rect 58161 39083 58219 39089
rect 58161 39080 58173 39083
rect 56192 39052 58173 39080
rect 56192 39040 56198 39052
rect 58161 39049 58173 39052
rect 58207 39049 58219 39083
rect 58161 39043 58219 39049
rect 1857 38947 1915 38953
rect 1857 38913 1869 38947
rect 1903 38944 1915 38947
rect 1903 38916 2452 38944
rect 1903 38913 1915 38916
rect 1857 38907 1915 38913
rect 2424 38817 2452 38916
rect 57882 38904 57888 38956
rect 57940 38944 57946 38956
rect 58342 38944 58348 38956
rect 57940 38916 58348 38944
rect 57940 38904 57946 38916
rect 58342 38904 58348 38916
rect 58400 38904 58406 38956
rect 2409 38811 2467 38817
rect 2409 38777 2421 38811
rect 2455 38808 2467 38811
rect 18230 38808 18236 38820
rect 2455 38780 18236 38808
rect 2455 38777 2467 38780
rect 2409 38771 2467 38777
rect 18230 38768 18236 38780
rect 18288 38768 18294 38820
rect 1670 38740 1676 38752
rect 1631 38712 1676 38740
rect 1670 38700 1676 38712
rect 1728 38700 1734 38752
rect 55401 38743 55459 38749
rect 55401 38709 55413 38743
rect 55447 38740 55459 38743
rect 56686 38740 56692 38752
rect 55447 38712 56692 38740
rect 55447 38709 55459 38712
rect 55401 38703 55459 38709
rect 56686 38700 56692 38712
rect 56744 38700 56750 38752
rect 57514 38740 57520 38752
rect 57475 38712 57520 38740
rect 57514 38700 57520 38712
rect 57572 38700 57578 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 55490 38496 55496 38548
rect 55548 38536 55554 38548
rect 56226 38536 56232 38548
rect 55548 38508 56232 38536
rect 55548 38496 55554 38508
rect 56226 38496 56232 38508
rect 56284 38496 56290 38548
rect 56686 38360 56692 38412
rect 56744 38400 56750 38412
rect 56744 38372 57178 38400
rect 56744 38360 56750 38372
rect 57425 38335 57483 38341
rect 57425 38301 57437 38335
rect 57471 38332 57483 38335
rect 57606 38332 57612 38344
rect 57471 38304 57612 38332
rect 57471 38301 57483 38304
rect 57425 38295 57483 38301
rect 57606 38292 57612 38304
rect 57664 38292 57670 38344
rect 57882 38332 57888 38344
rect 57716 38304 57888 38332
rect 55769 38267 55827 38273
rect 55769 38233 55781 38267
rect 55815 38264 55827 38267
rect 57716 38264 57744 38304
rect 57882 38292 57888 38304
rect 57940 38292 57946 38344
rect 58250 38292 58256 38344
rect 58308 38332 58314 38344
rect 59170 38332 59176 38344
rect 58308 38304 59176 38332
rect 58308 38292 58314 38304
rect 59170 38292 59176 38304
rect 59228 38292 59234 38344
rect 55815 38236 57744 38264
rect 57793 38267 57851 38273
rect 55815 38233 55827 38236
rect 55769 38227 55827 38233
rect 57793 38233 57805 38267
rect 57839 38264 57851 38267
rect 57974 38264 57980 38276
rect 57839 38236 57980 38264
rect 57839 38233 57851 38236
rect 57793 38227 57851 38233
rect 57974 38224 57980 38236
rect 58032 38224 58038 38276
rect 58161 38267 58219 38273
rect 58161 38233 58173 38267
rect 58207 38264 58219 38267
rect 58802 38264 58808 38276
rect 58207 38236 58808 38264
rect 58207 38233 58219 38236
rect 58161 38227 58219 38233
rect 58802 38224 58808 38236
rect 58860 38224 58866 38276
rect 56594 38156 56600 38208
rect 56652 38196 56658 38208
rect 56873 38199 56931 38205
rect 56873 38196 56885 38199
rect 56652 38168 56885 38196
rect 56652 38156 56658 38168
rect 56873 38165 56885 38168
rect 56919 38165 56931 38199
rect 56873 38159 56931 38165
rect 57057 38199 57115 38205
rect 57057 38165 57069 38199
rect 57103 38196 57115 38199
rect 59170 38196 59176 38208
rect 57103 38168 59176 38196
rect 57103 38165 57115 38168
rect 57057 38159 57115 38165
rect 59170 38156 59176 38168
rect 59228 38156 59234 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 54757 37995 54815 38001
rect 54757 37961 54769 37995
rect 54803 37992 54815 37995
rect 55766 37992 55772 38004
rect 54803 37964 55772 37992
rect 54803 37961 54815 37964
rect 54757 37955 54815 37961
rect 55766 37952 55772 37964
rect 55824 37952 55830 38004
rect 55861 37995 55919 38001
rect 55861 37961 55873 37995
rect 55907 37992 55919 37995
rect 55950 37992 55956 38004
rect 55907 37964 55956 37992
rect 55907 37961 55919 37964
rect 55861 37955 55919 37961
rect 55950 37952 55956 37964
rect 56008 37952 56014 38004
rect 56597 37995 56655 38001
rect 56597 37961 56609 37995
rect 56643 37992 56655 37995
rect 56778 37992 56784 38004
rect 56643 37964 56784 37992
rect 56643 37961 56655 37964
rect 56597 37955 56655 37961
rect 56778 37952 56784 37964
rect 56836 37952 56842 38004
rect 57517 37995 57575 38001
rect 57517 37961 57529 37995
rect 57563 37992 57575 37995
rect 57882 37992 57888 38004
rect 57563 37964 57888 37992
rect 57563 37961 57575 37964
rect 57517 37955 57575 37961
rect 57882 37952 57888 37964
rect 57940 37992 57946 38004
rect 58066 37992 58072 38004
rect 57940 37964 58072 37992
rect 57940 37952 57946 37964
rect 58066 37952 58072 37964
rect 58124 37952 58130 38004
rect 58161 37995 58219 38001
rect 58161 37961 58173 37995
rect 58207 37961 58219 37995
rect 58161 37955 58219 37961
rect 55125 37927 55183 37933
rect 55125 37893 55137 37927
rect 55171 37924 55183 37927
rect 58176 37924 58204 37955
rect 55171 37896 58204 37924
rect 55171 37893 55183 37896
rect 55125 37887 55183 37893
rect 1857 37859 1915 37865
rect 1857 37825 1869 37859
rect 1903 37856 1915 37859
rect 54021 37859 54079 37865
rect 1903 37828 2452 37856
rect 1903 37825 1915 37828
rect 1857 37819 1915 37825
rect 1670 37720 1676 37732
rect 1631 37692 1676 37720
rect 1670 37680 1676 37692
rect 1728 37680 1734 37732
rect 2424 37661 2452 37828
rect 54021 37825 54033 37859
rect 54067 37856 54079 37859
rect 55490 37856 55496 37868
rect 54067 37828 55496 37856
rect 54067 37825 54079 37828
rect 54021 37819 54079 37825
rect 55490 37816 55496 37828
rect 55548 37816 55554 37868
rect 55585 37859 55643 37865
rect 55585 37825 55597 37859
rect 55631 37856 55643 37859
rect 56778 37856 56784 37868
rect 55631 37828 56784 37856
rect 55631 37825 55643 37828
rect 55585 37819 55643 37825
rect 56778 37816 56784 37828
rect 56836 37816 56842 37868
rect 57514 37816 57520 37868
rect 57572 37856 57578 37868
rect 58342 37856 58348 37868
rect 57572 37828 58348 37856
rect 57572 37816 57578 37828
rect 58342 37816 58348 37828
rect 58400 37816 58406 37868
rect 56686 37788 56692 37800
rect 56074 37760 56692 37788
rect 56686 37748 56692 37760
rect 56744 37748 56750 37800
rect 2409 37655 2467 37661
rect 2409 37621 2421 37655
rect 2455 37652 2467 37655
rect 2590 37652 2596 37664
rect 2455 37624 2596 37652
rect 2455 37621 2467 37624
rect 2409 37615 2467 37621
rect 2590 37612 2596 37624
rect 2648 37612 2654 37664
rect 54573 37655 54631 37661
rect 54573 37621 54585 37655
rect 54619 37652 54631 37655
rect 54662 37652 54668 37664
rect 54619 37624 54668 37652
rect 54619 37621 54631 37624
rect 54573 37615 54631 37621
rect 54662 37612 54668 37624
rect 54720 37612 54726 37664
rect 55858 37612 55864 37664
rect 55916 37652 55922 37664
rect 59814 37652 59820 37664
rect 55916 37624 59820 37652
rect 55916 37612 55922 37624
rect 59814 37612 59820 37624
rect 59872 37612 59878 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 2590 37408 2596 37460
rect 2648 37448 2654 37460
rect 15194 37448 15200 37460
rect 2648 37420 15200 37448
rect 2648 37408 2654 37420
rect 15194 37408 15200 37420
rect 15252 37408 15258 37460
rect 56226 37448 56232 37460
rect 56187 37420 56232 37448
rect 56226 37408 56232 37420
rect 56284 37408 56290 37460
rect 56873 37383 56931 37389
rect 56873 37349 56885 37383
rect 56919 37380 56931 37383
rect 56962 37380 56968 37392
rect 56919 37352 56968 37380
rect 56919 37349 56931 37352
rect 56873 37343 56931 37349
rect 56962 37340 56968 37352
rect 57020 37340 57026 37392
rect 54389 37315 54447 37321
rect 54389 37281 54401 37315
rect 54435 37312 54447 37315
rect 56686 37312 56692 37324
rect 54435 37284 56692 37312
rect 54435 37281 54447 37284
rect 54389 37275 54447 37281
rect 56686 37272 56692 37284
rect 56744 37312 56750 37324
rect 56744 37284 57178 37312
rect 56744 37272 56750 37284
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37244 1915 37247
rect 57882 37244 57888 37256
rect 1903 37216 2452 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 1670 37108 1676 37120
rect 1631 37080 1676 37108
rect 1670 37068 1676 37080
rect 1728 37068 1734 37120
rect 2424 37117 2452 37216
rect 57256 37216 57744 37244
rect 57843 37216 57888 37244
rect 56226 37136 56232 37188
rect 56284 37176 56290 37188
rect 57256 37176 57284 37216
rect 57422 37176 57428 37188
rect 56284 37148 57284 37176
rect 57383 37148 57428 37176
rect 56284 37136 56290 37148
rect 57422 37136 57428 37148
rect 57480 37136 57486 37188
rect 57716 37176 57744 37216
rect 57882 37204 57888 37216
rect 57940 37204 57946 37256
rect 57793 37179 57851 37185
rect 57793 37176 57805 37179
rect 57716 37148 57805 37176
rect 57793 37145 57805 37148
rect 57839 37176 57851 37179
rect 57974 37176 57980 37188
rect 57839 37148 57980 37176
rect 57839 37145 57851 37148
rect 57793 37139 57851 37145
rect 57974 37136 57980 37148
rect 58032 37136 58038 37188
rect 58161 37179 58219 37185
rect 58161 37145 58173 37179
rect 58207 37176 58219 37179
rect 59538 37176 59544 37188
rect 58207 37148 59544 37176
rect 58207 37145 58219 37148
rect 58161 37139 58219 37145
rect 59538 37136 59544 37148
rect 59596 37136 59602 37188
rect 2409 37111 2467 37117
rect 2409 37077 2421 37111
rect 2455 37108 2467 37111
rect 2498 37108 2504 37120
rect 2455 37080 2504 37108
rect 2455 37077 2467 37080
rect 2409 37071 2467 37077
rect 2498 37068 2504 37080
rect 2556 37068 2562 37120
rect 57057 37111 57115 37117
rect 57057 37077 57069 37111
rect 57103 37108 57115 37111
rect 58066 37108 58072 37120
rect 57103 37080 58072 37108
rect 57103 37077 57115 37080
rect 57057 37071 57115 37077
rect 58066 37068 58072 37080
rect 58124 37068 58130 37120
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 56686 36904 56692 36916
rect 56647 36876 56692 36904
rect 56686 36864 56692 36876
rect 56744 36864 56750 36916
rect 57422 36864 57428 36916
rect 57480 36904 57486 36916
rect 58161 36907 58219 36913
rect 58161 36904 58173 36907
rect 57480 36876 58173 36904
rect 57480 36864 57486 36876
rect 58161 36873 58173 36876
rect 58207 36873 58219 36907
rect 58161 36867 58219 36873
rect 57517 36771 57575 36777
rect 57517 36737 57529 36771
rect 57563 36768 57575 36771
rect 58342 36768 58348 36780
rect 57563 36740 58348 36768
rect 57563 36737 57575 36740
rect 57517 36731 57575 36737
rect 58342 36728 58348 36740
rect 58400 36728 58406 36780
rect 58986 36524 58992 36576
rect 59044 36564 59050 36576
rect 59354 36564 59360 36576
rect 59044 36536 59360 36564
rect 59044 36524 59050 36536
rect 59354 36524 59360 36536
rect 59412 36524 59418 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1857 36159 1915 36165
rect 1857 36125 1869 36159
rect 1903 36156 1915 36159
rect 57149 36159 57207 36165
rect 1903 36128 2452 36156
rect 1903 36125 1915 36128
rect 1857 36119 1915 36125
rect 1670 36020 1676 36032
rect 1631 35992 1676 36020
rect 1670 35980 1676 35992
rect 1728 35980 1734 36032
rect 2424 36029 2452 36128
rect 57149 36125 57161 36159
rect 57195 36156 57207 36159
rect 58342 36156 58348 36168
rect 57195 36128 58348 36156
rect 57195 36125 57207 36128
rect 57149 36119 57207 36125
rect 58342 36116 58348 36128
rect 58400 36116 58406 36168
rect 2409 36023 2467 36029
rect 2409 35989 2421 36023
rect 2455 36020 2467 36023
rect 7558 36020 7564 36032
rect 2455 35992 7564 36020
rect 2455 35989 2467 35992
rect 2409 35983 2467 35989
rect 7558 35980 7564 35992
rect 7616 35980 7622 36032
rect 57698 36020 57704 36032
rect 57659 35992 57704 36020
rect 57698 35980 57704 35992
rect 57756 35980 57762 36032
rect 58158 36020 58164 36032
rect 58119 35992 58164 36020
rect 58158 35980 58164 35992
rect 58216 35980 58222 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 56229 35819 56287 35825
rect 56229 35785 56241 35819
rect 56275 35816 56287 35819
rect 56686 35816 56692 35828
rect 56275 35788 56692 35816
rect 56275 35785 56287 35788
rect 56229 35779 56287 35785
rect 56686 35776 56692 35788
rect 56744 35816 56750 35828
rect 57422 35816 57428 35828
rect 56744 35788 57428 35816
rect 56744 35776 56750 35788
rect 57422 35776 57428 35788
rect 57480 35776 57486 35828
rect 57517 35819 57575 35825
rect 57517 35785 57529 35819
rect 57563 35816 57575 35819
rect 57974 35816 57980 35828
rect 57563 35788 57980 35816
rect 57563 35785 57575 35788
rect 57517 35779 57575 35785
rect 57974 35776 57980 35788
rect 58032 35816 58038 35828
rect 58526 35816 58532 35828
rect 58032 35788 58532 35816
rect 58032 35776 58038 35788
rect 58526 35776 58532 35788
rect 58584 35776 58590 35828
rect 1857 35683 1915 35689
rect 1857 35649 1869 35683
rect 1903 35680 1915 35683
rect 2409 35683 2467 35689
rect 2409 35680 2421 35683
rect 1903 35652 2421 35680
rect 1903 35649 1915 35652
rect 1857 35643 1915 35649
rect 2409 35649 2421 35652
rect 2455 35680 2467 35683
rect 7006 35680 7012 35692
rect 2455 35652 7012 35680
rect 2455 35649 2467 35652
rect 2409 35643 2467 35649
rect 7006 35640 7012 35652
rect 7064 35640 7070 35692
rect 57698 35640 57704 35692
rect 57756 35680 57762 35692
rect 58342 35680 58348 35692
rect 57756 35652 58348 35680
rect 57756 35640 57762 35652
rect 58342 35640 58348 35652
rect 58400 35640 58406 35692
rect 1670 35476 1676 35488
rect 1631 35448 1676 35476
rect 1670 35436 1676 35448
rect 1728 35436 1734 35488
rect 57606 35436 57612 35488
rect 57664 35476 57670 35488
rect 58161 35479 58219 35485
rect 58161 35476 58173 35479
rect 57664 35448 58173 35476
rect 57664 35436 57670 35448
rect 58161 35445 58173 35448
rect 58207 35445 58219 35479
rect 58161 35439 58219 35445
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 53926 35232 53932 35284
rect 53984 35272 53990 35284
rect 55861 35275 55919 35281
rect 55861 35272 55873 35275
rect 53984 35244 55873 35272
rect 53984 35232 53990 35244
rect 55861 35241 55873 35244
rect 55907 35272 55919 35275
rect 56226 35272 56232 35284
rect 55907 35244 56232 35272
rect 55907 35241 55919 35244
rect 55861 35235 55919 35241
rect 56226 35232 56232 35244
rect 56284 35232 56290 35284
rect 57146 35232 57152 35284
rect 57204 35272 57210 35284
rect 58710 35272 58716 35284
rect 57204 35244 58716 35272
rect 57204 35232 57210 35244
rect 58710 35232 58716 35244
rect 58768 35232 58774 35284
rect 3510 35164 3516 35216
rect 3568 35204 3574 35216
rect 11238 35204 11244 35216
rect 3568 35176 11244 35204
rect 3568 35164 3574 35176
rect 11238 35164 11244 35176
rect 11296 35164 11302 35216
rect 56244 35136 56272 35232
rect 57974 35204 57980 35216
rect 57440 35176 57980 35204
rect 57146 35145 57152 35148
rect 56965 35139 57023 35145
rect 56965 35136 56977 35139
rect 56244 35108 56977 35136
rect 56965 35105 56977 35108
rect 57011 35105 57023 35139
rect 56965 35099 57023 35105
rect 57124 35139 57152 35145
rect 57124 35105 57136 35139
rect 57124 35099 57152 35105
rect 57146 35096 57152 35099
rect 57204 35096 57210 35148
rect 57241 35139 57299 35145
rect 57241 35105 57253 35139
rect 57287 35136 57299 35139
rect 57440 35136 57468 35176
rect 57974 35164 57980 35176
rect 58032 35164 58038 35216
rect 57287 35108 57468 35136
rect 57287 35105 57299 35108
rect 57241 35099 57299 35105
rect 57514 35096 57520 35148
rect 57572 35136 57578 35148
rect 58158 35136 58164 35148
rect 57572 35108 57617 35136
rect 58119 35108 58164 35136
rect 57572 35096 57578 35108
rect 58158 35096 58164 35108
rect 58216 35096 58222 35148
rect 59078 35096 59084 35148
rect 59136 35096 59142 35148
rect 54570 35068 54576 35080
rect 54531 35040 54576 35068
rect 54570 35028 54576 35040
rect 54628 35028 54634 35080
rect 54754 35028 54760 35080
rect 54812 35068 54818 35080
rect 54849 35071 54907 35077
rect 54849 35068 54861 35071
rect 54812 35040 54861 35068
rect 54812 35028 54818 35040
rect 54849 35037 54861 35040
rect 54895 35037 54907 35071
rect 54849 35031 54907 35037
rect 57977 35071 58035 35077
rect 57977 35037 57989 35071
rect 58023 35068 58035 35071
rect 58802 35068 58808 35080
rect 58023 35040 58808 35068
rect 58023 35037 58035 35040
rect 57977 35031 58035 35037
rect 58802 35028 58808 35040
rect 58860 35028 58866 35080
rect 52362 34960 52368 35012
rect 52420 35000 52426 35012
rect 56321 35003 56379 35009
rect 56321 35000 56333 35003
rect 52420 34972 56333 35000
rect 52420 34960 52426 34972
rect 56321 34969 56333 34972
rect 56367 34969 56379 35003
rect 56321 34963 56379 34969
rect 59096 34944 59124 35096
rect 59078 34892 59084 34944
rect 59136 34892 59142 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 53926 34728 53932 34740
rect 53887 34700 53932 34728
rect 53926 34688 53932 34700
rect 53984 34688 53990 34740
rect 54389 34731 54447 34737
rect 54389 34697 54401 34731
rect 54435 34728 54447 34731
rect 54754 34728 54760 34740
rect 54435 34700 54760 34728
rect 54435 34697 54447 34700
rect 54389 34691 54447 34697
rect 54754 34688 54760 34700
rect 54812 34688 54818 34740
rect 55214 34688 55220 34740
rect 55272 34728 55278 34740
rect 57238 34728 57244 34740
rect 55272 34700 57244 34728
rect 55272 34688 55278 34700
rect 57238 34688 57244 34700
rect 57296 34688 57302 34740
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34561 1915 34595
rect 52362 34592 52368 34604
rect 52323 34564 52368 34592
rect 1857 34555 1915 34561
rect 1872 34524 1900 34555
rect 52362 34552 52368 34564
rect 52420 34552 52426 34604
rect 2409 34527 2467 34533
rect 2409 34524 2421 34527
rect 1872 34496 2421 34524
rect 2409 34493 2421 34496
rect 2455 34524 2467 34527
rect 8202 34524 8208 34536
rect 2455 34496 8208 34524
rect 2455 34493 2467 34496
rect 2409 34487 2467 34493
rect 8202 34484 8208 34496
rect 8260 34484 8266 34536
rect 51442 34484 51448 34536
rect 51500 34524 51506 34536
rect 52089 34527 52147 34533
rect 52089 34524 52101 34527
rect 51500 34496 52101 34524
rect 51500 34484 51506 34496
rect 52089 34493 52101 34496
rect 52135 34493 52147 34527
rect 53944 34524 53972 34688
rect 57606 34660 57612 34672
rect 56244 34632 57612 34660
rect 55214 34601 55220 34604
rect 55192 34595 55220 34601
rect 55192 34561 55204 34595
rect 55192 34555 55220 34561
rect 55214 34552 55220 34555
rect 55272 34552 55278 34604
rect 56244 34601 56272 34632
rect 57606 34620 57612 34632
rect 57664 34620 57670 34672
rect 56229 34595 56287 34601
rect 55876 34564 56180 34592
rect 55033 34527 55091 34533
rect 55033 34524 55045 34527
rect 53944 34496 55045 34524
rect 52089 34487 52147 34493
rect 55033 34493 55045 34496
rect 55079 34493 55091 34527
rect 55033 34487 55091 34493
rect 55309 34527 55367 34533
rect 55309 34493 55321 34527
rect 55355 34524 55367 34527
rect 55876 34524 55904 34564
rect 56042 34524 56048 34536
rect 55355 34496 55904 34524
rect 56003 34496 56048 34524
rect 55355 34493 55367 34496
rect 55309 34487 55367 34493
rect 56042 34484 56048 34496
rect 56100 34484 56106 34536
rect 56152 34524 56180 34564
rect 56229 34561 56241 34595
rect 56275 34561 56287 34595
rect 56229 34555 56287 34561
rect 57517 34595 57575 34601
rect 57517 34561 57529 34595
rect 57563 34592 57575 34595
rect 57882 34592 57888 34604
rect 57563 34564 57888 34592
rect 57563 34561 57575 34564
rect 57517 34555 57575 34561
rect 57882 34552 57888 34564
rect 57940 34592 57946 34604
rect 58161 34595 58219 34601
rect 58161 34592 58173 34595
rect 57940 34564 58173 34592
rect 57940 34552 57946 34564
rect 58161 34561 58173 34564
rect 58207 34561 58219 34595
rect 58161 34555 58219 34561
rect 56781 34527 56839 34533
rect 56781 34524 56793 34527
rect 56152 34496 56793 34524
rect 56781 34493 56793 34496
rect 56827 34524 56839 34527
rect 58434 34524 58440 34536
rect 56827 34496 58440 34524
rect 56827 34493 56839 34496
rect 56781 34487 56839 34493
rect 58434 34484 58440 34496
rect 58492 34484 58498 34536
rect 1670 34456 1676 34468
rect 1631 34428 1676 34456
rect 1670 34416 1676 34428
rect 1728 34416 1734 34468
rect 55582 34416 55588 34468
rect 55640 34456 55646 34468
rect 56686 34456 56692 34468
rect 55640 34428 56692 34456
rect 55640 34416 55646 34428
rect 56686 34416 56692 34428
rect 56744 34416 56750 34468
rect 56962 34416 56968 34468
rect 57020 34456 57026 34468
rect 57514 34456 57520 34468
rect 57020 34428 57520 34456
rect 57020 34416 57026 34428
rect 57514 34416 57520 34428
rect 57572 34416 57578 34468
rect 58342 34388 58348 34400
rect 58303 34360 58348 34388
rect 58342 34348 58348 34360
rect 58400 34348 58406 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 54297 34187 54355 34193
rect 54297 34153 54309 34187
rect 54343 34184 54355 34187
rect 55582 34184 55588 34196
rect 54343 34156 55588 34184
rect 54343 34153 54355 34156
rect 54297 34147 54355 34153
rect 55582 34144 55588 34156
rect 55640 34144 55646 34196
rect 56594 34076 56600 34128
rect 56652 34116 56658 34128
rect 58161 34119 58219 34125
rect 58161 34116 58173 34119
rect 56652 34088 58173 34116
rect 56652 34076 56658 34088
rect 58161 34085 58173 34088
rect 58207 34085 58219 34119
rect 58161 34079 58219 34085
rect 1857 33983 1915 33989
rect 1857 33949 1869 33983
rect 1903 33980 1915 33983
rect 2682 33980 2688 33992
rect 1903 33952 2688 33980
rect 1903 33949 1915 33952
rect 1857 33943 1915 33949
rect 2682 33940 2688 33952
rect 2740 33940 2746 33992
rect 57149 33983 57207 33989
rect 57149 33949 57161 33983
rect 57195 33980 57207 33983
rect 58345 33983 58403 33989
rect 58345 33980 58357 33983
rect 57195 33952 58357 33980
rect 57195 33949 57207 33952
rect 57149 33943 57207 33949
rect 58345 33949 58357 33952
rect 58391 33980 58403 33983
rect 58434 33980 58440 33992
rect 58391 33952 58440 33980
rect 58391 33949 58403 33952
rect 58345 33943 58403 33949
rect 58434 33940 58440 33952
rect 58492 33940 58498 33992
rect 1670 33844 1676 33856
rect 1631 33816 1676 33844
rect 1670 33804 1676 33816
rect 1728 33804 1734 33856
rect 57701 33847 57759 33853
rect 57701 33813 57713 33847
rect 57747 33844 57759 33847
rect 57882 33844 57888 33856
rect 57747 33816 57888 33844
rect 57747 33813 57759 33816
rect 57701 33807 57759 33813
rect 57882 33804 57888 33816
rect 57940 33804 57946 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 56226 33640 56232 33652
rect 56187 33612 56232 33640
rect 56226 33600 56232 33612
rect 56284 33600 56290 33652
rect 56686 33640 56692 33652
rect 56647 33612 56692 33640
rect 56686 33600 56692 33612
rect 56744 33600 56750 33652
rect 57422 33600 57428 33652
rect 57480 33640 57486 33652
rect 57517 33643 57575 33649
rect 57517 33640 57529 33643
rect 57480 33612 57529 33640
rect 57480 33600 57486 33612
rect 57517 33609 57529 33612
rect 57563 33640 57575 33643
rect 58250 33640 58256 33652
rect 57563 33612 58256 33640
rect 57563 33609 57575 33612
rect 57517 33603 57575 33609
rect 58250 33600 58256 33612
rect 58308 33600 58314 33652
rect 57882 33464 57888 33516
rect 57940 33504 57946 33516
rect 58345 33507 58403 33513
rect 58345 33504 58357 33507
rect 57940 33476 58357 33504
rect 57940 33464 57946 33476
rect 58345 33473 58357 33476
rect 58391 33473 58403 33507
rect 58345 33467 58403 33473
rect 57974 33260 57980 33312
rect 58032 33300 58038 33312
rect 58161 33303 58219 33309
rect 58161 33300 58173 33303
rect 58032 33272 58173 33300
rect 58032 33260 58038 33272
rect 58161 33269 58173 33272
rect 58207 33269 58219 33303
rect 58161 33263 58219 33269
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 55861 33099 55919 33105
rect 55861 33065 55873 33099
rect 55907 33096 55919 33099
rect 56134 33096 56140 33108
rect 55907 33068 56140 33096
rect 55907 33065 55919 33068
rect 55861 33059 55919 33065
rect 56134 33056 56140 33068
rect 56192 33096 56198 33108
rect 56686 33096 56692 33108
rect 56192 33068 56692 33096
rect 56192 33056 56198 33068
rect 56686 33056 56692 33068
rect 56744 33096 56750 33108
rect 57698 33096 57704 33108
rect 56744 33068 57704 33096
rect 56744 33056 56750 33068
rect 57698 33056 57704 33068
rect 57756 33056 57762 33108
rect 58618 33028 58624 33040
rect 57624 33000 58624 33028
rect 56226 32920 56232 32972
rect 56284 32960 56290 32972
rect 57149 32963 57207 32969
rect 57149 32960 57161 32963
rect 56284 32932 57161 32960
rect 56284 32920 56290 32932
rect 57149 32929 57161 32932
rect 57195 32929 57207 32963
rect 57149 32923 57207 32929
rect 57308 32963 57366 32969
rect 57308 32929 57320 32963
rect 57354 32960 57366 32963
rect 57624 32960 57652 33000
rect 58618 32988 58624 33000
rect 58676 32988 58682 33040
rect 57354 32932 57652 32960
rect 57354 32929 57366 32932
rect 57308 32923 57366 32929
rect 57698 32920 57704 32972
rect 57756 32960 57762 32972
rect 58342 32960 58348 32972
rect 57756 32932 57801 32960
rect 58303 32932 58348 32960
rect 57756 32920 57762 32932
rect 58342 32920 58348 32932
rect 58400 32920 58406 32972
rect 1857 32895 1915 32901
rect 1857 32861 1869 32895
rect 1903 32892 1915 32895
rect 2222 32892 2228 32904
rect 1903 32864 2228 32892
rect 1903 32861 1915 32864
rect 1857 32855 1915 32861
rect 2222 32852 2228 32864
rect 2280 32852 2286 32904
rect 57422 32892 57428 32904
rect 57383 32864 57428 32892
rect 57422 32852 57428 32864
rect 57480 32852 57486 32904
rect 58161 32895 58219 32901
rect 58161 32861 58173 32895
rect 58207 32892 58219 32895
rect 58618 32892 58624 32904
rect 58207 32864 58624 32892
rect 58207 32861 58219 32864
rect 58161 32855 58219 32861
rect 58618 32852 58624 32864
rect 58676 32852 58682 32904
rect 1670 32756 1676 32768
rect 1631 32728 1676 32756
rect 1670 32716 1676 32728
rect 1728 32716 1734 32768
rect 55858 32716 55864 32768
rect 55916 32756 55922 32768
rect 56505 32759 56563 32765
rect 56505 32756 56517 32759
rect 55916 32728 56517 32756
rect 55916 32716 55922 32728
rect 56505 32725 56517 32728
rect 56551 32725 56563 32759
rect 56505 32719 56563 32725
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 56229 32555 56287 32561
rect 56229 32521 56241 32555
rect 56275 32552 56287 32555
rect 56962 32552 56968 32564
rect 56275 32524 56968 32552
rect 56275 32521 56287 32524
rect 56229 32515 56287 32521
rect 56962 32512 56968 32524
rect 57020 32512 57026 32564
rect 57333 32555 57391 32561
rect 57333 32521 57345 32555
rect 57379 32552 57391 32555
rect 59722 32552 59728 32564
rect 57379 32524 59728 32552
rect 57379 32521 57391 32524
rect 57333 32515 57391 32521
rect 59722 32512 59728 32524
rect 59780 32512 59786 32564
rect 3418 32444 3424 32496
rect 3476 32484 3482 32496
rect 16942 32484 16948 32496
rect 3476 32456 16948 32484
rect 3476 32444 3482 32456
rect 16942 32444 16948 32456
rect 17000 32444 17006 32496
rect 56594 32484 56600 32496
rect 56555 32456 56600 32484
rect 56594 32444 56600 32456
rect 56652 32444 56658 32496
rect 1857 32419 1915 32425
rect 1857 32385 1869 32419
rect 1903 32416 1915 32419
rect 4614 32416 4620 32428
rect 1903 32388 4620 32416
rect 1903 32385 1915 32388
rect 1857 32379 1915 32385
rect 4614 32376 4620 32388
rect 4672 32376 4678 32428
rect 55125 32419 55183 32425
rect 55125 32385 55137 32419
rect 55171 32416 55183 32419
rect 55858 32416 55864 32428
rect 55171 32388 55864 32416
rect 55171 32385 55183 32388
rect 55125 32379 55183 32385
rect 55858 32376 55864 32388
rect 55916 32376 55922 32428
rect 56226 32376 56232 32428
rect 56284 32416 56290 32428
rect 56965 32419 57023 32425
rect 56965 32416 56977 32419
rect 56284 32388 56977 32416
rect 56284 32376 56290 32388
rect 56965 32385 56977 32388
rect 57011 32385 57023 32419
rect 56965 32379 57023 32385
rect 57057 32419 57115 32425
rect 57057 32385 57069 32419
rect 57103 32416 57115 32419
rect 58158 32416 58164 32428
rect 57103 32388 58164 32416
rect 57103 32385 57115 32388
rect 57057 32379 57115 32385
rect 58158 32376 58164 32388
rect 58216 32376 58222 32428
rect 58342 32416 58348 32428
rect 58303 32388 58348 32416
rect 58342 32376 58348 32388
rect 58400 32376 58406 32428
rect 49050 32308 49056 32360
rect 49108 32348 49114 32360
rect 54849 32351 54907 32357
rect 54849 32348 54861 32351
rect 49108 32320 54861 32348
rect 49108 32308 49114 32320
rect 54849 32317 54861 32320
rect 54895 32317 54907 32351
rect 54849 32311 54907 32317
rect 56686 32308 56692 32360
rect 56744 32308 56750 32360
rect 1670 32212 1676 32224
rect 1631 32184 1676 32212
rect 1670 32172 1676 32184
rect 1728 32172 1734 32224
rect 55950 32172 55956 32224
rect 56008 32212 56014 32224
rect 56045 32215 56103 32221
rect 56045 32212 56057 32215
rect 56008 32184 56057 32212
rect 56008 32172 56014 32184
rect 56045 32181 56057 32184
rect 56091 32181 56103 32215
rect 56045 32175 56103 32181
rect 58161 32215 58219 32221
rect 58161 32181 58173 32215
rect 58207 32212 58219 32215
rect 58250 32212 58256 32224
rect 58207 32184 58256 32212
rect 58207 32181 58219 32184
rect 58161 32175 58219 32181
rect 58250 32172 58256 32184
rect 58308 32172 58314 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 55677 32011 55735 32017
rect 55677 31977 55689 32011
rect 55723 32008 55735 32011
rect 56226 32008 56232 32020
rect 55723 31980 56232 32008
rect 55723 31977 55735 31980
rect 55677 31971 55735 31977
rect 56226 31968 56232 31980
rect 56284 31968 56290 32020
rect 58342 32008 58348 32020
rect 58303 31980 58348 32008
rect 58342 31968 58348 31980
rect 58400 31968 58406 32020
rect 57701 31943 57759 31949
rect 57701 31909 57713 31943
rect 57747 31940 57759 31943
rect 58158 31940 58164 31952
rect 57747 31912 58164 31940
rect 57747 31909 57759 31912
rect 57701 31903 57759 31909
rect 58158 31900 58164 31912
rect 58216 31940 58222 31952
rect 59630 31940 59636 31952
rect 58216 31912 59636 31940
rect 58216 31900 58222 31912
rect 59630 31900 59636 31912
rect 59688 31900 59694 31952
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 56965 31467 57023 31473
rect 56965 31433 56977 31467
rect 57011 31464 57023 31467
rect 58434 31464 58440 31476
rect 57011 31436 58440 31464
rect 57011 31433 57023 31436
rect 56965 31427 57023 31433
rect 58434 31424 58440 31436
rect 58492 31464 58498 31476
rect 59262 31464 59268 31476
rect 58492 31436 59268 31464
rect 58492 31424 58498 31436
rect 59262 31424 59268 31436
rect 59320 31424 59326 31476
rect 1857 31331 1915 31337
rect 1857 31297 1869 31331
rect 1903 31328 1915 31331
rect 4062 31328 4068 31340
rect 1903 31300 4068 31328
rect 1903 31297 1915 31300
rect 1857 31291 1915 31297
rect 4062 31288 4068 31300
rect 4120 31288 4126 31340
rect 57517 31331 57575 31337
rect 57517 31297 57529 31331
rect 57563 31328 57575 31331
rect 58158 31328 58164 31340
rect 57563 31300 58164 31328
rect 57563 31297 57575 31300
rect 57517 31291 57575 31297
rect 58158 31288 58164 31300
rect 58216 31288 58222 31340
rect 1670 31192 1676 31204
rect 1631 31164 1676 31192
rect 1670 31152 1676 31164
rect 1728 31152 1734 31204
rect 58342 31124 58348 31136
rect 58303 31096 58348 31124
rect 58342 31084 58348 31096
rect 58400 31084 58406 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 57606 30744 57612 30796
rect 57664 30744 57670 30796
rect 1857 30719 1915 30725
rect 1857 30685 1869 30719
rect 1903 30716 1915 30719
rect 2314 30716 2320 30728
rect 1903 30688 2320 30716
rect 1903 30685 1915 30688
rect 1857 30679 1915 30685
rect 2314 30676 2320 30688
rect 2372 30676 2378 30728
rect 57149 30719 57207 30725
rect 57149 30685 57161 30719
rect 57195 30716 57207 30719
rect 57974 30716 57980 30728
rect 57195 30688 57980 30716
rect 57195 30685 57207 30688
rect 57149 30679 57207 30685
rect 57974 30676 57980 30688
rect 58032 30676 58038 30728
rect 57054 30648 57060 30660
rect 56612 30620 57060 30648
rect 1670 30580 1676 30592
rect 1631 30552 1676 30580
rect 1670 30540 1676 30552
rect 1728 30540 1734 30592
rect 56612 30589 56640 30620
rect 57054 30608 57060 30620
rect 57112 30608 57118 30660
rect 57238 30608 57244 30660
rect 57296 30648 57302 30660
rect 57517 30651 57575 30657
rect 57517 30648 57529 30651
rect 57296 30620 57529 30648
rect 57296 30608 57302 30620
rect 57517 30617 57529 30620
rect 57563 30617 57575 30651
rect 57517 30611 57575 30617
rect 57609 30651 57667 30657
rect 57609 30617 57621 30651
rect 57655 30648 57667 30651
rect 58434 30648 58440 30660
rect 57655 30620 58440 30648
rect 57655 30617 57667 30620
rect 57609 30611 57667 30617
rect 58434 30608 58440 30620
rect 58492 30608 58498 30660
rect 56597 30583 56655 30589
rect 56597 30549 56609 30583
rect 56643 30549 56655 30583
rect 56778 30580 56784 30592
rect 56739 30552 56784 30580
rect 56597 30543 56655 30549
rect 56778 30540 56784 30552
rect 56836 30540 56842 30592
rect 56962 30540 56968 30592
rect 57020 30580 57026 30592
rect 57885 30583 57943 30589
rect 57885 30580 57897 30583
rect 57020 30552 57897 30580
rect 57020 30540 57026 30552
rect 57885 30549 57897 30552
rect 57931 30549 57943 30583
rect 57885 30543 57943 30549
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 56413 30243 56471 30249
rect 56413 30209 56425 30243
rect 56459 30240 56471 30243
rect 58158 30240 58164 30252
rect 56459 30212 58164 30240
rect 56459 30209 56471 30212
rect 56413 30203 56471 30209
rect 58158 30200 58164 30212
rect 58216 30200 58222 30252
rect 56870 30036 56876 30048
rect 56831 30008 56876 30036
rect 56870 29996 56876 30008
rect 56928 30036 56934 30048
rect 57238 30036 57244 30048
rect 56928 30008 57244 30036
rect 56928 29996 56934 30008
rect 57238 29996 57244 30008
rect 57296 29996 57302 30048
rect 57517 30039 57575 30045
rect 57517 30005 57529 30039
rect 57563 30036 57575 30039
rect 57606 30036 57612 30048
rect 57563 30008 57612 30036
rect 57563 30005 57575 30008
rect 57517 29999 57575 30005
rect 57606 29996 57612 30008
rect 57664 29996 57670 30048
rect 58345 30039 58403 30045
rect 58345 30005 58357 30039
rect 58391 30036 58403 30039
rect 58434 30036 58440 30048
rect 58391 30008 58440 30036
rect 58391 30005 58403 30008
rect 58345 29999 58403 30005
rect 58434 29996 58440 30008
rect 58492 29996 58498 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 56870 29656 56876 29708
rect 56928 29696 56934 29708
rect 57057 29699 57115 29705
rect 57057 29696 57069 29699
rect 56928 29668 57069 29696
rect 56928 29656 56934 29668
rect 57057 29665 57069 29668
rect 57103 29665 57115 29699
rect 57514 29696 57520 29708
rect 57057 29659 57115 29665
rect 57348 29668 57520 29696
rect 1857 29631 1915 29637
rect 1857 29597 1869 29631
rect 1903 29628 1915 29631
rect 2409 29631 2467 29637
rect 2409 29628 2421 29631
rect 1903 29600 2421 29628
rect 1903 29597 1915 29600
rect 1857 29591 1915 29597
rect 2409 29597 2421 29600
rect 2455 29628 2467 29631
rect 14642 29628 14648 29640
rect 2455 29600 14648 29628
rect 2455 29597 2467 29600
rect 2409 29591 2467 29597
rect 14642 29588 14648 29600
rect 14700 29588 14706 29640
rect 57238 29637 57244 29640
rect 57195 29631 57244 29637
rect 57195 29597 57207 29631
rect 57241 29597 57244 29631
rect 57195 29591 57244 29597
rect 57238 29588 57244 29591
rect 57296 29588 57302 29640
rect 57348 29637 57376 29668
rect 57514 29656 57520 29668
rect 57572 29656 57578 29708
rect 57606 29656 57612 29708
rect 57664 29696 57670 29708
rect 58250 29696 58256 29708
rect 57664 29668 57709 29696
rect 58211 29668 58256 29696
rect 57664 29656 57670 29668
rect 58250 29656 58256 29668
rect 58308 29656 58314 29708
rect 57333 29631 57391 29637
rect 57333 29597 57345 29631
rect 57379 29597 57391 29631
rect 57333 29591 57391 29597
rect 58069 29631 58127 29637
rect 58069 29597 58081 29631
rect 58115 29628 58127 29631
rect 58710 29628 58716 29640
rect 58115 29600 58716 29628
rect 58115 29597 58127 29600
rect 58069 29591 58127 29597
rect 58710 29588 58716 29600
rect 58768 29588 58774 29640
rect 1670 29492 1676 29504
rect 1631 29464 1676 29492
rect 1670 29452 1676 29464
rect 1728 29452 1734 29504
rect 9950 29492 9956 29504
rect 9911 29464 9956 29492
rect 9950 29452 9956 29464
rect 10008 29452 10014 29504
rect 10597 29495 10655 29501
rect 10597 29461 10609 29495
rect 10643 29492 10655 29495
rect 10686 29492 10692 29504
rect 10643 29464 10692 29492
rect 10643 29461 10655 29464
rect 10597 29455 10655 29461
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 56413 29495 56471 29501
rect 56413 29461 56425 29495
rect 56459 29492 56471 29495
rect 57422 29492 57428 29504
rect 56459 29464 57428 29492
rect 56459 29461 56471 29464
rect 56413 29455 56471 29461
rect 57422 29452 57428 29464
rect 57480 29452 57486 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 3050 29248 3056 29300
rect 3108 29288 3114 29300
rect 9309 29291 9367 29297
rect 9309 29288 9321 29291
rect 3108 29260 9321 29288
rect 3108 29248 3114 29260
rect 9309 29257 9321 29260
rect 9355 29288 9367 29291
rect 9950 29288 9956 29300
rect 9355 29260 9956 29288
rect 9355 29257 9367 29260
rect 9309 29251 9367 29257
rect 9950 29248 9956 29260
rect 10008 29248 10014 29300
rect 10686 29288 10692 29300
rect 10647 29260 10692 29288
rect 10686 29248 10692 29260
rect 10744 29248 10750 29300
rect 58161 29291 58219 29297
rect 58161 29257 58173 29291
rect 58207 29288 58219 29291
rect 58986 29288 58992 29300
rect 58207 29260 58992 29288
rect 58207 29257 58219 29260
rect 58161 29251 58219 29257
rect 58986 29248 58992 29260
rect 59044 29248 59050 29300
rect 10704 29220 10732 29248
rect 9140 29192 10732 29220
rect 56965 29223 57023 29229
rect 1857 29155 1915 29161
rect 1857 29121 1869 29155
rect 1903 29152 1915 29155
rect 6914 29152 6920 29164
rect 1903 29124 2452 29152
rect 6875 29124 6920 29152
rect 1903 29121 1915 29124
rect 1857 29115 1915 29121
rect 1670 29016 1676 29028
rect 1631 28988 1676 29016
rect 1670 28976 1676 28988
rect 1728 28976 1734 29028
rect 2424 29025 2452 29124
rect 6914 29112 6920 29124
rect 6972 29152 6978 29164
rect 8294 29152 8300 29164
rect 6972 29124 8300 29152
rect 6972 29112 6978 29124
rect 8294 29112 8300 29124
rect 8352 29112 8358 29164
rect 7006 29084 7012 29096
rect 6919 29056 7012 29084
rect 7006 29044 7012 29056
rect 7064 29044 7070 29096
rect 7193 29087 7251 29093
rect 7193 29053 7205 29087
rect 7239 29084 7251 29087
rect 7834 29084 7840 29096
rect 7239 29056 7840 29084
rect 7239 29053 7251 29056
rect 7193 29047 7251 29053
rect 7834 29044 7840 29056
rect 7892 29044 7898 29096
rect 9140 29093 9168 29192
rect 56965 29189 56977 29223
rect 57011 29220 57023 29223
rect 57514 29220 57520 29232
rect 57011 29192 57520 29220
rect 57011 29189 57023 29192
rect 56965 29183 57023 29189
rect 57514 29180 57520 29192
rect 57572 29220 57578 29232
rect 59354 29220 59360 29232
rect 57572 29192 59360 29220
rect 57572 29180 57578 29192
rect 59354 29180 59360 29192
rect 59412 29180 59418 29232
rect 57882 29112 57888 29164
rect 57940 29152 57946 29164
rect 58345 29155 58403 29161
rect 58345 29152 58357 29155
rect 57940 29124 58357 29152
rect 57940 29112 57946 29124
rect 58345 29121 58357 29124
rect 58391 29121 58403 29155
rect 58345 29115 58403 29121
rect 9125 29087 9183 29093
rect 9125 29053 9137 29087
rect 9171 29053 9183 29087
rect 9125 29047 9183 29053
rect 9214 29044 9220 29096
rect 9272 29084 9278 29096
rect 9272 29056 9365 29084
rect 9272 29044 9278 29056
rect 57238 29044 57244 29096
rect 57296 29084 57302 29096
rect 59446 29084 59452 29096
rect 57296 29056 59452 29084
rect 57296 29044 57302 29056
rect 59446 29044 59452 29056
rect 59504 29044 59510 29096
rect 2409 29019 2467 29025
rect 2409 28985 2421 29019
rect 2455 29016 2467 29019
rect 6362 29016 6368 29028
rect 2455 28988 6368 29016
rect 2455 28985 2467 28988
rect 2409 28979 2467 28985
rect 6362 28976 6368 28988
rect 6420 28976 6426 29028
rect 7024 29016 7052 29044
rect 7742 29016 7748 29028
rect 7024 28988 7748 29016
rect 7742 28976 7748 28988
rect 7800 28976 7806 29028
rect 9232 29016 9260 29044
rect 10226 29016 10232 29028
rect 9232 28988 10232 29016
rect 10226 28976 10232 28988
rect 10284 28976 10290 29028
rect 57514 29016 57520 29028
rect 57475 28988 57520 29016
rect 57514 28976 57520 28988
rect 57572 28976 57578 29028
rect 6546 28948 6552 28960
rect 6507 28920 6552 28948
rect 6546 28908 6552 28920
rect 6604 28908 6610 28960
rect 9677 28951 9735 28957
rect 9677 28917 9689 28951
rect 9723 28948 9735 28951
rect 10042 28948 10048 28960
rect 9723 28920 10048 28948
rect 9723 28917 9735 28920
rect 9677 28911 9735 28917
rect 10042 28908 10048 28920
rect 10100 28908 10106 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 3602 28704 3608 28756
rect 3660 28744 3666 28756
rect 6914 28744 6920 28756
rect 3660 28716 6920 28744
rect 3660 28704 3666 28716
rect 6914 28704 6920 28716
rect 6972 28704 6978 28756
rect 9950 28704 9956 28756
rect 10008 28744 10014 28756
rect 12437 28747 12495 28753
rect 12437 28744 12449 28747
rect 10008 28716 12449 28744
rect 10008 28704 10014 28716
rect 12437 28713 12449 28716
rect 12483 28744 12495 28747
rect 12483 28716 13400 28744
rect 12483 28713 12495 28716
rect 12437 28707 12495 28713
rect 10505 28611 10563 28617
rect 10505 28577 10517 28611
rect 10551 28608 10563 28611
rect 10686 28608 10692 28620
rect 10551 28580 10692 28608
rect 10551 28577 10563 28580
rect 10505 28571 10563 28577
rect 10686 28568 10692 28580
rect 10744 28568 10750 28620
rect 13173 28611 13231 28617
rect 13173 28577 13185 28611
rect 13219 28608 13231 28611
rect 13219 28580 13308 28608
rect 13219 28577 13231 28580
rect 13173 28571 13231 28577
rect 6546 28540 6552 28552
rect 6507 28512 6552 28540
rect 6546 28500 6552 28512
rect 6604 28500 6610 28552
rect 8294 28500 8300 28552
rect 8352 28540 8358 28552
rect 10229 28543 10287 28549
rect 10229 28540 10241 28543
rect 8352 28512 10241 28540
rect 8352 28500 8358 28512
rect 10229 28509 10241 28512
rect 10275 28540 10287 28543
rect 11609 28543 11667 28549
rect 11609 28540 11621 28543
rect 10275 28512 11621 28540
rect 10275 28509 10287 28512
rect 10229 28503 10287 28509
rect 11609 28509 11621 28512
rect 11655 28509 11667 28543
rect 11609 28503 11667 28509
rect 8202 28432 8208 28484
rect 8260 28472 8266 28484
rect 13280 28472 13308 28580
rect 13372 28549 13400 28716
rect 57790 28704 57796 28756
rect 57848 28744 57854 28756
rect 58161 28747 58219 28753
rect 58161 28744 58173 28747
rect 57848 28716 58173 28744
rect 57848 28704 57854 28716
rect 58161 28713 58173 28716
rect 58207 28713 58219 28747
rect 58161 28707 58219 28713
rect 13722 28676 13728 28688
rect 13683 28648 13728 28676
rect 13722 28636 13728 28648
rect 13780 28636 13786 28688
rect 57149 28679 57207 28685
rect 57149 28645 57161 28679
rect 57195 28676 57207 28679
rect 57882 28676 57888 28688
rect 57195 28648 57888 28676
rect 57195 28645 57207 28648
rect 57149 28639 57207 28645
rect 57882 28636 57888 28648
rect 57940 28636 57946 28688
rect 13357 28543 13415 28549
rect 13357 28509 13369 28543
rect 13403 28509 13415 28543
rect 13814 28540 13820 28552
rect 13357 28503 13415 28509
rect 13464 28512 13820 28540
rect 13464 28472 13492 28512
rect 13814 28500 13820 28512
rect 13872 28500 13878 28552
rect 58342 28540 58348 28552
rect 58303 28512 58348 28540
rect 58342 28500 58348 28512
rect 58400 28500 58406 28552
rect 8260 28444 12434 28472
rect 13280 28444 13492 28472
rect 8260 28432 8266 28444
rect 6454 28364 6460 28416
rect 6512 28404 6518 28416
rect 6733 28407 6791 28413
rect 6733 28404 6745 28407
rect 6512 28376 6745 28404
rect 6512 28364 6518 28376
rect 6733 28373 6745 28376
rect 6779 28373 6791 28407
rect 6733 28367 6791 28373
rect 7469 28407 7527 28413
rect 7469 28373 7481 28407
rect 7515 28404 7527 28407
rect 7834 28404 7840 28416
rect 7515 28376 7840 28404
rect 7515 28373 7527 28376
rect 7469 28367 7527 28373
rect 7834 28364 7840 28376
rect 7892 28364 7898 28416
rect 9858 28404 9864 28416
rect 9819 28376 9864 28404
rect 9858 28364 9864 28376
rect 9916 28364 9922 28416
rect 10318 28404 10324 28416
rect 10279 28376 10324 28404
rect 10318 28364 10324 28376
rect 10376 28404 10382 28416
rect 10870 28404 10876 28416
rect 10376 28376 10876 28404
rect 10376 28364 10382 28376
rect 10870 28364 10876 28376
rect 10928 28404 10934 28416
rect 11057 28407 11115 28413
rect 11057 28404 11069 28407
rect 10928 28376 11069 28404
rect 10928 28364 10934 28376
rect 11057 28373 11069 28376
rect 11103 28373 11115 28407
rect 12406 28404 12434 28444
rect 13265 28407 13323 28413
rect 13265 28404 13277 28407
rect 12406 28376 13277 28404
rect 11057 28367 11115 28373
rect 13265 28373 13277 28376
rect 13311 28404 13323 28407
rect 14277 28407 14335 28413
rect 14277 28404 14289 28407
rect 13311 28376 14289 28404
rect 13311 28373 13323 28376
rect 13265 28367 13323 28373
rect 14277 28373 14289 28376
rect 14323 28404 14335 28407
rect 14366 28404 14372 28416
rect 14323 28376 14372 28404
rect 14323 28373 14335 28376
rect 14277 28367 14335 28373
rect 14366 28364 14372 28376
rect 14424 28364 14430 28416
rect 56870 28364 56876 28416
rect 56928 28404 56934 28416
rect 57146 28404 57152 28416
rect 56928 28376 57152 28404
rect 56928 28364 56934 28376
rect 57146 28364 57152 28376
rect 57204 28404 57210 28416
rect 57609 28407 57667 28413
rect 57609 28404 57621 28407
rect 57204 28376 57621 28404
rect 57204 28364 57210 28376
rect 57609 28373 57621 28376
rect 57655 28373 57667 28407
rect 57609 28367 57667 28373
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 2406 28160 2412 28212
rect 2464 28200 2470 28212
rect 10318 28200 10324 28212
rect 2464 28172 10324 28200
rect 2464 28160 2470 28172
rect 10318 28160 10324 28172
rect 10376 28160 10382 28212
rect 57517 28203 57575 28209
rect 57517 28169 57529 28203
rect 57563 28200 57575 28203
rect 58342 28200 58348 28212
rect 57563 28172 58348 28200
rect 57563 28169 57575 28172
rect 57517 28163 57575 28169
rect 58342 28160 58348 28172
rect 58400 28160 58406 28212
rect 1857 28067 1915 28073
rect 1857 28033 1869 28067
rect 1903 28064 1915 28067
rect 9858 28064 9864 28076
rect 1903 28036 2452 28064
rect 9819 28036 9864 28064
rect 1903 28033 1915 28036
rect 1857 28027 1915 28033
rect 1670 27928 1676 27940
rect 1631 27900 1676 27928
rect 1670 27888 1676 27900
rect 1728 27888 1734 27940
rect 2424 27869 2452 28036
rect 9858 28024 9864 28036
rect 9916 28024 9922 28076
rect 10042 28024 10048 28076
rect 10100 28064 10106 28076
rect 10321 28067 10379 28073
rect 10321 28064 10333 28067
rect 10100 28036 10333 28064
rect 10100 28024 10106 28036
rect 10321 28033 10333 28036
rect 10367 28033 10379 28067
rect 10321 28027 10379 28033
rect 13722 28024 13728 28076
rect 13780 28064 13786 28076
rect 15381 28067 15439 28073
rect 15381 28064 15393 28067
rect 13780 28036 15393 28064
rect 13780 28024 13786 28036
rect 15381 28033 15393 28036
rect 15427 28033 15439 28067
rect 58342 28064 58348 28076
rect 58303 28036 58348 28064
rect 15381 28027 15439 28033
rect 58342 28024 58348 28036
rect 58400 28024 58406 28076
rect 58161 27931 58219 27937
rect 58161 27897 58173 27931
rect 58207 27928 58219 27931
rect 59814 27928 59820 27940
rect 58207 27900 59820 27928
rect 58207 27897 58219 27900
rect 58161 27891 58219 27897
rect 59814 27888 59820 27900
rect 59872 27888 59878 27940
rect 2409 27863 2467 27869
rect 2409 27829 2421 27863
rect 2455 27860 2467 27863
rect 4890 27860 4896 27872
rect 2455 27832 4896 27860
rect 2455 27829 2467 27832
rect 2409 27823 2467 27829
rect 4890 27820 4896 27832
rect 4948 27820 4954 27872
rect 5350 27820 5356 27872
rect 5408 27860 5414 27872
rect 5905 27863 5963 27869
rect 5905 27860 5917 27863
rect 5408 27832 5917 27860
rect 5408 27820 5414 27832
rect 5905 27829 5917 27832
rect 5951 27829 5963 27863
rect 5905 27823 5963 27829
rect 7101 27863 7159 27869
rect 7101 27829 7113 27863
rect 7147 27860 7159 27863
rect 8294 27860 8300 27872
rect 7147 27832 8300 27860
rect 7147 27829 7159 27832
rect 7101 27823 7159 27829
rect 8294 27820 8300 27832
rect 8352 27820 8358 27872
rect 9677 27863 9735 27869
rect 9677 27829 9689 27863
rect 9723 27860 9735 27863
rect 9766 27860 9772 27872
rect 9723 27832 9772 27860
rect 9723 27829 9735 27832
rect 9677 27823 9735 27829
rect 9766 27820 9772 27832
rect 9824 27820 9830 27872
rect 10505 27863 10563 27869
rect 10505 27829 10517 27863
rect 10551 27860 10563 27863
rect 11606 27860 11612 27872
rect 10551 27832 11612 27860
rect 10551 27829 10563 27832
rect 10505 27823 10563 27829
rect 11606 27820 11612 27832
rect 11664 27820 11670 27872
rect 13814 27860 13820 27872
rect 13775 27832 13820 27860
rect 13814 27820 13820 27832
rect 13872 27820 13878 27872
rect 14461 27863 14519 27869
rect 14461 27829 14473 27863
rect 14507 27860 14519 27863
rect 15010 27860 15016 27872
rect 14507 27832 15016 27860
rect 14507 27829 14519 27832
rect 14461 27823 14519 27829
rect 15010 27820 15016 27832
rect 15068 27820 15074 27872
rect 15562 27860 15568 27872
rect 15523 27832 15568 27860
rect 15562 27820 15568 27832
rect 15620 27820 15626 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 5718 27656 5724 27668
rect 5679 27628 5724 27656
rect 5718 27616 5724 27628
rect 5776 27616 5782 27668
rect 6840 27628 7052 27656
rect 2409 27591 2467 27597
rect 2409 27557 2421 27591
rect 2455 27588 2467 27591
rect 6840 27588 6868 27628
rect 2455 27560 6868 27588
rect 6917 27591 6975 27597
rect 2455 27557 2467 27560
rect 2409 27551 2467 27557
rect 6917 27557 6929 27591
rect 6963 27557 6975 27591
rect 6917 27551 6975 27557
rect 1857 27455 1915 27461
rect 1857 27421 1869 27455
rect 1903 27452 1915 27455
rect 2424 27452 2452 27551
rect 5169 27523 5227 27529
rect 5169 27489 5181 27523
rect 5215 27520 5227 27523
rect 6178 27520 6184 27532
rect 5215 27492 6184 27520
rect 5215 27489 5227 27492
rect 5169 27483 5227 27489
rect 6178 27480 6184 27492
rect 6236 27520 6242 27532
rect 6273 27523 6331 27529
rect 6273 27520 6285 27523
rect 6236 27492 6285 27520
rect 6236 27480 6242 27492
rect 6273 27489 6285 27492
rect 6319 27489 6331 27523
rect 6273 27483 6331 27489
rect 5350 27452 5356 27464
rect 1903 27424 2452 27452
rect 5311 27424 5356 27452
rect 1903 27421 1915 27424
rect 1857 27415 1915 27421
rect 5350 27412 5356 27424
rect 5408 27412 5414 27464
rect 5442 27412 5448 27464
rect 5500 27452 5506 27464
rect 6549 27455 6607 27461
rect 6549 27452 6561 27455
rect 5500 27424 6561 27452
rect 5500 27412 5506 27424
rect 6549 27421 6561 27424
rect 6595 27421 6607 27455
rect 6932 27452 6960 27551
rect 7024 27520 7052 27628
rect 9490 27616 9496 27668
rect 9548 27656 9554 27668
rect 10505 27659 10563 27665
rect 10505 27656 10517 27659
rect 9548 27628 10517 27656
rect 9548 27616 9554 27628
rect 10505 27625 10517 27628
rect 10551 27656 10563 27659
rect 10686 27656 10692 27668
rect 10551 27628 10692 27656
rect 10551 27625 10563 27628
rect 10505 27619 10563 27625
rect 10686 27616 10692 27628
rect 10744 27616 10750 27668
rect 58342 27656 58348 27668
rect 57716 27628 58348 27656
rect 7561 27591 7619 27597
rect 7561 27557 7573 27591
rect 7607 27588 7619 27591
rect 8110 27588 8116 27600
rect 7607 27560 8116 27588
rect 7607 27557 7619 27560
rect 7561 27551 7619 27557
rect 8110 27548 8116 27560
rect 8168 27548 8174 27600
rect 7650 27520 7656 27532
rect 7024 27492 7656 27520
rect 7650 27480 7656 27492
rect 7708 27480 7714 27532
rect 7377 27455 7435 27461
rect 7377 27452 7389 27455
rect 6932 27424 7389 27452
rect 6549 27415 6607 27421
rect 7377 27421 7389 27424
rect 7423 27421 7435 27455
rect 10704 27452 10732 27616
rect 14182 27588 14188 27600
rect 13372 27560 14188 27588
rect 13372 27532 13400 27560
rect 14182 27548 14188 27560
rect 14240 27588 14246 27600
rect 57716 27597 57744 27628
rect 58342 27616 58348 27628
rect 58400 27616 58406 27668
rect 14277 27591 14335 27597
rect 14277 27588 14289 27591
rect 14240 27560 14289 27588
rect 14240 27548 14246 27560
rect 14277 27557 14289 27560
rect 14323 27557 14335 27591
rect 14277 27551 14335 27557
rect 57701 27591 57759 27597
rect 57701 27557 57713 27591
rect 57747 27557 57759 27591
rect 57701 27551 57759 27557
rect 58066 27548 58072 27600
rect 58124 27588 58130 27600
rect 58161 27591 58219 27597
rect 58161 27588 58173 27591
rect 58124 27560 58173 27588
rect 58124 27548 58130 27560
rect 58161 27557 58173 27560
rect 58207 27557 58219 27591
rect 58161 27551 58219 27557
rect 13354 27520 13360 27532
rect 13315 27492 13360 27520
rect 13354 27480 13360 27492
rect 13412 27480 13418 27532
rect 13541 27523 13599 27529
rect 13541 27489 13553 27523
rect 13587 27520 13599 27523
rect 13998 27520 14004 27532
rect 13587 27492 14004 27520
rect 13587 27489 13599 27492
rect 13541 27483 13599 27489
rect 13556 27452 13584 27483
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 57149 27523 57207 27529
rect 57149 27489 57161 27523
rect 57195 27520 57207 27523
rect 57974 27520 57980 27532
rect 57195 27492 57980 27520
rect 57195 27489 57207 27492
rect 57149 27483 57207 27489
rect 57974 27480 57980 27492
rect 58032 27520 58038 27532
rect 59078 27520 59084 27532
rect 58032 27492 59084 27520
rect 58032 27480 58038 27492
rect 59078 27480 59084 27492
rect 59136 27480 59142 27532
rect 58342 27452 58348 27464
rect 10704 27424 13584 27452
rect 58303 27424 58348 27452
rect 7377 27415 7435 27421
rect 58342 27412 58348 27424
rect 58400 27412 58406 27464
rect 5258 27384 5264 27396
rect 5171 27356 5264 27384
rect 5258 27344 5264 27356
rect 5316 27384 5322 27396
rect 5902 27384 5908 27396
rect 5316 27356 5908 27384
rect 5316 27344 5322 27356
rect 5902 27344 5908 27356
rect 5960 27344 5966 27396
rect 7834 27344 7840 27396
rect 7892 27384 7898 27396
rect 10594 27384 10600 27396
rect 7892 27356 10600 27384
rect 7892 27344 7898 27356
rect 10594 27344 10600 27356
rect 10652 27344 10658 27396
rect 10778 27344 10784 27396
rect 10836 27384 10842 27396
rect 12161 27387 12219 27393
rect 12161 27384 12173 27387
rect 10836 27356 12173 27384
rect 10836 27344 10842 27356
rect 12161 27353 12173 27356
rect 12207 27384 12219 27387
rect 12207 27356 13308 27384
rect 12207 27353 12219 27356
rect 12161 27347 12219 27353
rect 1670 27316 1676 27328
rect 1631 27288 1676 27316
rect 1670 27276 1676 27288
rect 1728 27276 1734 27328
rect 1946 27276 1952 27328
rect 2004 27316 2010 27328
rect 6457 27319 6515 27325
rect 6457 27316 6469 27319
rect 2004 27288 6469 27316
rect 2004 27276 2010 27288
rect 6457 27285 6469 27288
rect 6503 27316 6515 27319
rect 8113 27319 8171 27325
rect 8113 27316 8125 27319
rect 6503 27288 8125 27316
rect 6503 27285 6515 27288
rect 6457 27279 6515 27285
rect 8113 27285 8125 27288
rect 8159 27316 8171 27319
rect 8754 27316 8760 27328
rect 8159 27288 8760 27316
rect 8159 27285 8171 27288
rect 8113 27279 8171 27285
rect 8754 27276 8760 27288
rect 8812 27276 8818 27328
rect 9214 27276 9220 27328
rect 9272 27316 9278 27328
rect 9861 27319 9919 27325
rect 9861 27316 9873 27319
rect 9272 27288 9873 27316
rect 9272 27276 9278 27288
rect 9861 27285 9873 27288
rect 9907 27285 9919 27319
rect 9861 27279 9919 27285
rect 11514 27276 11520 27328
rect 11572 27316 11578 27328
rect 11609 27319 11667 27325
rect 11609 27316 11621 27319
rect 11572 27288 11621 27316
rect 11572 27276 11578 27288
rect 11609 27285 11621 27288
rect 11655 27285 11667 27319
rect 11609 27279 11667 27285
rect 12342 27276 12348 27328
rect 12400 27316 12406 27328
rect 13280 27325 13308 27356
rect 12897 27319 12955 27325
rect 12897 27316 12909 27319
rect 12400 27288 12909 27316
rect 12400 27276 12406 27288
rect 12897 27285 12909 27288
rect 12943 27285 12955 27319
rect 12897 27279 12955 27285
rect 13265 27319 13323 27325
rect 13265 27285 13277 27319
rect 13311 27316 13323 27319
rect 14829 27319 14887 27325
rect 14829 27316 14841 27319
rect 13311 27288 14841 27316
rect 13311 27285 13323 27288
rect 13265 27279 13323 27285
rect 14829 27285 14841 27288
rect 14875 27285 14887 27319
rect 14829 27279 14887 27285
rect 15010 27276 15016 27328
rect 15068 27316 15074 27328
rect 15381 27319 15439 27325
rect 15381 27316 15393 27319
rect 15068 27288 15393 27316
rect 15068 27276 15074 27288
rect 15381 27285 15393 27288
rect 15427 27285 15439 27319
rect 15381 27279 15439 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 5445 27115 5503 27121
rect 5445 27081 5457 27115
rect 5491 27112 5503 27115
rect 6178 27112 6184 27124
rect 5491 27084 6184 27112
rect 5491 27081 5503 27084
rect 5445 27075 5503 27081
rect 6178 27072 6184 27084
rect 6236 27072 6242 27124
rect 8849 27115 8907 27121
rect 8849 27081 8861 27115
rect 8895 27081 8907 27115
rect 9306 27112 9312 27124
rect 9267 27084 9312 27112
rect 8849 27075 8907 27081
rect 3970 27004 3976 27056
rect 4028 27044 4034 27056
rect 4341 27047 4399 27053
rect 4341 27044 4353 27047
rect 4028 27016 4353 27044
rect 4028 27004 4034 27016
rect 4341 27013 4353 27016
rect 4387 27044 4399 27047
rect 7834 27044 7840 27056
rect 4387 27016 7840 27044
rect 4387 27013 4399 27016
rect 4341 27007 4399 27013
rect 7834 27004 7840 27016
rect 7892 27004 7898 27056
rect 2590 26936 2596 26988
rect 2648 26976 2654 26988
rect 2648 26948 3832 26976
rect 2648 26936 2654 26948
rect 2498 26868 2504 26920
rect 2556 26908 2562 26920
rect 3804 26917 3832 26948
rect 5718 26936 5724 26988
rect 5776 26976 5782 26988
rect 6549 26979 6607 26985
rect 6549 26976 6561 26979
rect 5776 26948 6561 26976
rect 5776 26936 5782 26948
rect 6549 26945 6561 26948
rect 6595 26945 6607 26979
rect 6549 26939 6607 26945
rect 8205 26979 8263 26985
rect 8205 26945 8217 26979
rect 8251 26976 8263 26979
rect 8864 26976 8892 27075
rect 9306 27072 9312 27084
rect 9364 27072 9370 27124
rect 11149 27115 11207 27121
rect 11149 27081 11161 27115
rect 11195 27081 11207 27115
rect 11149 27075 11207 27081
rect 9214 27044 9220 27056
rect 9175 27016 9220 27044
rect 9214 27004 9220 27016
rect 9272 27004 9278 27056
rect 8251 26948 8892 26976
rect 8251 26945 8263 26948
rect 8205 26939 8263 26945
rect 3789 26911 3847 26917
rect 2556 26880 2774 26908
rect 2556 26868 2562 26880
rect 2746 26840 2774 26880
rect 3789 26877 3801 26911
rect 3835 26908 3847 26911
rect 9232 26908 9260 27004
rect 10318 26936 10324 26988
rect 10376 26976 10382 26988
rect 10778 26976 10784 26988
rect 10376 26948 10784 26976
rect 10376 26936 10382 26948
rect 10778 26936 10784 26948
rect 10836 26936 10842 26988
rect 11164 26976 11192 27075
rect 12066 27072 12072 27124
rect 12124 27112 12130 27124
rect 14553 27115 14611 27121
rect 14553 27112 14565 27115
rect 12124 27084 14565 27112
rect 12124 27072 12130 27084
rect 14553 27081 14565 27084
rect 14599 27081 14611 27115
rect 58342 27112 58348 27124
rect 58303 27084 58348 27112
rect 14553 27075 14611 27081
rect 58342 27072 58348 27084
rect 58400 27072 58406 27124
rect 13446 27044 13452 27056
rect 13407 27016 13452 27044
rect 13446 27004 13452 27016
rect 13504 27004 13510 27056
rect 13814 27004 13820 27056
rect 13872 27044 13878 27056
rect 15102 27044 15108 27056
rect 13872 27016 15108 27044
rect 13872 27004 13878 27016
rect 15102 27004 15108 27016
rect 15160 27044 15166 27056
rect 15197 27047 15255 27053
rect 15197 27044 15209 27047
rect 15160 27016 15209 27044
rect 15160 27004 15166 27016
rect 15197 27013 15209 27016
rect 15243 27013 15255 27047
rect 15197 27007 15255 27013
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11164 26948 11713 26976
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 12342 26976 12348 26988
rect 12303 26948 12348 26976
rect 11701 26939 11759 26945
rect 12342 26936 12348 26948
rect 12400 26936 12406 26988
rect 13357 26979 13415 26985
rect 13357 26945 13369 26979
rect 13403 26945 13415 26979
rect 14734 26976 14740 26988
rect 14695 26948 14740 26976
rect 13357 26939 13415 26945
rect 9490 26908 9496 26920
rect 3835 26880 9260 26908
rect 9451 26880 9496 26908
rect 3835 26877 3847 26880
rect 3789 26871 3847 26877
rect 9490 26868 9496 26880
rect 9548 26868 9554 26920
rect 10594 26908 10600 26920
rect 10555 26880 10600 26908
rect 10594 26868 10600 26880
rect 10652 26868 10658 26920
rect 10689 26911 10747 26917
rect 10689 26877 10701 26911
rect 10735 26908 10747 26911
rect 11514 26908 11520 26920
rect 10735 26880 11520 26908
rect 10735 26877 10747 26880
rect 10689 26871 10747 26877
rect 2746 26812 5396 26840
rect 2041 26775 2099 26781
rect 2041 26741 2053 26775
rect 2087 26772 2099 26775
rect 2866 26772 2872 26784
rect 2087 26744 2872 26772
rect 2087 26741 2099 26744
rect 2041 26735 2099 26741
rect 2866 26732 2872 26744
rect 2924 26732 2930 26784
rect 5368 26772 5396 26812
rect 5442 26800 5448 26852
rect 5500 26840 5506 26852
rect 7193 26843 7251 26849
rect 7193 26840 7205 26843
rect 5500 26812 7205 26840
rect 5500 26800 5506 26812
rect 7193 26809 7205 26812
rect 7239 26809 7251 26843
rect 7193 26803 7251 26809
rect 7558 26800 7564 26852
rect 7616 26840 7622 26852
rect 10704 26840 10732 26871
rect 11514 26868 11520 26880
rect 11572 26908 11578 26920
rect 11974 26908 11980 26920
rect 11572 26880 11980 26908
rect 11572 26868 11578 26880
rect 11974 26868 11980 26880
rect 12032 26868 12038 26920
rect 13372 26908 13400 26939
rect 14734 26936 14740 26948
rect 14792 26936 14798 26988
rect 13446 26908 13452 26920
rect 13372 26880 13452 26908
rect 13446 26868 13452 26880
rect 13504 26868 13510 26920
rect 13633 26911 13691 26917
rect 13633 26877 13645 26911
rect 13679 26908 13691 26911
rect 13998 26908 14004 26920
rect 13679 26880 14004 26908
rect 13679 26877 13691 26880
rect 13633 26871 13691 26877
rect 13998 26868 14004 26880
rect 14056 26908 14062 26920
rect 15010 26908 15016 26920
rect 14056 26880 15016 26908
rect 14056 26868 14062 26880
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 17037 26911 17095 26917
rect 17037 26877 17049 26911
rect 17083 26908 17095 26911
rect 17494 26908 17500 26920
rect 17083 26880 17500 26908
rect 17083 26877 17095 26880
rect 17037 26871 17095 26877
rect 17494 26868 17500 26880
rect 17552 26868 17558 26920
rect 7616 26812 10732 26840
rect 11885 26843 11943 26849
rect 7616 26800 7622 26812
rect 11885 26809 11897 26843
rect 11931 26840 11943 26843
rect 13354 26840 13360 26852
rect 11931 26812 13360 26840
rect 11931 26809 11943 26812
rect 11885 26803 11943 26809
rect 13354 26800 13360 26812
rect 13412 26800 13418 26852
rect 5626 26772 5632 26784
rect 5368 26744 5632 26772
rect 5626 26732 5632 26744
rect 5684 26732 5690 26784
rect 5902 26772 5908 26784
rect 5863 26744 5908 26772
rect 5902 26732 5908 26744
rect 5960 26732 5966 26784
rect 6733 26775 6791 26781
rect 6733 26741 6745 26775
rect 6779 26772 6791 26775
rect 6822 26772 6828 26784
rect 6779 26744 6828 26772
rect 6779 26741 6791 26744
rect 6733 26735 6791 26741
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 8389 26775 8447 26781
rect 8389 26741 8401 26775
rect 8435 26772 8447 26775
rect 8478 26772 8484 26784
rect 8435 26744 8484 26772
rect 8435 26741 8447 26744
rect 8389 26735 8447 26741
rect 8478 26732 8484 26744
rect 8536 26732 8542 26784
rect 12529 26775 12587 26781
rect 12529 26741 12541 26775
rect 12575 26772 12587 26775
rect 12710 26772 12716 26784
rect 12575 26744 12716 26772
rect 12575 26741 12587 26744
rect 12529 26735 12587 26741
rect 12710 26732 12716 26744
rect 12768 26732 12774 26784
rect 12986 26772 12992 26784
rect 12947 26744 12992 26772
rect 12986 26732 12992 26744
rect 13044 26732 13050 26784
rect 15746 26772 15752 26784
rect 15707 26744 15752 26772
rect 15746 26732 15752 26744
rect 15804 26732 15810 26784
rect 17586 26772 17592 26784
rect 17547 26744 17592 26772
rect 17586 26732 17592 26744
rect 17644 26732 17650 26784
rect 56965 26775 57023 26781
rect 56965 26741 56977 26775
rect 57011 26772 57023 26775
rect 57146 26772 57152 26784
rect 57011 26744 57152 26772
rect 57011 26741 57023 26744
rect 56965 26735 57023 26741
rect 57146 26732 57152 26744
rect 57204 26732 57210 26784
rect 57514 26772 57520 26784
rect 57427 26744 57520 26772
rect 57514 26732 57520 26744
rect 57572 26772 57578 26784
rect 57790 26772 57796 26784
rect 57572 26744 57796 26772
rect 57572 26732 57578 26744
rect 57790 26732 57796 26744
rect 57848 26732 57854 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 4062 26528 4068 26580
rect 4120 26568 4126 26580
rect 8662 26568 8668 26580
rect 4120 26540 8668 26568
rect 4120 26528 4126 26540
rect 1670 26500 1676 26512
rect 1631 26472 1676 26500
rect 1670 26460 1676 26472
rect 1728 26460 1734 26512
rect 2130 26392 2136 26444
rect 2188 26432 2194 26444
rect 2777 26435 2835 26441
rect 2777 26432 2789 26435
rect 2188 26404 2789 26432
rect 2188 26392 2194 26404
rect 2777 26401 2789 26404
rect 2823 26432 2835 26435
rect 3970 26432 3976 26444
rect 2823 26404 3976 26432
rect 2823 26401 2835 26404
rect 2777 26395 2835 26401
rect 3970 26392 3976 26404
rect 4028 26432 4034 26444
rect 4264 26441 4292 26540
rect 8662 26528 8668 26540
rect 8720 26528 8726 26580
rect 9306 26528 9312 26580
rect 9364 26568 9370 26580
rect 9950 26568 9956 26580
rect 9364 26540 9956 26568
rect 9364 26528 9370 26540
rect 9950 26528 9956 26540
rect 10008 26568 10014 26580
rect 10045 26571 10103 26577
rect 10045 26568 10057 26571
rect 10008 26540 10057 26568
rect 10008 26528 10014 26540
rect 10045 26537 10057 26540
rect 10091 26537 10103 26571
rect 10045 26531 10103 26537
rect 10594 26528 10600 26580
rect 10652 26568 10658 26580
rect 11333 26571 11391 26577
rect 11333 26568 11345 26571
rect 10652 26540 11345 26568
rect 10652 26528 10658 26540
rect 11333 26537 11345 26540
rect 11379 26568 11391 26571
rect 12621 26571 12679 26577
rect 11379 26540 12434 26568
rect 11379 26537 11391 26540
rect 11333 26531 11391 26537
rect 4709 26503 4767 26509
rect 4709 26469 4721 26503
rect 4755 26469 4767 26503
rect 4709 26463 4767 26469
rect 5905 26503 5963 26509
rect 5905 26469 5917 26503
rect 5951 26500 5963 26503
rect 8202 26500 8208 26512
rect 5951 26472 8208 26500
rect 5951 26469 5963 26472
rect 5905 26463 5963 26469
rect 4065 26435 4123 26441
rect 4065 26432 4077 26435
rect 4028 26404 4077 26432
rect 4028 26392 4034 26404
rect 4065 26401 4077 26404
rect 4111 26401 4123 26435
rect 4065 26395 4123 26401
rect 4249 26435 4307 26441
rect 4249 26401 4261 26435
rect 4295 26401 4307 26435
rect 4249 26395 4307 26401
rect 1857 26367 1915 26373
rect 1857 26333 1869 26367
rect 1903 26364 1915 26367
rect 2866 26364 2872 26376
rect 1903 26336 2872 26364
rect 1903 26333 1915 26336
rect 1857 26327 1915 26333
rect 2866 26324 2872 26336
rect 2924 26324 2930 26376
rect 2961 26367 3019 26373
rect 2961 26333 2973 26367
rect 3007 26364 3019 26367
rect 4614 26364 4620 26376
rect 3007 26336 4620 26364
rect 3007 26333 3019 26336
rect 2961 26327 3019 26333
rect 4614 26324 4620 26336
rect 4672 26324 4678 26376
rect 4724 26364 4752 26463
rect 8202 26460 8208 26472
rect 8260 26460 8266 26512
rect 8294 26460 8300 26512
rect 8352 26500 8358 26512
rect 8573 26503 8631 26509
rect 8573 26500 8585 26503
rect 8352 26472 8585 26500
rect 8352 26460 8358 26472
rect 8573 26469 8585 26472
rect 8619 26500 8631 26503
rect 9490 26500 9496 26512
rect 8619 26472 9496 26500
rect 8619 26469 8631 26472
rect 8573 26463 8631 26469
rect 9490 26460 9496 26472
rect 9548 26460 9554 26512
rect 12069 26503 12127 26509
rect 12069 26469 12081 26503
rect 12115 26500 12127 26503
rect 12158 26500 12164 26512
rect 12115 26472 12164 26500
rect 12115 26469 12127 26472
rect 12069 26463 12127 26469
rect 12158 26460 12164 26472
rect 12216 26460 12222 26512
rect 12406 26500 12434 26540
rect 12621 26537 12633 26571
rect 12667 26568 12679 26571
rect 13262 26568 13268 26580
rect 12667 26540 13268 26568
rect 12667 26537 12679 26540
rect 12621 26531 12679 26537
rect 13262 26528 13268 26540
rect 13320 26528 13326 26580
rect 14734 26568 14740 26580
rect 14695 26540 14740 26568
rect 14734 26528 14740 26540
rect 14792 26528 14798 26580
rect 15010 26528 15016 26580
rect 15068 26568 15074 26580
rect 15068 26540 17816 26568
rect 15068 26528 15074 26540
rect 13814 26500 13820 26512
rect 12406 26472 13820 26500
rect 13814 26460 13820 26472
rect 13872 26460 13878 26512
rect 15102 26460 15108 26512
rect 15160 26500 15166 26512
rect 15160 26472 15332 26500
rect 15160 26460 15166 26472
rect 6178 26392 6184 26444
rect 6236 26432 6242 26444
rect 6457 26435 6515 26441
rect 6457 26432 6469 26435
rect 6236 26404 6469 26432
rect 6236 26392 6242 26404
rect 6457 26401 6469 26404
rect 6503 26401 6515 26435
rect 6638 26432 6644 26444
rect 6599 26404 6644 26432
rect 6457 26395 6515 26401
rect 5721 26367 5779 26373
rect 5721 26364 5733 26367
rect 4724 26336 5733 26364
rect 5721 26333 5733 26336
rect 5767 26333 5779 26367
rect 6472 26364 6500 26395
rect 6638 26392 6644 26404
rect 6696 26432 6702 26444
rect 7561 26435 7619 26441
rect 7561 26432 7573 26435
rect 6696 26404 7573 26432
rect 6696 26392 6702 26404
rect 7561 26401 7573 26404
rect 7607 26401 7619 26435
rect 10410 26432 10416 26444
rect 7561 26395 7619 26401
rect 8496 26404 10416 26432
rect 6546 26364 6552 26376
rect 6472 26336 6552 26364
rect 5721 26327 5779 26333
rect 6546 26324 6552 26336
rect 6604 26324 6610 26376
rect 2038 26256 2044 26308
rect 2096 26296 2102 26308
rect 2590 26296 2596 26308
rect 2096 26268 2596 26296
rect 2096 26256 2102 26268
rect 2590 26256 2596 26268
rect 2648 26296 2654 26308
rect 3053 26299 3111 26305
rect 3053 26296 3065 26299
rect 2648 26268 3065 26296
rect 2648 26256 2654 26268
rect 3053 26265 3065 26268
rect 3099 26265 3111 26299
rect 3053 26259 3111 26265
rect 4341 26299 4399 26305
rect 4341 26265 4353 26299
rect 4387 26296 4399 26299
rect 5261 26299 5319 26305
rect 5261 26296 5273 26299
rect 4387 26268 5273 26296
rect 4387 26265 4399 26268
rect 4341 26259 4399 26265
rect 5261 26265 5273 26268
rect 5307 26296 5319 26299
rect 5442 26296 5448 26308
rect 5307 26268 5448 26296
rect 5307 26265 5319 26268
rect 5261 26259 5319 26265
rect 5442 26256 5448 26268
rect 5500 26256 5506 26308
rect 5626 26256 5632 26308
rect 5684 26296 5690 26308
rect 8496 26296 8524 26404
rect 10410 26392 10416 26404
rect 10468 26432 10474 26444
rect 15304 26441 15332 26472
rect 17586 26460 17592 26512
rect 17644 26460 17650 26512
rect 13633 26435 13691 26441
rect 13633 26432 13645 26435
rect 10468 26404 13645 26432
rect 10468 26392 10474 26404
rect 13633 26401 13645 26404
rect 13679 26432 13691 26435
rect 15197 26435 15255 26441
rect 15197 26432 15209 26435
rect 13679 26404 15209 26432
rect 13679 26401 13691 26404
rect 13633 26395 13691 26401
rect 15197 26401 15209 26404
rect 15243 26401 15255 26435
rect 15197 26395 15255 26401
rect 15289 26435 15347 26441
rect 15289 26401 15301 26435
rect 15335 26432 15347 26435
rect 16485 26435 16543 26441
rect 16485 26432 16497 26435
rect 15335 26404 16497 26432
rect 15335 26401 15347 26404
rect 15289 26395 15347 26401
rect 16485 26401 16497 26404
rect 16531 26401 16543 26435
rect 17604 26432 17632 26460
rect 17788 26441 17816 26540
rect 57974 26500 57980 26512
rect 57624 26472 57980 26500
rect 57330 26441 57336 26444
rect 16485 26395 16543 26401
rect 16684 26404 17632 26432
rect 17773 26435 17831 26441
rect 11885 26367 11943 26373
rect 11885 26333 11897 26367
rect 11931 26364 11943 26367
rect 12986 26364 12992 26376
rect 11931 26336 12992 26364
rect 11931 26333 11943 26336
rect 11885 26327 11943 26333
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 13173 26367 13231 26373
rect 13173 26333 13185 26367
rect 13219 26364 13231 26367
rect 13446 26364 13452 26376
rect 13219 26336 13452 26364
rect 13219 26333 13231 26336
rect 13173 26327 13231 26333
rect 13446 26324 13452 26336
rect 13504 26364 13510 26376
rect 15105 26367 15163 26373
rect 15105 26364 15117 26367
rect 13504 26336 15117 26364
rect 13504 26324 13510 26336
rect 15105 26333 15117 26336
rect 15151 26364 15163 26367
rect 15470 26364 15476 26376
rect 15151 26336 15476 26364
rect 15151 26333 15163 26336
rect 15105 26327 15163 26333
rect 15470 26324 15476 26336
rect 15528 26364 15534 26376
rect 15746 26364 15752 26376
rect 15528 26336 15752 26364
rect 15528 26324 15534 26336
rect 15746 26324 15752 26336
rect 15804 26324 15810 26376
rect 16500 26364 16528 26395
rect 16684 26364 16712 26404
rect 17773 26401 17785 26435
rect 17819 26432 17831 26435
rect 57308 26435 57336 26441
rect 17819 26404 18460 26432
rect 17819 26401 17831 26404
rect 17773 26395 17831 26401
rect 16500 26336 16712 26364
rect 16758 26324 16764 26376
rect 16816 26364 16822 26376
rect 17589 26367 17647 26373
rect 17589 26364 17601 26367
rect 16816 26336 17601 26364
rect 16816 26324 16822 26336
rect 17589 26333 17601 26336
rect 17635 26333 17647 26367
rect 17589 26327 17647 26333
rect 9122 26296 9128 26308
rect 5684 26268 8524 26296
rect 9083 26268 9128 26296
rect 5684 26256 5690 26268
rect 9122 26256 9128 26268
rect 9180 26256 9186 26308
rect 18432 26305 18460 26404
rect 57308 26401 57320 26435
rect 57308 26395 57336 26401
rect 57330 26392 57336 26395
rect 57388 26392 57394 26444
rect 57425 26435 57483 26441
rect 57425 26401 57437 26435
rect 57471 26432 57483 26435
rect 57624 26432 57652 26472
rect 57974 26460 57980 26472
rect 58032 26460 58038 26512
rect 57471 26404 57652 26432
rect 57701 26435 57759 26441
rect 57471 26401 57483 26404
rect 57425 26395 57483 26401
rect 57701 26401 57713 26435
rect 57747 26432 57759 26435
rect 57790 26432 57796 26444
rect 57747 26404 57796 26432
rect 57747 26401 57759 26404
rect 57701 26395 57759 26401
rect 57790 26392 57796 26404
rect 57848 26392 57854 26444
rect 58345 26435 58403 26441
rect 58345 26401 58357 26435
rect 58391 26432 58403 26435
rect 58434 26432 58440 26444
rect 58391 26404 58440 26432
rect 58391 26401 58403 26404
rect 58345 26395 58403 26401
rect 58434 26392 58440 26404
rect 58492 26392 58498 26444
rect 44545 26367 44603 26373
rect 44545 26333 44557 26367
rect 44591 26364 44603 26367
rect 56505 26367 56563 26373
rect 56505 26364 56517 26367
rect 44591 26336 56517 26364
rect 44591 26333 44603 26336
rect 44545 26327 44603 26333
rect 56505 26333 56517 26336
rect 56551 26333 56563 26367
rect 56505 26327 56563 26333
rect 57146 26324 57152 26376
rect 57204 26364 57210 26376
rect 58161 26367 58219 26373
rect 57204 26336 57249 26364
rect 57204 26324 57210 26336
rect 58161 26333 58173 26367
rect 58207 26364 58219 26367
rect 58207 26336 58480 26364
rect 58207 26333 58219 26336
rect 58161 26327 58219 26333
rect 58452 26308 58480 26336
rect 16301 26299 16359 26305
rect 11164 26268 11376 26296
rect 3421 26231 3479 26237
rect 3421 26197 3433 26231
rect 3467 26228 3479 26231
rect 3694 26228 3700 26240
rect 3467 26200 3700 26228
rect 3467 26197 3479 26200
rect 3421 26191 3479 26197
rect 3694 26188 3700 26200
rect 3752 26188 3758 26240
rect 6730 26228 6736 26240
rect 6691 26200 6736 26228
rect 6730 26188 6736 26200
rect 6788 26188 6794 26240
rect 7101 26231 7159 26237
rect 7101 26197 7113 26231
rect 7147 26228 7159 26231
rect 7190 26228 7196 26240
rect 7147 26200 7196 26228
rect 7147 26197 7159 26200
rect 7101 26191 7159 26197
rect 7190 26188 7196 26200
rect 7248 26188 7254 26240
rect 9140 26228 9168 26256
rect 11164 26228 11192 26268
rect 9140 26200 11192 26228
rect 11348 26228 11376 26268
rect 16301 26265 16313 26299
rect 16347 26296 16359 26299
rect 18417 26299 18475 26305
rect 16347 26268 17540 26296
rect 16347 26265 16359 26268
rect 16301 26259 16359 26265
rect 17512 26240 17540 26268
rect 18417 26265 18429 26299
rect 18463 26296 18475 26299
rect 19426 26296 19432 26308
rect 18463 26268 19432 26296
rect 18463 26265 18475 26268
rect 18417 26259 18475 26265
rect 19426 26256 19432 26268
rect 19484 26256 19490 26308
rect 58434 26256 58440 26308
rect 58492 26256 58498 26308
rect 14090 26228 14096 26240
rect 11348 26200 14096 26228
rect 14090 26188 14096 26200
rect 14148 26188 14154 26240
rect 15930 26228 15936 26240
rect 15891 26200 15936 26228
rect 15930 26188 15936 26200
rect 15988 26188 15994 26240
rect 16390 26228 16396 26240
rect 16351 26200 16396 26228
rect 16390 26188 16396 26200
rect 16448 26188 16454 26240
rect 17034 26188 17040 26240
rect 17092 26228 17098 26240
rect 17129 26231 17187 26237
rect 17129 26228 17141 26231
rect 17092 26200 17141 26228
rect 17092 26188 17098 26200
rect 17129 26197 17141 26200
rect 17175 26197 17187 26231
rect 17494 26228 17500 26240
rect 17455 26200 17500 26228
rect 17129 26191 17187 26197
rect 17494 26188 17500 26200
rect 17552 26228 17558 26240
rect 44358 26228 44364 26240
rect 17552 26200 17577 26228
rect 44319 26200 44364 26228
rect 17552 26188 17558 26200
rect 44358 26188 44364 26200
rect 44416 26188 44422 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 2774 25984 2780 26036
rect 2832 26024 2838 26036
rect 2832 25996 10272 26024
rect 2832 25984 2838 25996
rect 1854 25916 1860 25968
rect 1912 25956 1918 25968
rect 8113 25959 8171 25965
rect 8113 25956 8125 25959
rect 1912 25928 8125 25956
rect 1912 25916 1918 25928
rect 8113 25925 8125 25928
rect 8159 25956 8171 25959
rect 9122 25956 9128 25968
rect 8159 25928 9128 25956
rect 8159 25925 8171 25928
rect 8113 25919 8171 25925
rect 9122 25916 9128 25928
rect 9180 25916 9186 25968
rect 1762 25848 1768 25900
rect 1820 25888 1826 25900
rect 2409 25891 2467 25897
rect 2409 25888 2421 25891
rect 1820 25860 2421 25888
rect 1820 25848 1826 25860
rect 2409 25857 2421 25860
rect 2455 25857 2467 25891
rect 3694 25888 3700 25900
rect 3655 25860 3700 25888
rect 2409 25851 2467 25857
rect 3694 25848 3700 25860
rect 3752 25848 3758 25900
rect 3970 25848 3976 25900
rect 4028 25888 4034 25900
rect 4801 25891 4859 25897
rect 4801 25888 4813 25891
rect 4028 25860 4813 25888
rect 4028 25848 4034 25860
rect 4801 25857 4813 25860
rect 4847 25857 4859 25891
rect 7190 25888 7196 25900
rect 7151 25860 7196 25888
rect 4801 25851 4859 25857
rect 7190 25848 7196 25860
rect 7248 25848 7254 25900
rect 8205 25891 8263 25897
rect 8205 25888 8217 25891
rect 7300 25860 8217 25888
rect 2130 25820 2136 25832
rect 2091 25792 2136 25820
rect 2130 25780 2136 25792
rect 2188 25780 2194 25832
rect 2314 25780 2320 25832
rect 2372 25820 2378 25832
rect 2682 25820 2688 25832
rect 2372 25792 2688 25820
rect 2372 25780 2378 25792
rect 2682 25780 2688 25792
rect 2740 25780 2746 25832
rect 3326 25780 3332 25832
rect 3384 25820 3390 25832
rect 7300 25820 7328 25860
rect 8205 25857 8217 25860
rect 8251 25888 8263 25891
rect 8386 25888 8392 25900
rect 8251 25860 8392 25888
rect 8251 25857 8263 25860
rect 8205 25851 8263 25857
rect 8386 25848 8392 25860
rect 8444 25848 8450 25900
rect 9677 25891 9735 25897
rect 9677 25857 9689 25891
rect 9723 25888 9735 25891
rect 9723 25860 10180 25888
rect 9723 25857 9735 25860
rect 9677 25851 9735 25857
rect 8021 25823 8079 25829
rect 8021 25820 8033 25823
rect 3384 25792 7328 25820
rect 7392 25792 8033 25820
rect 3384 25780 3390 25792
rect 6546 25712 6552 25764
rect 6604 25752 6610 25764
rect 6733 25755 6791 25761
rect 6733 25752 6745 25755
rect 6604 25724 6745 25752
rect 6604 25712 6610 25724
rect 6733 25721 6745 25724
rect 6779 25752 6791 25755
rect 7392 25752 7420 25792
rect 8021 25789 8033 25792
rect 8067 25820 8079 25823
rect 8294 25820 8300 25832
rect 8067 25792 8300 25820
rect 8067 25789 8079 25792
rect 8021 25783 8079 25789
rect 8294 25780 8300 25792
rect 8352 25780 8358 25832
rect 9306 25752 9312 25764
rect 6779 25724 7420 25752
rect 8404 25724 9312 25752
rect 6779 25721 6791 25724
rect 6733 25715 6791 25721
rect 2406 25644 2412 25696
rect 2464 25684 2470 25696
rect 2777 25687 2835 25693
rect 2777 25684 2789 25687
rect 2464 25656 2789 25684
rect 2464 25644 2470 25656
rect 2777 25653 2789 25656
rect 2823 25653 2835 25687
rect 3878 25684 3884 25696
rect 3839 25656 3884 25684
rect 2777 25647 2835 25653
rect 3878 25644 3884 25656
rect 3936 25644 3942 25696
rect 7377 25687 7435 25693
rect 7377 25653 7389 25687
rect 7423 25684 7435 25687
rect 8404 25684 8432 25724
rect 9306 25712 9312 25724
rect 9364 25712 9370 25764
rect 10152 25761 10180 25860
rect 10244 25820 10272 25996
rect 15378 25984 15384 26036
rect 15436 26024 15442 26036
rect 16390 26024 16396 26036
rect 15436 25996 16396 26024
rect 15436 25984 15442 25996
rect 16390 25984 16396 25996
rect 16448 25984 16454 26036
rect 56042 25984 56048 26036
rect 56100 26024 56106 26036
rect 57333 26027 57391 26033
rect 57333 26024 57345 26027
rect 56100 25996 57345 26024
rect 56100 25984 56106 25996
rect 57333 25993 57345 25996
rect 57379 25993 57391 26027
rect 57333 25987 57391 25993
rect 58161 26027 58219 26033
rect 58161 25993 58173 26027
rect 58207 26024 58219 26027
rect 58802 26024 58808 26036
rect 58207 25996 58808 26024
rect 58207 25993 58219 25996
rect 58161 25987 58219 25993
rect 58802 25984 58808 25996
rect 58860 25984 58866 26036
rect 56321 25959 56379 25965
rect 56321 25925 56333 25959
rect 56367 25956 56379 25959
rect 56367 25928 58388 25956
rect 56367 25925 56379 25928
rect 56321 25919 56379 25925
rect 58360 25900 58388 25928
rect 10318 25848 10324 25900
rect 10376 25888 10382 25900
rect 10505 25891 10563 25897
rect 10505 25888 10517 25891
rect 10376 25860 10517 25888
rect 10376 25848 10382 25860
rect 10505 25857 10517 25860
rect 10551 25857 10563 25891
rect 10505 25851 10563 25857
rect 10594 25848 10600 25900
rect 10652 25888 10658 25900
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 10652 25860 11713 25888
rect 10652 25848 10658 25860
rect 11701 25857 11713 25860
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 13357 25891 13415 25897
rect 13357 25857 13369 25891
rect 13403 25888 13415 25891
rect 14185 25891 14243 25897
rect 13403 25860 13860 25888
rect 13403 25857 13415 25860
rect 13357 25851 13415 25857
rect 10686 25820 10692 25832
rect 10244 25792 10692 25820
rect 10686 25780 10692 25792
rect 10744 25820 10750 25832
rect 10744 25792 10837 25820
rect 10744 25780 10750 25792
rect 13832 25761 13860 25860
rect 14185 25857 14197 25891
rect 14231 25888 14243 25891
rect 15470 25888 15476 25900
rect 14231 25860 15476 25888
rect 14231 25857 14243 25860
rect 14185 25851 14243 25857
rect 15470 25848 15476 25860
rect 15528 25848 15534 25900
rect 15930 25848 15936 25900
rect 15988 25888 15994 25900
rect 16025 25891 16083 25897
rect 16025 25888 16037 25891
rect 15988 25860 16037 25888
rect 15988 25848 15994 25860
rect 16025 25857 16037 25860
rect 16071 25857 16083 25891
rect 17034 25888 17040 25900
rect 16995 25860 17040 25888
rect 16025 25851 16083 25857
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 56873 25891 56931 25897
rect 56873 25857 56885 25891
rect 56919 25888 56931 25891
rect 57514 25888 57520 25900
rect 56919 25860 57520 25888
rect 56919 25857 56931 25860
rect 56873 25851 56931 25857
rect 57514 25848 57520 25860
rect 57572 25848 57578 25900
rect 58342 25888 58348 25900
rect 58303 25860 58348 25888
rect 58342 25848 58348 25860
rect 58400 25848 58406 25900
rect 14274 25820 14280 25832
rect 14235 25792 14280 25820
rect 14274 25780 14280 25792
rect 14332 25780 14338 25832
rect 14458 25820 14464 25832
rect 14419 25792 14464 25820
rect 14458 25780 14464 25792
rect 14516 25780 14522 25832
rect 10137 25755 10195 25761
rect 10137 25721 10149 25755
rect 10183 25721 10195 25755
rect 10137 25715 10195 25721
rect 13817 25755 13875 25761
rect 13817 25721 13829 25755
rect 13863 25721 13875 25755
rect 13817 25715 13875 25721
rect 13998 25712 14004 25764
rect 14056 25752 14062 25764
rect 15841 25755 15899 25761
rect 15841 25752 15853 25755
rect 14056 25724 15853 25752
rect 14056 25712 14062 25724
rect 15841 25721 15853 25724
rect 15887 25721 15899 25755
rect 15841 25715 15899 25721
rect 7423 25656 8432 25684
rect 8573 25687 8631 25693
rect 7423 25653 7435 25656
rect 7377 25647 7435 25653
rect 8573 25653 8585 25687
rect 8619 25684 8631 25687
rect 9122 25684 9128 25696
rect 8619 25656 9128 25684
rect 8619 25653 8631 25656
rect 8573 25647 8631 25653
rect 9122 25644 9128 25656
rect 9180 25644 9186 25696
rect 9398 25644 9404 25696
rect 9456 25684 9462 25696
rect 9493 25687 9551 25693
rect 9493 25684 9505 25687
rect 9456 25656 9505 25684
rect 9456 25644 9462 25656
rect 9493 25653 9505 25656
rect 9539 25653 9551 25687
rect 13170 25684 13176 25696
rect 13131 25656 13176 25684
rect 9493 25647 9551 25653
rect 13170 25644 13176 25656
rect 13228 25644 13234 25696
rect 15378 25684 15384 25696
rect 15339 25656 15384 25684
rect 15378 25644 15384 25656
rect 15436 25644 15442 25696
rect 15930 25644 15936 25696
rect 15988 25684 15994 25696
rect 16853 25687 16911 25693
rect 16853 25684 16865 25687
rect 15988 25656 16865 25684
rect 15988 25644 15994 25656
rect 16853 25653 16865 25656
rect 16899 25653 16911 25687
rect 16853 25647 16911 25653
rect 17494 25644 17500 25696
rect 17552 25684 17558 25696
rect 17589 25687 17647 25693
rect 17589 25684 17601 25687
rect 17552 25656 17601 25684
rect 17552 25644 17558 25656
rect 17589 25653 17601 25656
rect 17635 25684 17647 25687
rect 19242 25684 19248 25696
rect 17635 25656 19248 25684
rect 17635 25653 17647 25656
rect 17589 25647 17647 25653
rect 19242 25644 19248 25656
rect 19300 25644 19306 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1670 25480 1676 25492
rect 1631 25452 1676 25480
rect 1670 25440 1676 25452
rect 1728 25440 1734 25492
rect 3142 25480 3148 25492
rect 3055 25452 3148 25480
rect 3142 25440 3148 25452
rect 3200 25480 3206 25492
rect 5350 25480 5356 25492
rect 3200 25452 5356 25480
rect 3200 25440 3206 25452
rect 5350 25440 5356 25452
rect 5408 25440 5414 25492
rect 6730 25440 6736 25492
rect 6788 25480 6794 25492
rect 7377 25483 7435 25489
rect 7377 25480 7389 25483
rect 6788 25452 7389 25480
rect 6788 25440 6794 25452
rect 7377 25449 7389 25452
rect 7423 25449 7435 25483
rect 7377 25443 7435 25449
rect 8386 25440 8392 25492
rect 8444 25480 8450 25492
rect 8481 25483 8539 25489
rect 8481 25480 8493 25483
rect 8444 25452 8493 25480
rect 8444 25440 8450 25452
rect 8481 25449 8493 25452
rect 8527 25449 8539 25483
rect 8481 25443 8539 25449
rect 10686 25440 10692 25492
rect 10744 25480 10750 25492
rect 11701 25483 11759 25489
rect 11701 25480 11713 25483
rect 10744 25452 11713 25480
rect 10744 25440 10750 25452
rect 11701 25449 11713 25452
rect 11747 25480 11759 25483
rect 14458 25480 14464 25492
rect 11747 25452 14464 25480
rect 11747 25449 11759 25452
rect 11701 25443 11759 25449
rect 14458 25440 14464 25452
rect 14516 25480 14522 25492
rect 14516 25452 16574 25480
rect 14516 25440 14522 25452
rect 2593 25415 2651 25421
rect 2593 25381 2605 25415
rect 2639 25412 2651 25415
rect 5534 25412 5540 25424
rect 2639 25384 5540 25412
rect 2639 25381 2651 25384
rect 2593 25375 2651 25381
rect 5534 25372 5540 25384
rect 5592 25372 5598 25424
rect 3234 25304 3240 25356
rect 3292 25344 3298 25356
rect 6748 25344 6776 25440
rect 9309 25415 9367 25421
rect 9309 25381 9321 25415
rect 9355 25412 9367 25415
rect 15286 25412 15292 25424
rect 9355 25384 15292 25412
rect 9355 25381 9367 25384
rect 9309 25375 9367 25381
rect 15286 25372 15292 25384
rect 15344 25372 15350 25424
rect 3292 25316 6776 25344
rect 3292 25304 3298 25316
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25276 1915 25279
rect 2222 25276 2228 25288
rect 1903 25248 2228 25276
rect 1903 25245 1915 25248
rect 1857 25239 1915 25245
rect 2222 25236 2228 25248
rect 2280 25236 2286 25288
rect 2406 25276 2412 25288
rect 2367 25248 2412 25276
rect 2406 25236 2412 25248
rect 2464 25236 2470 25288
rect 9122 25276 9128 25288
rect 9083 25248 9128 25276
rect 9122 25236 9128 25248
rect 9180 25236 9186 25288
rect 16546 25208 16574 25452
rect 58894 25412 58900 25424
rect 57624 25384 58900 25412
rect 57330 25353 57336 25356
rect 57308 25347 57336 25353
rect 57308 25313 57320 25347
rect 57308 25307 57336 25313
rect 57330 25304 57336 25307
rect 57388 25304 57394 25356
rect 57425 25347 57483 25353
rect 57425 25313 57437 25347
rect 57471 25344 57483 25347
rect 57624 25344 57652 25384
rect 58894 25372 58900 25384
rect 58952 25372 58958 25424
rect 57471 25316 57652 25344
rect 57701 25347 57759 25353
rect 57471 25313 57483 25316
rect 57425 25307 57483 25313
rect 57701 25313 57713 25347
rect 57747 25344 57759 25347
rect 57790 25344 57796 25356
rect 57747 25316 57796 25344
rect 57747 25313 57759 25316
rect 57701 25307 57759 25313
rect 57790 25304 57796 25316
rect 57848 25304 57854 25356
rect 58250 25304 58256 25356
rect 58308 25344 58314 25356
rect 58345 25347 58403 25353
rect 58345 25344 58357 25347
rect 58308 25316 58357 25344
rect 58308 25304 58314 25316
rect 58345 25313 58357 25316
rect 58391 25313 58403 25347
rect 58345 25307 58403 25313
rect 57146 25236 57152 25288
rect 57204 25276 57210 25288
rect 58158 25276 58164 25288
rect 57204 25248 57249 25276
rect 58119 25248 58164 25276
rect 57204 25236 57210 25248
rect 58158 25236 58164 25248
rect 58216 25236 58222 25288
rect 17402 25208 17408 25220
rect 16546 25180 17408 25208
rect 17402 25168 17408 25180
rect 17460 25168 17466 25220
rect 1762 25100 1768 25152
rect 1820 25140 1826 25152
rect 3142 25140 3148 25152
rect 1820 25112 3148 25140
rect 1820 25100 1826 25112
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 10318 25100 10324 25152
rect 10376 25140 10382 25152
rect 11149 25143 11207 25149
rect 11149 25140 11161 25143
rect 10376 25112 11161 25140
rect 10376 25100 10382 25112
rect 11149 25109 11161 25112
rect 11195 25109 11207 25143
rect 11149 25103 11207 25109
rect 14274 25100 14280 25152
rect 14332 25140 14338 25152
rect 15013 25143 15071 25149
rect 15013 25140 15025 25143
rect 14332 25112 15025 25140
rect 14332 25100 14338 25112
rect 15013 25109 15025 25112
rect 15059 25109 15071 25143
rect 15013 25103 15071 25109
rect 15470 25100 15476 25152
rect 15528 25140 15534 25152
rect 15565 25143 15623 25149
rect 15565 25140 15577 25143
rect 15528 25112 15577 25140
rect 15528 25100 15534 25112
rect 15565 25109 15577 25112
rect 15611 25109 15623 25143
rect 16758 25140 16764 25152
rect 16719 25112 16764 25140
rect 15565 25103 15623 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 56505 25143 56563 25149
rect 56505 25109 56517 25143
rect 56551 25140 56563 25143
rect 57974 25140 57980 25152
rect 56551 25112 57980 25140
rect 56551 25109 56563 25112
rect 56505 25103 56563 25109
rect 57974 25100 57980 25112
rect 58032 25100 58038 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 2406 24800 2412 24812
rect 1903 24772 2412 24800
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 2406 24760 2412 24772
rect 2464 24760 2470 24812
rect 58342 24800 58348 24812
rect 58303 24772 58348 24800
rect 58342 24760 58348 24772
rect 58400 24760 58406 24812
rect 2130 24692 2136 24744
rect 2188 24732 2194 24744
rect 2590 24732 2596 24744
rect 2188 24704 2596 24732
rect 2188 24692 2194 24704
rect 2590 24692 2596 24704
rect 2648 24732 2654 24744
rect 2869 24735 2927 24741
rect 2869 24732 2881 24735
rect 2648 24704 2881 24732
rect 2648 24692 2654 24704
rect 2869 24701 2881 24704
rect 2915 24701 2927 24735
rect 2869 24695 2927 24701
rect 1670 24664 1676 24676
rect 1631 24636 1676 24664
rect 1670 24624 1676 24636
rect 1728 24624 1734 24676
rect 56686 24624 56692 24676
rect 56744 24664 56750 24676
rect 57425 24667 57483 24673
rect 57425 24664 57437 24667
rect 56744 24636 57437 24664
rect 56744 24624 56750 24636
rect 57425 24633 57437 24636
rect 57471 24664 57483 24667
rect 57790 24664 57796 24676
rect 57471 24636 57796 24664
rect 57471 24633 57483 24636
rect 57425 24627 57483 24633
rect 57790 24624 57796 24636
rect 57848 24624 57854 24676
rect 58161 24667 58219 24673
rect 58161 24633 58173 24667
rect 58207 24664 58219 24667
rect 58618 24664 58624 24676
rect 58207 24636 58624 24664
rect 58207 24633 58219 24636
rect 58161 24627 58219 24633
rect 58618 24624 58624 24636
rect 58676 24624 58682 24676
rect 2222 24556 2228 24608
rect 2280 24596 2286 24608
rect 2317 24599 2375 24605
rect 2317 24596 2329 24599
rect 2280 24568 2329 24596
rect 2280 24556 2286 24568
rect 2317 24565 2329 24568
rect 2363 24565 2375 24599
rect 3510 24596 3516 24608
rect 3423 24568 3516 24596
rect 2317 24559 2375 24565
rect 3510 24556 3516 24568
rect 3568 24596 3574 24608
rect 14274 24596 14280 24608
rect 3568 24568 14280 24596
rect 3568 24556 3574 24568
rect 14274 24556 14280 24568
rect 14332 24596 14338 24608
rect 14642 24596 14648 24608
rect 14332 24568 14648 24596
rect 14332 24556 14338 24568
rect 14642 24556 14648 24568
rect 14700 24556 14706 24608
rect 56965 24599 57023 24605
rect 56965 24565 56977 24599
rect 57011 24596 57023 24599
rect 57146 24596 57152 24608
rect 57011 24568 57152 24596
rect 57011 24565 57023 24568
rect 56965 24559 57023 24565
rect 57146 24556 57152 24568
rect 57204 24596 57210 24608
rect 57330 24596 57336 24608
rect 57204 24568 57336 24596
rect 57204 24556 57210 24568
rect 57330 24556 57336 24568
rect 57388 24556 57394 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 2590 24352 2596 24404
rect 2648 24392 2654 24404
rect 2869 24395 2927 24401
rect 2869 24392 2881 24395
rect 2648 24364 2881 24392
rect 2648 24352 2654 24364
rect 2869 24361 2881 24364
rect 2915 24361 2927 24395
rect 2869 24355 2927 24361
rect 19426 24352 19432 24404
rect 19484 24392 19490 24404
rect 19521 24395 19579 24401
rect 19521 24392 19533 24395
rect 19484 24364 19533 24392
rect 19484 24352 19490 24364
rect 19521 24361 19533 24364
rect 19567 24361 19579 24395
rect 19521 24355 19579 24361
rect 57701 24395 57759 24401
rect 57701 24361 57713 24395
rect 57747 24392 57759 24395
rect 58342 24392 58348 24404
rect 57747 24364 58348 24392
rect 57747 24361 57759 24364
rect 57701 24355 57759 24361
rect 58342 24352 58348 24364
rect 58400 24352 58406 24404
rect 57238 24284 57244 24336
rect 57296 24324 57302 24336
rect 58161 24327 58219 24333
rect 58161 24324 58173 24327
rect 57296 24296 58173 24324
rect 57296 24284 57302 24296
rect 58161 24293 58173 24296
rect 58207 24293 58219 24327
rect 58161 24287 58219 24293
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24188 1915 24191
rect 3510 24188 3516 24200
rect 1903 24160 3516 24188
rect 1903 24157 1915 24160
rect 1857 24151 1915 24157
rect 3510 24148 3516 24160
rect 3568 24148 3574 24200
rect 57149 24191 57207 24197
rect 57149 24157 57161 24191
rect 57195 24188 57207 24191
rect 58342 24188 58348 24200
rect 57195 24160 58348 24188
rect 57195 24157 57207 24160
rect 57149 24151 57207 24157
rect 58342 24148 58348 24160
rect 58400 24148 58406 24200
rect 6362 24080 6368 24132
rect 6420 24120 6426 24132
rect 18598 24120 18604 24132
rect 6420 24092 18604 24120
rect 6420 24080 6426 24092
rect 18598 24080 18604 24092
rect 18656 24080 18662 24132
rect 19797 24123 19855 24129
rect 19797 24089 19809 24123
rect 19843 24089 19855 24123
rect 19797 24083 19855 24089
rect 1670 24052 1676 24064
rect 1631 24024 1676 24052
rect 1670 24012 1676 24024
rect 1728 24012 1734 24064
rect 2406 24052 2412 24064
rect 2367 24024 2412 24052
rect 2406 24012 2412 24024
rect 2464 24012 2470 24064
rect 19812 24052 19840 24083
rect 20438 24052 20444 24064
rect 19812 24024 20444 24052
rect 20438 24012 20444 24024
rect 20496 24012 20502 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 2406 23808 2412 23860
rect 2464 23848 2470 23860
rect 18414 23848 18420 23860
rect 2464 23820 18420 23848
rect 2464 23808 2470 23820
rect 18414 23808 18420 23820
rect 18472 23808 18478 23860
rect 58345 23851 58403 23857
rect 58345 23817 58357 23851
rect 58391 23848 58403 23851
rect 58894 23848 58900 23860
rect 58391 23820 58900 23848
rect 58391 23817 58403 23820
rect 58345 23811 58403 23817
rect 58894 23808 58900 23820
rect 58952 23808 58958 23860
rect 3237 23783 3295 23789
rect 3237 23780 3249 23783
rect 2746 23752 3249 23780
rect 2317 23715 2375 23721
rect 2317 23681 2329 23715
rect 2363 23712 2375 23715
rect 2746 23712 2774 23752
rect 3237 23749 3249 23752
rect 3283 23780 3295 23783
rect 3326 23780 3332 23792
rect 3283 23752 3332 23780
rect 3283 23749 3295 23752
rect 3237 23743 3295 23749
rect 3326 23740 3332 23752
rect 3384 23740 3390 23792
rect 5074 23740 5080 23792
rect 5132 23740 5138 23792
rect 5534 23780 5540 23792
rect 5495 23752 5540 23780
rect 5534 23740 5540 23752
rect 5592 23740 5598 23792
rect 8938 23740 8944 23792
rect 8996 23740 9002 23792
rect 9306 23740 9312 23792
rect 9364 23780 9370 23792
rect 9401 23783 9459 23789
rect 9401 23780 9413 23783
rect 9364 23752 9413 23780
rect 9364 23740 9370 23752
rect 9401 23749 9413 23752
rect 9447 23749 9459 23783
rect 9401 23743 9459 23749
rect 2363 23684 2774 23712
rect 2363 23681 2375 23684
rect 2317 23675 2375 23681
rect 6638 23672 6644 23724
rect 6696 23712 6702 23724
rect 6696 23684 7972 23712
rect 6696 23672 6702 23684
rect 2130 23644 2136 23656
rect 2091 23616 2136 23644
rect 2130 23604 2136 23616
rect 2188 23604 2194 23656
rect 2225 23647 2283 23653
rect 2225 23613 2237 23647
rect 2271 23644 2283 23647
rect 2406 23644 2412 23656
rect 2271 23616 2412 23644
rect 2271 23613 2283 23616
rect 2225 23607 2283 23613
rect 2406 23604 2412 23616
rect 2464 23644 2470 23656
rect 2590 23644 2596 23656
rect 2464 23616 2596 23644
rect 2464 23604 2470 23616
rect 2590 23604 2596 23616
rect 2648 23604 2654 23656
rect 2682 23604 2688 23656
rect 2740 23644 2746 23656
rect 7944 23653 7972 23684
rect 4065 23647 4123 23653
rect 4065 23644 4077 23647
rect 2740 23616 4077 23644
rect 2740 23604 2746 23616
rect 4065 23613 4077 23616
rect 4111 23613 4123 23647
rect 4065 23607 4123 23613
rect 5813 23647 5871 23653
rect 5813 23613 5825 23647
rect 5859 23644 5871 23647
rect 7929 23647 7987 23653
rect 5859 23616 6684 23644
rect 5859 23613 5871 23616
rect 5813 23607 5871 23613
rect 6656 23588 6684 23616
rect 7929 23613 7941 23647
rect 7975 23613 7987 23647
rect 7929 23607 7987 23613
rect 9677 23647 9735 23653
rect 9677 23613 9689 23647
rect 9723 23644 9735 23647
rect 10134 23644 10140 23656
rect 9723 23616 10140 23644
rect 9723 23613 9735 23616
rect 9677 23607 9735 23613
rect 6638 23536 6644 23588
rect 6696 23576 6702 23588
rect 6696 23548 8064 23576
rect 6696 23536 6702 23548
rect 2314 23468 2320 23520
rect 2372 23508 2378 23520
rect 2685 23511 2743 23517
rect 2685 23508 2697 23511
rect 2372 23480 2697 23508
rect 2372 23468 2378 23480
rect 2685 23477 2697 23480
rect 2731 23477 2743 23511
rect 8036 23508 8064 23548
rect 9692 23508 9720 23607
rect 10134 23604 10140 23616
rect 10192 23604 10198 23656
rect 8036 23480 9720 23508
rect 2685 23471 2743 23477
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 4062 23304 4068 23316
rect 1872 23276 4068 23304
rect 1872 23109 1900 23276
rect 4062 23264 4068 23276
rect 4120 23264 4126 23316
rect 10226 23264 10232 23316
rect 10284 23304 10290 23316
rect 10689 23307 10747 23313
rect 10689 23304 10701 23307
rect 10284 23276 10701 23304
rect 10284 23264 10290 23276
rect 10689 23273 10701 23276
rect 10735 23273 10747 23307
rect 10689 23267 10747 23273
rect 2501 23239 2559 23245
rect 2501 23205 2513 23239
rect 2547 23205 2559 23239
rect 2501 23199 2559 23205
rect 2516 23168 2544 23199
rect 2590 23196 2596 23248
rect 2648 23236 2654 23248
rect 4893 23239 4951 23245
rect 4893 23236 4905 23239
rect 2648 23208 4905 23236
rect 2648 23196 2654 23208
rect 4893 23205 4905 23208
rect 4939 23205 4951 23239
rect 4893 23199 4951 23205
rect 6365 23171 6423 23177
rect 6365 23168 6377 23171
rect 2516 23140 6377 23168
rect 6365 23137 6377 23140
rect 6411 23137 6423 23171
rect 6638 23168 6644 23180
rect 6599 23140 6644 23168
rect 6365 23131 6423 23137
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 11606 23128 11612 23180
rect 11664 23168 11670 23180
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 11664 23140 12173 23168
rect 11664 23128 11670 23140
rect 12161 23137 12173 23140
rect 12207 23137 12219 23171
rect 12161 23131 12219 23137
rect 57974 23128 57980 23180
rect 58032 23168 58038 23180
rect 58069 23171 58127 23177
rect 58069 23168 58081 23171
rect 58032 23140 58081 23168
rect 58032 23128 58038 23140
rect 58069 23137 58081 23140
rect 58115 23137 58127 23171
rect 58069 23131 58127 23137
rect 1857 23103 1915 23109
rect 1857 23069 1869 23103
rect 1903 23069 1915 23103
rect 2314 23100 2320 23112
rect 2275 23072 2320 23100
rect 1857 23063 1915 23069
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 2682 23060 2688 23112
rect 2740 23100 2746 23112
rect 2961 23103 3019 23109
rect 2961 23100 2973 23103
rect 2740 23072 2973 23100
rect 2740 23060 2746 23072
rect 2961 23069 2973 23072
rect 3007 23069 3019 23103
rect 2961 23063 3019 23069
rect 12434 23060 12440 23112
rect 12492 23100 12498 23112
rect 12492 23072 12537 23100
rect 12492 23060 12498 23072
rect 53098 23060 53104 23112
rect 53156 23100 53162 23112
rect 57793 23103 57851 23109
rect 57793 23100 57805 23103
rect 53156 23072 57805 23100
rect 53156 23060 53162 23072
rect 57793 23069 57805 23072
rect 57839 23069 57851 23103
rect 57793 23063 57851 23069
rect 5350 22992 5356 23044
rect 5408 22992 5414 23044
rect 11882 23032 11888 23044
rect 11730 23004 11888 23032
rect 11882 22992 11888 23004
rect 11940 22992 11946 23044
rect 1670 22964 1676 22976
rect 1631 22936 1676 22964
rect 1670 22924 1676 22936
rect 1728 22924 1734 22976
rect 3142 22964 3148 22976
rect 3103 22936 3148 22964
rect 3142 22924 3148 22936
rect 3200 22924 3206 22976
rect 4062 22964 4068 22976
rect 3975 22936 4068 22964
rect 4062 22924 4068 22936
rect 4120 22964 4126 22976
rect 10594 22964 10600 22976
rect 4120 22936 10600 22964
rect 4120 22924 4126 22936
rect 10594 22924 10600 22936
rect 10652 22924 10658 22976
rect 18414 22964 18420 22976
rect 18375 22936 18420 22964
rect 18414 22924 18420 22936
rect 18472 22924 18478 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 2225 22763 2283 22769
rect 2225 22729 2237 22763
rect 2271 22760 2283 22763
rect 2498 22760 2504 22772
rect 2271 22732 2504 22760
rect 2271 22729 2283 22732
rect 2225 22723 2283 22729
rect 2498 22720 2504 22732
rect 2556 22720 2562 22772
rect 2682 22760 2688 22772
rect 2643 22732 2688 22760
rect 2682 22720 2688 22732
rect 2740 22720 2746 22772
rect 3234 22760 3240 22772
rect 3195 22732 3240 22760
rect 3234 22720 3240 22732
rect 3292 22720 3298 22772
rect 8389 22763 8447 22769
rect 8389 22729 8401 22763
rect 8435 22760 8447 22763
rect 8570 22760 8576 22772
rect 8435 22732 8576 22760
rect 8435 22729 8447 22732
rect 8389 22723 8447 22729
rect 8570 22720 8576 22732
rect 8628 22720 8634 22772
rect 11698 22720 11704 22772
rect 11756 22760 11762 22772
rect 11882 22760 11888 22772
rect 11756 22732 11888 22760
rect 11756 22720 11762 22732
rect 11882 22720 11888 22732
rect 11940 22760 11946 22772
rect 14182 22760 14188 22772
rect 11940 22732 12848 22760
rect 11940 22720 11946 22732
rect 2317 22695 2375 22701
rect 2317 22661 2329 22695
rect 2363 22692 2375 22695
rect 3252 22692 3280 22720
rect 2363 22664 3280 22692
rect 2363 22661 2375 22664
rect 2317 22655 2375 22661
rect 2130 22556 2136 22568
rect 2091 22528 2136 22556
rect 2130 22516 2136 22528
rect 2188 22516 2194 22568
rect 3252 22556 3280 22664
rect 5074 22652 5080 22704
rect 5132 22692 5138 22704
rect 5350 22692 5356 22704
rect 5132 22664 5356 22692
rect 5132 22652 5138 22664
rect 5350 22652 5356 22664
rect 5408 22692 5414 22704
rect 12710 22692 12716 22704
rect 5408 22664 8694 22692
rect 12671 22664 12716 22692
rect 5408 22652 5414 22664
rect 12710 22652 12716 22664
rect 12768 22652 12774 22704
rect 12820 22692 12848 22732
rect 13096 22732 13860 22760
rect 14143 22732 14188 22760
rect 13096 22692 13124 22732
rect 12820 22664 13202 22692
rect 13832 22636 13860 22732
rect 14182 22720 14188 22732
rect 14240 22720 14246 22772
rect 18785 22763 18843 22769
rect 18785 22729 18797 22763
rect 18831 22729 18843 22763
rect 18785 22723 18843 22729
rect 10134 22584 10140 22636
rect 10192 22624 10198 22636
rect 12434 22624 12440 22636
rect 10192 22596 10237 22624
rect 12395 22596 12440 22624
rect 10192 22584 10198 22596
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 13814 22584 13820 22636
rect 13872 22584 13878 22636
rect 18325 22627 18383 22633
rect 18325 22593 18337 22627
rect 18371 22624 18383 22627
rect 18800 22624 18828 22723
rect 56778 22720 56784 22772
rect 56836 22760 56842 22772
rect 58161 22763 58219 22769
rect 58161 22760 58173 22763
rect 56836 22732 58173 22760
rect 56836 22720 56842 22732
rect 58161 22729 58173 22732
rect 58207 22729 58219 22763
rect 58161 22723 58219 22729
rect 19153 22695 19211 22701
rect 19153 22661 19165 22695
rect 19199 22692 19211 22695
rect 19242 22692 19248 22704
rect 19199 22664 19248 22692
rect 19199 22661 19211 22664
rect 19153 22655 19211 22661
rect 19242 22652 19248 22664
rect 19300 22652 19306 22704
rect 18371 22596 18828 22624
rect 57517 22627 57575 22633
rect 18371 22593 18383 22596
rect 18325 22587 18383 22593
rect 57517 22593 57529 22627
rect 57563 22624 57575 22627
rect 58342 22624 58348 22636
rect 57563 22596 58348 22624
rect 57563 22593 57575 22596
rect 57517 22587 57575 22593
rect 58342 22584 58348 22596
rect 58400 22584 58406 22636
rect 3326 22556 3332 22568
rect 3252 22528 3332 22556
rect 3326 22516 3332 22528
rect 3384 22516 3390 22568
rect 8202 22516 8208 22568
rect 8260 22556 8266 22568
rect 9861 22559 9919 22565
rect 9861 22556 9873 22559
rect 8260 22528 9873 22556
rect 8260 22516 8266 22528
rect 9861 22525 9873 22528
rect 9907 22525 9919 22559
rect 9861 22519 9919 22525
rect 18414 22516 18420 22568
rect 18472 22556 18478 22568
rect 19245 22559 19303 22565
rect 19245 22556 19257 22559
rect 18472 22528 19257 22556
rect 18472 22516 18478 22528
rect 19245 22525 19257 22528
rect 19291 22525 19303 22559
rect 19245 22519 19303 22525
rect 19429 22559 19487 22565
rect 19429 22525 19441 22559
rect 19475 22556 19487 22559
rect 19475 22528 20116 22556
rect 19475 22525 19487 22528
rect 19429 22519 19487 22525
rect 17402 22448 17408 22500
rect 17460 22488 17466 22500
rect 19444 22488 19472 22519
rect 17460 22460 19472 22488
rect 17460 22448 17466 22460
rect 15654 22380 15660 22432
rect 15712 22420 15718 22432
rect 20088 22429 20116 22528
rect 18141 22423 18199 22429
rect 18141 22420 18153 22423
rect 15712 22392 18153 22420
rect 15712 22380 15718 22392
rect 18141 22389 18153 22392
rect 18187 22389 18199 22423
rect 18141 22383 18199 22389
rect 20073 22423 20131 22429
rect 20073 22389 20085 22423
rect 20119 22420 20131 22423
rect 20346 22420 20352 22432
rect 20119 22392 20352 22420
rect 20119 22389 20131 22392
rect 20073 22383 20131 22389
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1670 22216 1676 22228
rect 1631 22188 1676 22216
rect 1670 22176 1676 22188
rect 1728 22176 1734 22228
rect 3142 22176 3148 22228
rect 3200 22216 3206 22228
rect 6285 22219 6343 22225
rect 6285 22216 6297 22219
rect 3200 22188 6297 22216
rect 3200 22176 3206 22188
rect 6285 22185 6297 22188
rect 6331 22185 6343 22219
rect 6285 22179 6343 22185
rect 15276 22219 15334 22225
rect 15276 22185 15288 22219
rect 15322 22216 15334 22219
rect 15930 22216 15936 22228
rect 15322 22188 15936 22216
rect 15322 22185 15334 22188
rect 15276 22179 15334 22185
rect 15930 22176 15936 22188
rect 15988 22176 15994 22228
rect 2130 22040 2136 22092
rect 2188 22080 2194 22092
rect 2777 22083 2835 22089
rect 2777 22080 2789 22083
rect 2188 22052 2789 22080
rect 2188 22040 2194 22052
rect 2777 22049 2789 22052
rect 2823 22049 2835 22083
rect 16758 22080 16764 22092
rect 16719 22052 16764 22080
rect 2777 22043 2835 22049
rect 16758 22040 16764 22052
rect 16816 22040 16822 22092
rect 1854 22012 1860 22024
rect 1815 21984 1860 22012
rect 1854 21972 1860 21984
rect 1912 21972 1918 22024
rect 6549 22015 6607 22021
rect 6549 21981 6561 22015
rect 6595 22012 6607 22015
rect 6638 22012 6644 22024
rect 6595 21984 6644 22012
rect 6595 21981 6607 21984
rect 6549 21975 6607 21981
rect 2746 21916 4844 21944
rect 2498 21836 2504 21888
rect 2556 21876 2562 21888
rect 2746 21876 2774 21916
rect 4816 21885 4844 21916
rect 5258 21904 5264 21956
rect 5316 21904 5322 21956
rect 5994 21904 6000 21956
rect 6052 21944 6058 21956
rect 6564 21944 6592 21975
rect 6638 21972 6644 21984
rect 6696 21972 6702 22024
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 21981 15071 22015
rect 15013 21975 15071 21981
rect 57701 22015 57759 22021
rect 57701 21981 57713 22015
rect 57747 22012 57759 22015
rect 58342 22012 58348 22024
rect 57747 21984 58348 22012
rect 57747 21981 57759 21984
rect 57701 21975 57759 21981
rect 6052 21916 6592 21944
rect 15028 21944 15056 21975
rect 58342 21972 58348 21984
rect 58400 21972 58406 22024
rect 15194 21944 15200 21956
rect 15028 21916 15200 21944
rect 6052 21904 6058 21916
rect 15194 21904 15200 21916
rect 15252 21904 15258 21956
rect 16022 21904 16028 21956
rect 16080 21904 16086 21956
rect 2556 21848 2774 21876
rect 4801 21879 4859 21885
rect 2556 21836 2562 21848
rect 4801 21845 4813 21879
rect 4847 21845 4859 21879
rect 4801 21839 4859 21845
rect 18693 21879 18751 21885
rect 18693 21845 18705 21879
rect 18739 21876 18751 21879
rect 19242 21876 19248 21888
rect 18739 21848 19248 21876
rect 18739 21845 18751 21848
rect 18693 21839 18751 21845
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 58161 21879 58219 21885
rect 58161 21845 58173 21879
rect 58207 21876 58219 21879
rect 58710 21876 58716 21888
rect 58207 21848 58716 21876
rect 58207 21845 58219 21848
rect 58161 21839 58219 21845
rect 58710 21836 58716 21848
rect 58768 21836 58774 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 2866 21632 2872 21684
rect 2924 21672 2930 21684
rect 16206 21672 16212 21684
rect 2924 21644 16212 21672
rect 2924 21632 2930 21644
rect 16206 21632 16212 21644
rect 16264 21632 16270 21684
rect 58158 21672 58164 21684
rect 58119 21644 58164 21672
rect 58158 21632 58164 21644
rect 58216 21632 58222 21684
rect 13814 21564 13820 21616
rect 13872 21604 13878 21616
rect 13872 21576 14122 21604
rect 13872 21564 13878 21576
rect 15194 21564 15200 21616
rect 15252 21604 15258 21616
rect 15252 21576 15608 21604
rect 15252 21564 15258 21576
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21536 1915 21539
rect 2590 21536 2596 21548
rect 1903 21508 2596 21536
rect 1903 21505 1915 21508
rect 1857 21499 1915 21505
rect 2590 21496 2596 21508
rect 2648 21496 2654 21548
rect 15580 21545 15608 21576
rect 17586 21564 17592 21616
rect 17644 21604 17650 21616
rect 19337 21607 19395 21613
rect 19337 21604 19349 21607
rect 17644 21576 19349 21604
rect 17644 21564 17650 21576
rect 19337 21573 19349 21576
rect 19383 21573 19395 21607
rect 19337 21567 19395 21573
rect 15565 21539 15623 21545
rect 15565 21505 15577 21539
rect 15611 21505 15623 21539
rect 15565 21499 15623 21505
rect 19613 21539 19671 21545
rect 19613 21505 19625 21539
rect 19659 21536 19671 21539
rect 20162 21536 20168 21548
rect 19659 21508 20168 21536
rect 19659 21505 19671 21508
rect 19613 21499 19671 21505
rect 20162 21496 20168 21508
rect 20220 21496 20226 21548
rect 57517 21539 57575 21545
rect 57517 21505 57529 21539
rect 57563 21536 57575 21539
rect 58342 21536 58348 21548
rect 57563 21508 58348 21536
rect 57563 21505 57575 21508
rect 57517 21499 57575 21505
rect 58342 21496 58348 21508
rect 58400 21496 58406 21548
rect 11790 21428 11796 21480
rect 11848 21468 11854 21480
rect 13814 21468 13820 21480
rect 11848 21440 13820 21468
rect 11848 21428 11854 21440
rect 13814 21428 13820 21440
rect 13872 21428 13878 21480
rect 15286 21468 15292 21480
rect 15247 21440 15292 21468
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 1670 21400 1676 21412
rect 1631 21372 1676 21400
rect 1670 21360 1676 21372
rect 1728 21360 1734 21412
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 2869 21335 2927 21341
rect 2869 21332 2881 21335
rect 2832 21304 2881 21332
rect 2832 21292 2838 21304
rect 2869 21301 2881 21304
rect 2915 21332 2927 21335
rect 2958 21332 2964 21344
rect 2915 21304 2964 21332
rect 2915 21301 2927 21304
rect 2869 21295 2927 21301
rect 2958 21292 2964 21304
rect 3016 21292 3022 21344
rect 13817 21335 13875 21341
rect 13817 21301 13829 21335
rect 13863 21332 13875 21335
rect 14090 21332 14096 21344
rect 13863 21304 14096 21332
rect 13863 21301 13875 21304
rect 13817 21295 13875 21301
rect 14090 21292 14096 21304
rect 14148 21292 14154 21344
rect 20162 21332 20168 21344
rect 20123 21304 20168 21332
rect 20162 21292 20168 21304
rect 20220 21292 20226 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 11974 21128 11980 21140
rect 11935 21100 11980 21128
rect 11974 21088 11980 21100
rect 12032 21088 12038 21140
rect 14366 21088 14372 21140
rect 14424 21128 14430 21140
rect 17037 21131 17095 21137
rect 17037 21128 17049 21131
rect 14424 21100 17049 21128
rect 14424 21088 14430 21100
rect 17037 21097 17049 21100
rect 17083 21097 17095 21131
rect 18230 21128 18236 21140
rect 18191 21100 18236 21128
rect 17037 21091 17095 21097
rect 18230 21088 18236 21100
rect 18288 21128 18294 21140
rect 58161 21131 58219 21137
rect 18288 21100 19932 21128
rect 18288 21088 18294 21100
rect 2133 20995 2191 21001
rect 2133 20961 2145 20995
rect 2179 20992 2191 20995
rect 2958 20992 2964 21004
rect 2179 20964 2964 20992
rect 2179 20961 2191 20964
rect 2133 20955 2191 20961
rect 2958 20952 2964 20964
rect 3016 20952 3022 21004
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 13725 20995 13783 21001
rect 13725 20992 13737 20995
rect 12492 20964 13737 20992
rect 12492 20952 12498 20964
rect 13725 20961 13737 20964
rect 13771 20992 13783 20995
rect 15194 20992 15200 21004
rect 13771 20964 15200 20992
rect 13771 20961 13783 20964
rect 13725 20955 13783 20961
rect 15194 20952 15200 20964
rect 15252 20992 15258 21004
rect 15289 20995 15347 21001
rect 15289 20992 15301 20995
rect 15252 20964 15301 20992
rect 15252 20952 15258 20964
rect 15289 20961 15301 20964
rect 15335 20961 15347 20995
rect 15562 20992 15568 21004
rect 15523 20964 15568 20992
rect 15289 20955 15347 20961
rect 15562 20952 15568 20964
rect 15620 20952 15626 21004
rect 19904 21001 19932 21100
rect 58161 21097 58173 21131
rect 58207 21128 58219 21131
rect 58250 21128 58256 21140
rect 58207 21100 58256 21128
rect 58207 21097 58219 21100
rect 58161 21091 58219 21097
rect 58250 21088 58256 21100
rect 58308 21088 58314 21140
rect 19889 20995 19947 21001
rect 19889 20961 19901 20995
rect 19935 20961 19947 20995
rect 19889 20955 19947 20961
rect 20073 20995 20131 21001
rect 20073 20961 20085 20995
rect 20119 20992 20131 20995
rect 20162 20992 20168 21004
rect 20119 20964 20168 20992
rect 20119 20961 20131 20964
rect 20073 20955 20131 20961
rect 20162 20952 20168 20964
rect 20220 20992 20226 21004
rect 20622 20992 20628 21004
rect 20220 20964 20628 20992
rect 20220 20952 20226 20964
rect 20622 20952 20628 20964
rect 20680 20952 20686 21004
rect 2317 20927 2375 20933
rect 2317 20893 2329 20927
rect 2363 20924 2375 20927
rect 3050 20924 3056 20936
rect 2363 20896 3056 20924
rect 2363 20893 2375 20896
rect 2317 20887 2375 20893
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 12342 20884 12348 20936
rect 12400 20884 12406 20936
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20924 18935 20927
rect 19426 20924 19432 20936
rect 18923 20896 19432 20924
rect 18923 20893 18935 20896
rect 18877 20887 18935 20893
rect 19426 20884 19432 20896
rect 19484 20924 19490 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19484 20896 19809 20924
rect 19484 20884 19490 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 57701 20927 57759 20933
rect 57701 20893 57713 20927
rect 57747 20924 57759 20927
rect 58342 20924 58348 20936
rect 57747 20896 58348 20924
rect 57747 20893 57759 20896
rect 57701 20887 57759 20893
rect 58342 20884 58348 20896
rect 58400 20884 58406 20936
rect 1854 20816 1860 20868
rect 1912 20856 1918 20868
rect 2225 20859 2283 20865
rect 2225 20856 2237 20859
rect 1912 20828 2237 20856
rect 1912 20816 1918 20828
rect 2225 20825 2237 20828
rect 2271 20856 2283 20859
rect 4154 20856 4160 20868
rect 2271 20828 4160 20856
rect 2271 20825 2283 20828
rect 2225 20819 2283 20825
rect 4154 20816 4160 20828
rect 4212 20816 4218 20868
rect 13354 20816 13360 20868
rect 13412 20856 13418 20868
rect 13449 20859 13507 20865
rect 13449 20856 13461 20859
rect 13412 20828 13461 20856
rect 13412 20816 13418 20828
rect 13449 20825 13461 20828
rect 13495 20825 13507 20859
rect 13449 20819 13507 20825
rect 16022 20816 16028 20868
rect 16080 20816 16086 20868
rect 2682 20788 2688 20800
rect 2643 20760 2688 20788
rect 2682 20748 2688 20760
rect 2740 20748 2746 20800
rect 3050 20748 3056 20800
rect 3108 20788 3114 20800
rect 3237 20791 3295 20797
rect 3237 20788 3249 20791
rect 3108 20760 3249 20788
rect 3108 20748 3114 20760
rect 3237 20757 3249 20760
rect 3283 20788 3295 20791
rect 3418 20788 3424 20800
rect 3283 20760 3424 20788
rect 3283 20757 3295 20760
rect 3237 20751 3295 20757
rect 3418 20748 3424 20760
rect 3476 20788 3482 20800
rect 3786 20788 3792 20800
rect 3476 20760 3792 20788
rect 3476 20748 3482 20760
rect 3786 20748 3792 20760
rect 3844 20748 3850 20800
rect 4798 20748 4804 20800
rect 4856 20788 4862 20800
rect 10778 20788 10784 20800
rect 4856 20760 10784 20788
rect 4856 20748 4862 20760
rect 10778 20748 10784 20760
rect 10836 20748 10842 20800
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 19429 20791 19487 20797
rect 19429 20788 19441 20791
rect 19392 20760 19441 20788
rect 19392 20748 19398 20760
rect 19429 20757 19441 20760
rect 19475 20757 19487 20791
rect 20622 20788 20628 20800
rect 20583 20760 20628 20788
rect 19429 20751 19487 20757
rect 20622 20748 20628 20760
rect 20680 20748 20686 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 1670 20584 1676 20596
rect 1631 20556 1676 20584
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 4249 20587 4307 20593
rect 4249 20553 4261 20587
rect 4295 20584 4307 20587
rect 4706 20584 4712 20596
rect 4295 20556 4712 20584
rect 4295 20553 4307 20556
rect 4249 20547 4307 20553
rect 4706 20544 4712 20556
rect 4764 20544 4770 20596
rect 10870 20584 10876 20596
rect 10831 20556 10876 20584
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 11606 20544 11612 20596
rect 11664 20584 11670 20596
rect 14918 20584 14924 20596
rect 11664 20556 14924 20584
rect 11664 20544 11670 20556
rect 14918 20544 14924 20556
rect 14976 20544 14982 20596
rect 18782 20544 18788 20596
rect 18840 20584 18846 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 18840 20556 19441 20584
rect 18840 20544 18846 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 5258 20476 5264 20528
rect 5316 20476 5322 20528
rect 8938 20476 8944 20528
rect 8996 20516 9002 20528
rect 8996 20488 9890 20516
rect 8996 20476 9002 20488
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20448 1915 20451
rect 2130 20448 2136 20460
rect 1903 20420 2136 20448
rect 1903 20417 1915 20420
rect 1857 20411 1915 20417
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 2317 20451 2375 20457
rect 2317 20417 2329 20451
rect 2363 20448 2375 20451
rect 2682 20448 2688 20460
rect 2363 20420 2688 20448
rect 2363 20417 2375 20420
rect 2317 20411 2375 20417
rect 2682 20408 2688 20420
rect 2740 20408 2746 20460
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 19334 20448 19340 20460
rect 18739 20420 19340 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 19518 20448 19524 20460
rect 19479 20420 19524 20448
rect 19518 20408 19524 20420
rect 19576 20408 19582 20460
rect 3878 20340 3884 20392
rect 3936 20380 3942 20392
rect 5721 20383 5779 20389
rect 5721 20380 5733 20383
rect 3936 20352 5733 20380
rect 3936 20340 3942 20352
rect 5721 20349 5733 20352
rect 5767 20349 5779 20383
rect 5994 20380 6000 20392
rect 5955 20352 6000 20380
rect 5721 20343 5779 20349
rect 5994 20340 6000 20352
rect 6052 20340 6058 20392
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 9125 20383 9183 20389
rect 9125 20380 9137 20383
rect 8352 20352 9137 20380
rect 8352 20340 8358 20352
rect 9125 20349 9137 20352
rect 9171 20349 9183 20383
rect 9125 20343 9183 20349
rect 9401 20383 9459 20389
rect 9401 20349 9413 20383
rect 9447 20380 9459 20383
rect 9766 20380 9772 20392
rect 9447 20352 9772 20380
rect 9447 20349 9459 20352
rect 9401 20343 9459 20349
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 19245 20383 19303 20389
rect 19245 20349 19257 20383
rect 19291 20380 19303 20383
rect 19291 20352 20484 20380
rect 19291 20349 19303 20352
rect 19245 20343 19303 20349
rect 2501 20315 2559 20321
rect 2501 20281 2513 20315
rect 2547 20312 2559 20315
rect 4706 20312 4712 20324
rect 2547 20284 4712 20312
rect 2547 20281 2559 20284
rect 2501 20275 2559 20281
rect 4706 20272 4712 20284
rect 4764 20272 4770 20324
rect 20456 20256 20484 20352
rect 16022 20204 16028 20256
rect 16080 20244 16086 20256
rect 18509 20247 18567 20253
rect 18509 20244 18521 20247
rect 16080 20216 18521 20244
rect 16080 20204 16086 20216
rect 18509 20213 18521 20216
rect 18555 20213 18567 20247
rect 18509 20207 18567 20213
rect 19889 20247 19947 20253
rect 19889 20213 19901 20247
rect 19935 20244 19947 20247
rect 19978 20244 19984 20256
rect 19935 20216 19984 20244
rect 19935 20213 19947 20216
rect 19889 20207 19947 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 20438 20244 20444 20256
rect 20399 20216 20444 20244
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20040 17187 20043
rect 18414 20040 18420 20052
rect 17175 20012 18420 20040
rect 17175 20009 17187 20012
rect 17129 20003 17187 20009
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 18782 20040 18788 20052
rect 18743 20012 18788 20040
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15381 19907 15439 19913
rect 15381 19904 15393 19907
rect 15252 19876 15393 19904
rect 15252 19864 15258 19876
rect 15381 19873 15393 19876
rect 15427 19873 15439 19907
rect 15654 19904 15660 19916
rect 15615 19876 15660 19904
rect 15381 19867 15439 19873
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19836 1915 19839
rect 2038 19836 2044 19848
rect 1903 19808 2044 19836
rect 1903 19805 1915 19808
rect 1857 19799 1915 19805
rect 2038 19796 2044 19808
rect 2096 19796 2102 19848
rect 57701 19839 57759 19845
rect 57701 19805 57713 19839
rect 57747 19836 57759 19839
rect 58342 19836 58348 19848
rect 57747 19808 58348 19836
rect 57747 19805 57759 19808
rect 57701 19799 57759 19805
rect 58342 19796 58348 19808
rect 58400 19796 58406 19848
rect 5718 19768 5724 19780
rect 5631 19740 5724 19768
rect 5718 19728 5724 19740
rect 5776 19768 5782 19780
rect 6365 19771 6423 19777
rect 6365 19768 6377 19771
rect 5776 19740 6377 19768
rect 5776 19728 5782 19740
rect 6365 19737 6377 19740
rect 6411 19737 6423 19771
rect 6365 19731 6423 19737
rect 16114 19728 16120 19780
rect 16172 19728 16178 19780
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 5813 19703 5871 19709
rect 5813 19700 5825 19703
rect 5316 19672 5825 19700
rect 5316 19660 5322 19672
rect 5813 19669 5825 19672
rect 5859 19669 5871 19703
rect 19518 19700 19524 19712
rect 19431 19672 19524 19700
rect 5813 19663 5871 19669
rect 19518 19660 19524 19672
rect 19576 19700 19582 19712
rect 20530 19700 20536 19712
rect 19576 19672 20536 19700
rect 19576 19660 19582 19672
rect 20530 19660 20536 19672
rect 20588 19660 20594 19712
rect 58066 19660 58072 19712
rect 58124 19700 58130 19712
rect 58161 19703 58219 19709
rect 58161 19700 58173 19703
rect 58124 19672 58173 19700
rect 58124 19660 58130 19672
rect 58161 19669 58173 19672
rect 58207 19669 58219 19703
rect 58161 19663 58219 19669
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 4249 19499 4307 19505
rect 4249 19496 4261 19499
rect 4212 19468 4261 19496
rect 4212 19456 4218 19468
rect 4249 19465 4261 19468
rect 4295 19465 4307 19499
rect 4249 19459 4307 19465
rect 8754 19456 8760 19508
rect 8812 19496 8818 19508
rect 9493 19499 9551 19505
rect 9493 19496 9505 19499
rect 8812 19468 9505 19496
rect 8812 19456 8818 19468
rect 9493 19465 9505 19468
rect 9539 19465 9551 19499
rect 14642 19496 14648 19508
rect 14603 19468 14648 19496
rect 9493 19459 9551 19465
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 56594 19456 56600 19508
rect 56652 19496 56658 19508
rect 58161 19499 58219 19505
rect 58161 19496 58173 19499
rect 56652 19468 58173 19496
rect 56652 19456 56658 19468
rect 58161 19465 58173 19468
rect 58207 19465 58219 19499
rect 58161 19459 58219 19465
rect 5258 19388 5264 19440
rect 5316 19388 5322 19440
rect 8294 19428 8300 19440
rect 7760 19400 8300 19428
rect 1857 19363 1915 19369
rect 1857 19329 1869 19363
rect 1903 19360 1915 19363
rect 2222 19360 2228 19372
rect 1903 19332 2228 19360
rect 1903 19329 1915 19332
rect 1857 19323 1915 19329
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 5994 19320 6000 19372
rect 6052 19360 6058 19372
rect 7760 19369 7788 19400
rect 8294 19388 8300 19400
rect 8352 19388 8358 19440
rect 9030 19388 9036 19440
rect 9088 19388 9094 19440
rect 16114 19428 16120 19440
rect 14398 19414 16120 19428
rect 14384 19400 16120 19414
rect 7745 19363 7803 19369
rect 7745 19360 7757 19363
rect 6052 19332 7757 19360
rect 6052 19320 6058 19332
rect 7745 19329 7757 19332
rect 7791 19329 7803 19363
rect 7745 19323 7803 19329
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12618 19360 12624 19372
rect 12492 19332 12624 19360
rect 12492 19320 12498 19332
rect 12618 19320 12624 19332
rect 12676 19360 12682 19372
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12676 19332 12909 19360
rect 12676 19320 12682 19332
rect 12897 19329 12909 19332
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 4706 19252 4712 19304
rect 4764 19292 4770 19304
rect 5721 19295 5779 19301
rect 5721 19292 5733 19295
rect 4764 19264 5733 19292
rect 4764 19252 4770 19264
rect 5721 19261 5733 19264
rect 5767 19261 5779 19295
rect 5721 19255 5779 19261
rect 8021 19295 8079 19301
rect 8021 19261 8033 19295
rect 8067 19292 8079 19295
rect 8110 19292 8116 19304
rect 8067 19264 8116 19292
rect 8067 19261 8079 19264
rect 8021 19255 8079 19261
rect 8110 19252 8116 19264
rect 8168 19252 8174 19304
rect 13170 19292 13176 19304
rect 13131 19264 13176 19292
rect 13170 19252 13176 19264
rect 13228 19252 13234 19304
rect 1670 19156 1676 19168
rect 1631 19128 1676 19156
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 12342 19116 12348 19168
rect 12400 19156 12406 19168
rect 14384 19156 14412 19400
rect 16114 19388 16120 19400
rect 16172 19388 16178 19440
rect 58342 19360 58348 19372
rect 58303 19332 58348 19360
rect 58342 19320 58348 19332
rect 58400 19320 58406 19372
rect 57238 19292 57244 19304
rect 57199 19264 57244 19292
rect 57238 19252 57244 19264
rect 57296 19252 57302 19304
rect 57514 19292 57520 19304
rect 57475 19264 57520 19292
rect 57514 19252 57520 19264
rect 57572 19252 57578 19304
rect 12400 19128 14412 19156
rect 12400 19116 12406 19128
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 10873 18955 10931 18961
rect 10873 18952 10885 18955
rect 7708 18924 10885 18952
rect 7708 18912 7714 18924
rect 10873 18921 10885 18924
rect 10919 18921 10931 18955
rect 58342 18952 58348 18964
rect 58303 18924 58348 18952
rect 10873 18915 10931 18921
rect 1854 18748 1860 18760
rect 1815 18720 1860 18748
rect 1854 18708 1860 18720
rect 1912 18708 1918 18760
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18748 2375 18751
rect 2682 18748 2688 18760
rect 2363 18720 2688 18748
rect 2363 18717 2375 18720
rect 2317 18711 2375 18717
rect 2682 18708 2688 18720
rect 2740 18708 2746 18760
rect 1670 18612 1676 18624
rect 1631 18584 1676 18612
rect 1670 18572 1676 18584
rect 1728 18572 1734 18624
rect 2498 18612 2504 18624
rect 2459 18584 2504 18612
rect 2498 18572 2504 18584
rect 2556 18572 2562 18624
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 10888 18612 10916 18915
rect 58342 18912 58348 18924
rect 58400 18912 58406 18964
rect 20165 18887 20223 18893
rect 20165 18884 20177 18887
rect 16546 18856 20177 18884
rect 12618 18816 12624 18828
rect 12579 18788 12624 18816
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 15102 18816 15108 18828
rect 15063 18788 15108 18816
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 15381 18819 15439 18825
rect 15381 18785 15393 18819
rect 15427 18816 15439 18819
rect 16546 18816 16574 18856
rect 20165 18853 20177 18856
rect 20211 18853 20223 18887
rect 20165 18847 20223 18853
rect 17126 18816 17132 18828
rect 15427 18788 16574 18816
rect 17087 18788 17132 18816
rect 15427 18785 15439 18788
rect 15381 18779 15439 18785
rect 17126 18776 17132 18788
rect 17184 18776 17190 18828
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18748 19763 18751
rect 19978 18748 19984 18760
rect 19751 18720 19984 18748
rect 19751 18717 19763 18720
rect 19705 18711 19763 18717
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20254 18708 20260 18760
rect 20312 18748 20318 18760
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 20312 18720 20361 18748
rect 20312 18708 20318 18720
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 12250 18680 12256 18692
rect 11914 18652 12256 18680
rect 12250 18640 12256 18652
rect 12308 18640 12314 18692
rect 12345 18683 12403 18689
rect 12345 18649 12357 18683
rect 12391 18680 12403 18683
rect 15286 18680 15292 18692
rect 12391 18652 15292 18680
rect 12391 18649 12403 18652
rect 12345 18643 12403 18649
rect 15286 18640 15292 18652
rect 15344 18640 15350 18692
rect 16114 18640 16120 18692
rect 16172 18640 16178 18692
rect 21174 18680 21180 18692
rect 19444 18652 21180 18680
rect 19444 18612 19472 18652
rect 21174 18640 21180 18652
rect 21232 18640 21238 18692
rect 10888 18584 19472 18612
rect 19521 18615 19579 18621
rect 19521 18581 19533 18615
rect 19567 18612 19579 18615
rect 19978 18612 19984 18624
rect 19567 18584 19984 18612
rect 19567 18581 19579 18584
rect 19521 18575 19579 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 45830 18572 45836 18624
rect 45888 18612 45894 18624
rect 57238 18612 57244 18624
rect 45888 18584 57244 18612
rect 45888 18572 45894 18584
rect 57238 18572 57244 18584
rect 57296 18572 57302 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 2317 18411 2375 18417
rect 2317 18408 2329 18411
rect 2004 18380 2329 18408
rect 2004 18368 2010 18380
rect 2317 18377 2329 18380
rect 2363 18377 2375 18411
rect 2682 18408 2688 18420
rect 2643 18380 2688 18408
rect 2317 18371 2375 18377
rect 2332 18340 2360 18371
rect 2682 18368 2688 18380
rect 2740 18368 2746 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 7469 18411 7527 18417
rect 7469 18408 7481 18411
rect 5960 18380 7481 18408
rect 5960 18368 5966 18380
rect 7469 18377 7481 18380
rect 7515 18377 7527 18411
rect 12161 18411 12219 18417
rect 7469 18371 7527 18377
rect 7668 18380 8616 18408
rect 3145 18343 3203 18349
rect 3145 18340 3157 18343
rect 2332 18312 3157 18340
rect 3145 18309 3157 18312
rect 3191 18309 3203 18343
rect 7668 18340 7696 18380
rect 8588 18340 8616 18380
rect 12161 18377 12173 18411
rect 12207 18408 12219 18411
rect 12250 18408 12256 18420
rect 12207 18380 12256 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 17126 18368 17132 18420
rect 17184 18408 17190 18420
rect 18969 18411 19027 18417
rect 18969 18408 18981 18411
rect 17184 18380 18981 18408
rect 17184 18368 17190 18380
rect 18969 18377 18981 18380
rect 19015 18408 19027 18411
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 19015 18380 19809 18408
rect 19015 18377 19027 18380
rect 18969 18371 19027 18377
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 20254 18408 20260 18420
rect 20215 18380 20260 18408
rect 19797 18371 19855 18377
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 9030 18340 9036 18352
rect 5290 18312 7696 18340
rect 8510 18312 9036 18340
rect 3145 18303 3203 18309
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 14737 18343 14795 18349
rect 14737 18309 14749 18343
rect 14783 18340 14795 18343
rect 15102 18340 15108 18352
rect 14783 18312 15108 18340
rect 14783 18309 14795 18312
rect 14737 18303 14795 18309
rect 15102 18300 15108 18312
rect 15160 18300 15166 18352
rect 15286 18300 15292 18352
rect 15344 18340 15350 18352
rect 21450 18340 21456 18352
rect 15344 18312 21456 18340
rect 15344 18300 15350 18312
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 2958 18272 2964 18284
rect 2148 18244 2964 18272
rect 2148 18213 2176 18244
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 11054 18232 11060 18284
rect 11112 18272 11118 18284
rect 12345 18275 12403 18281
rect 12345 18272 12357 18275
rect 11112 18244 12357 18272
rect 11112 18232 11118 18244
rect 12345 18241 12357 18244
rect 12391 18241 12403 18275
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 12345 18235 12403 18241
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18272 19947 18275
rect 20162 18272 20168 18284
rect 19935 18244 20168 18272
rect 19935 18241 19947 18244
rect 19889 18235 19947 18241
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 57517 18275 57575 18281
rect 57517 18241 57529 18275
rect 57563 18272 57575 18275
rect 58342 18272 58348 18284
rect 57563 18244 58348 18272
rect 57563 18241 57575 18244
rect 57517 18235 57575 18241
rect 58342 18232 58348 18244
rect 58400 18232 58406 18284
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18173 2191 18207
rect 2133 18167 2191 18173
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2280 18176 2373 18204
rect 2280 18164 2286 18176
rect 2498 18164 2504 18216
rect 2556 18204 2562 18216
rect 5721 18207 5779 18213
rect 5721 18204 5733 18207
rect 2556 18176 5733 18204
rect 2556 18164 2562 18176
rect 5721 18173 5733 18176
rect 5767 18173 5779 18207
rect 5721 18167 5779 18173
rect 5997 18207 6055 18213
rect 5997 18173 6009 18207
rect 6043 18204 6055 18207
rect 6178 18204 6184 18216
rect 6043 18176 6184 18204
rect 6043 18173 6055 18176
rect 5997 18167 6055 18173
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 6822 18164 6828 18216
rect 6880 18204 6886 18216
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 6880 18176 8953 18204
rect 6880 18164 6886 18176
rect 8941 18173 8953 18176
rect 8987 18173 8999 18207
rect 9214 18204 9220 18216
rect 9175 18176 9220 18204
rect 8941 18167 8999 18173
rect 9214 18164 9220 18176
rect 9272 18164 9278 18216
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 19751 18176 20484 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 2240 18136 2268 18164
rect 4249 18139 4307 18145
rect 4249 18136 4261 18139
rect 2240 18108 4261 18136
rect 4249 18105 4261 18108
rect 4295 18105 4307 18139
rect 4249 18099 4307 18105
rect 20456 18080 20484 18176
rect 11054 18068 11060 18080
rect 11015 18040 11060 18068
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 20438 18028 20444 18080
rect 20496 18068 20502 18080
rect 20717 18071 20775 18077
rect 20717 18068 20729 18071
rect 20496 18040 20729 18068
rect 20496 18028 20502 18040
rect 20717 18037 20729 18040
rect 20763 18037 20775 18071
rect 20717 18031 20775 18037
rect 57422 18028 57428 18080
rect 57480 18068 57486 18080
rect 58161 18071 58219 18077
rect 58161 18068 58173 18071
rect 57480 18040 58173 18068
rect 57480 18028 57486 18040
rect 58161 18037 58173 18040
rect 58207 18037 58219 18071
rect 58161 18031 58219 18037
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 11885 17867 11943 17873
rect 11885 17833 11897 17867
rect 11931 17864 11943 17867
rect 15378 17864 15384 17876
rect 11931 17836 15384 17864
rect 11931 17833 11943 17836
rect 11885 17827 11943 17833
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 17129 17867 17187 17873
rect 17129 17833 17141 17867
rect 17175 17864 17187 17867
rect 18230 17864 18236 17876
rect 17175 17836 18236 17864
rect 17175 17833 17187 17836
rect 17129 17827 17187 17833
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 21450 17864 21456 17876
rect 21411 17836 21456 17864
rect 21450 17824 21456 17836
rect 21508 17824 21514 17876
rect 2958 17796 2964 17808
rect 2056 17768 2964 17796
rect 2056 17737 2084 17768
rect 2958 17756 2964 17768
rect 3016 17756 3022 17808
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 2130 17688 2136 17740
rect 2188 17728 2194 17740
rect 2225 17731 2283 17737
rect 2225 17728 2237 17731
rect 2188 17700 2237 17728
rect 2188 17688 2194 17700
rect 2225 17697 2237 17700
rect 2271 17728 2283 17731
rect 2406 17728 2412 17740
rect 2271 17700 2412 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 2406 17688 2412 17700
rect 2464 17688 2470 17740
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17728 13415 17731
rect 13998 17728 14004 17740
rect 13403 17700 14004 17728
rect 13403 17697 13415 17700
rect 13357 17691 13415 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 16022 17728 16028 17740
rect 15703 17700 16028 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17697 20315 17731
rect 20257 17691 20315 17697
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 3326 17660 3332 17672
rect 2363 17632 3332 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 1762 17552 1768 17604
rect 1820 17592 1826 17604
rect 2130 17592 2136 17604
rect 1820 17564 2136 17592
rect 1820 17552 1826 17564
rect 2130 17552 2136 17564
rect 2188 17552 2194 17604
rect 2682 17524 2688 17536
rect 2643 17496 2688 17524
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 3252 17533 3280 17632
rect 3326 17620 3332 17632
rect 3384 17620 3390 17672
rect 13633 17663 13691 17669
rect 13633 17629 13645 17663
rect 13679 17660 13691 17663
rect 15194 17660 15200 17672
rect 13679 17632 15200 17660
rect 13679 17629 13691 17632
rect 13633 17623 13691 17629
rect 15194 17620 15200 17632
rect 15252 17660 15258 17672
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 15252 17632 15393 17660
rect 15252 17620 15258 17632
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 15381 17623 15439 17629
rect 11698 17552 11704 17604
rect 11756 17592 11762 17604
rect 11756 17564 12190 17592
rect 11756 17552 11762 17564
rect 16666 17552 16672 17604
rect 16724 17552 16730 17604
rect 19981 17595 20039 17601
rect 19981 17561 19993 17595
rect 20027 17592 20039 17595
rect 20162 17592 20168 17604
rect 20027 17564 20168 17592
rect 20027 17561 20039 17564
rect 19981 17555 20039 17561
rect 20162 17552 20168 17564
rect 20220 17552 20226 17604
rect 3237 17527 3295 17533
rect 3237 17493 3249 17527
rect 3283 17524 3295 17527
rect 3970 17524 3976 17536
rect 3283 17496 3976 17524
rect 3283 17493 3295 17496
rect 3237 17487 3295 17493
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 19426 17484 19432 17536
rect 19484 17524 19490 17536
rect 19613 17527 19671 17533
rect 19613 17524 19625 17527
rect 19484 17496 19625 17524
rect 19484 17484 19490 17496
rect 19613 17493 19625 17496
rect 19659 17493 19671 17527
rect 20070 17524 20076 17536
rect 20031 17496 20076 17524
rect 19613 17487 19671 17493
rect 20070 17484 20076 17496
rect 20128 17484 20134 17536
rect 20272 17524 20300 17691
rect 21634 17660 21640 17672
rect 21595 17632 21640 17660
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 57701 17663 57759 17669
rect 57701 17629 57713 17663
rect 57747 17660 57759 17663
rect 58342 17660 58348 17672
rect 57747 17632 58348 17660
rect 57747 17629 57759 17632
rect 57701 17623 57759 17629
rect 58342 17620 58348 17632
rect 58400 17620 58406 17672
rect 20622 17524 20628 17536
rect 20272 17496 20628 17524
rect 20622 17484 20628 17496
rect 20680 17524 20686 17536
rect 20901 17527 20959 17533
rect 20901 17524 20913 17527
rect 20680 17496 20913 17524
rect 20680 17484 20686 17496
rect 20901 17493 20913 17496
rect 20947 17524 20959 17527
rect 23474 17524 23480 17536
rect 20947 17496 23480 17524
rect 20947 17493 20959 17496
rect 20901 17487 20959 17493
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 58161 17527 58219 17533
rect 58161 17493 58173 17527
rect 58207 17524 58219 17527
rect 58710 17524 58716 17536
rect 58207 17496 58716 17524
rect 58207 17493 58219 17496
rect 58161 17487 58219 17493
rect 58710 17484 58716 17496
rect 58768 17484 58774 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 1670 17320 1676 17332
rect 1631 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 8294 17320 8300 17332
rect 8255 17292 8300 17320
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 19521 17323 19579 17329
rect 19521 17320 19533 17323
rect 19392 17292 19533 17320
rect 19392 17280 19398 17292
rect 19521 17289 19533 17292
rect 19567 17320 19579 17323
rect 20070 17320 20076 17332
rect 19567 17292 20076 17320
rect 19567 17289 19579 17292
rect 19521 17283 19579 17289
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 4890 17212 4896 17264
rect 4948 17252 4954 17264
rect 16298 17252 16304 17264
rect 4948 17224 16304 17252
rect 4948 17212 4954 17224
rect 16298 17212 16304 17224
rect 16356 17212 16362 17264
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 2222 17184 2228 17196
rect 1903 17156 2228 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 2682 17184 2688 17196
rect 2363 17156 2688 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2682 17144 2688 17156
rect 2740 17144 2746 17196
rect 9582 17184 9588 17196
rect 9543 17156 9588 17184
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 2498 16980 2504 16992
rect 2459 16952 2504 16980
rect 2498 16940 2504 16952
rect 2556 16940 2562 16992
rect 2958 16980 2964 16992
rect 2919 16952 2964 16980
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 21174 16776 21180 16788
rect 21135 16748 21180 16776
rect 21174 16736 21180 16748
rect 21232 16736 21238 16788
rect 21634 16736 21640 16788
rect 21692 16776 21698 16788
rect 21729 16779 21787 16785
rect 21729 16776 21741 16779
rect 21692 16748 21741 16776
rect 21692 16736 21698 16748
rect 21729 16745 21741 16748
rect 21775 16745 21787 16779
rect 21729 16739 21787 16745
rect 20548 16680 22324 16708
rect 2498 16600 2504 16652
rect 2556 16640 2562 16652
rect 5905 16643 5963 16649
rect 5905 16640 5917 16643
rect 2556 16612 5917 16640
rect 2556 16600 2562 16612
rect 5905 16609 5917 16612
rect 5951 16609 5963 16643
rect 9122 16640 9128 16652
rect 9083 16612 9128 16640
rect 5905 16603 5963 16609
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 9398 16640 9404 16652
rect 9359 16612 9404 16640
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 1578 16532 1584 16584
rect 1636 16572 1642 16584
rect 1857 16575 1915 16581
rect 1857 16572 1869 16575
rect 1636 16544 1869 16572
rect 1636 16532 1642 16544
rect 1857 16541 1869 16544
rect 1903 16572 1915 16575
rect 2317 16575 2375 16581
rect 2317 16572 2329 16575
rect 1903 16544 2329 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 2317 16541 2329 16544
rect 2363 16541 2375 16575
rect 2317 16535 2375 16541
rect 6178 16532 6184 16584
rect 6236 16572 6242 16584
rect 9140 16572 9168 16600
rect 6236 16544 9168 16572
rect 6236 16532 6242 16544
rect 16942 16532 16948 16584
rect 17000 16572 17006 16584
rect 19334 16572 19340 16584
rect 17000 16544 19340 16572
rect 17000 16532 17006 16544
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 19613 16575 19671 16581
rect 19613 16572 19625 16575
rect 19484 16544 19625 16572
rect 19484 16532 19490 16544
rect 19613 16541 19625 16544
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16572 20315 16575
rect 20346 16572 20352 16584
rect 20303 16544 20352 16572
rect 20303 16541 20315 16544
rect 20257 16535 20315 16541
rect 20346 16532 20352 16544
rect 20404 16532 20410 16584
rect 20438 16532 20444 16584
rect 20496 16572 20502 16584
rect 20548 16581 20576 16680
rect 21174 16600 21180 16652
rect 21232 16640 21238 16652
rect 22296 16649 22324 16680
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 21232 16612 22201 16640
rect 21232 16600 21238 16612
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 22189 16603 22247 16609
rect 22281 16643 22339 16649
rect 22281 16609 22293 16643
rect 22327 16609 22339 16643
rect 22281 16603 22339 16609
rect 20533 16575 20591 16581
rect 20533 16572 20545 16575
rect 20496 16544 20545 16572
rect 20496 16532 20502 16544
rect 20533 16541 20545 16544
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 57701 16575 57759 16581
rect 57701 16541 57713 16575
rect 57747 16572 57759 16575
rect 58342 16572 58348 16584
rect 57747 16544 58348 16572
rect 57747 16541 57759 16544
rect 57701 16535 57759 16541
rect 58342 16532 58348 16544
rect 58400 16532 58406 16584
rect 5350 16464 5356 16516
rect 5408 16464 5414 16516
rect 9030 16464 9036 16516
rect 9088 16504 9094 16516
rect 9088 16476 9890 16504
rect 9088 16464 9094 16476
rect 1670 16436 1676 16448
rect 1631 16408 1676 16436
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 2406 16396 2412 16448
rect 2464 16436 2470 16448
rect 4433 16439 4491 16445
rect 4433 16436 4445 16439
rect 2464 16408 4445 16436
rect 2464 16396 2470 16408
rect 4433 16405 4445 16408
rect 4479 16405 4491 16439
rect 4433 16399 4491 16405
rect 10686 16396 10692 16448
rect 10744 16436 10750 16448
rect 10873 16439 10931 16445
rect 10873 16436 10885 16439
rect 10744 16408 10885 16436
rect 10744 16396 10750 16408
rect 10873 16405 10885 16408
rect 10919 16405 10931 16439
rect 19426 16436 19432 16448
rect 19387 16408 19432 16436
rect 10873 16399 10931 16405
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 22097 16439 22155 16445
rect 22097 16405 22109 16439
rect 22143 16436 22155 16439
rect 22278 16436 22284 16448
rect 22143 16408 22284 16436
rect 22143 16405 22155 16408
rect 22097 16399 22155 16405
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 56778 16396 56784 16448
rect 56836 16436 56842 16448
rect 58161 16439 58219 16445
rect 58161 16436 58173 16439
rect 56836 16408 58173 16436
rect 56836 16396 56842 16408
rect 58161 16405 58173 16408
rect 58207 16405 58219 16439
rect 58161 16399 58219 16405
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 9122 16232 9128 16244
rect 8343 16204 9128 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 3326 16096 3332 16108
rect 1903 16068 3332 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 9582 16096 9588 16108
rect 9495 16068 9588 16096
rect 9582 16056 9588 16068
rect 9640 16096 9646 16108
rect 12986 16096 12992 16108
rect 9640 16068 12992 16096
rect 9640 16056 9646 16068
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 58342 16096 58348 16108
rect 58303 16068 58348 16096
rect 58342 16056 58348 16068
rect 58400 16056 58406 16108
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 2958 15892 2964 15904
rect 2915 15864 2964 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 3326 15892 3332 15904
rect 3287 15864 3332 15892
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 12526 15852 12532 15904
rect 12584 15892 12590 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 12584 15864 14289 15892
rect 12584 15852 12590 15864
rect 14277 15861 14289 15864
rect 14323 15892 14335 15895
rect 15194 15892 15200 15904
rect 14323 15864 15200 15892
rect 14323 15861 14335 15864
rect 14277 15855 14335 15861
rect 15194 15852 15200 15864
rect 15252 15892 15258 15904
rect 15378 15892 15384 15904
rect 15252 15864 15384 15892
rect 15252 15852 15258 15864
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 57790 15852 57796 15904
rect 57848 15892 57854 15904
rect 58161 15895 58219 15901
rect 58161 15892 58173 15895
rect 57848 15864 58173 15892
rect 57848 15852 57854 15864
rect 58161 15861 58173 15864
rect 58207 15861 58219 15895
rect 58161 15855 58219 15861
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2038 15648 2044 15700
rect 2096 15648 2102 15700
rect 3234 15688 3240 15700
rect 3195 15660 3240 15688
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 10410 15648 10416 15700
rect 10468 15688 10474 15700
rect 10505 15691 10563 15697
rect 10505 15688 10517 15691
rect 10468 15660 10517 15688
rect 10468 15648 10474 15660
rect 10505 15657 10517 15660
rect 10551 15657 10563 15691
rect 10505 15651 10563 15657
rect 16942 15648 16948 15700
rect 17000 15688 17006 15700
rect 17129 15691 17187 15697
rect 17129 15688 17141 15691
rect 17000 15660 17141 15688
rect 17000 15648 17006 15660
rect 17129 15657 17141 15660
rect 17175 15657 17187 15691
rect 58342 15688 58348 15700
rect 58303 15660 58348 15688
rect 17129 15651 17187 15657
rect 58342 15648 58348 15660
rect 58400 15648 58406 15700
rect 2056 15620 2084 15648
rect 4341 15623 4399 15629
rect 4341 15620 4353 15623
rect 2056 15592 4353 15620
rect 2240 15561 2268 15592
rect 4341 15589 4353 15592
rect 4387 15589 4399 15623
rect 4341 15583 4399 15589
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15521 2191 15555
rect 2133 15515 2191 15521
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15521 2283 15555
rect 2225 15515 2283 15521
rect 2148 15484 2176 15515
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 5813 15555 5871 15561
rect 5813 15552 5825 15555
rect 4304 15524 5825 15552
rect 4304 15512 4310 15524
rect 5813 15521 5825 15524
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 6089 15555 6147 15561
rect 6089 15521 6101 15555
rect 6135 15552 6147 15555
rect 6178 15552 6184 15564
rect 6135 15524 6184 15552
rect 6135 15521 6147 15524
rect 6089 15515 6147 15521
rect 6178 15512 6184 15524
rect 6236 15552 6242 15564
rect 6822 15552 6828 15564
rect 6236 15524 6828 15552
rect 6236 15512 6242 15524
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 15378 15552 15384 15564
rect 15339 15524 15384 15552
rect 15378 15512 15384 15524
rect 15436 15512 15442 15564
rect 15657 15555 15715 15561
rect 15657 15521 15669 15555
rect 15703 15552 15715 15555
rect 19426 15552 19432 15564
rect 15703 15524 19432 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 2958 15484 2964 15496
rect 2148 15456 2964 15484
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12526 15484 12532 15496
rect 12299 15456 12532 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 2317 15419 2375 15425
rect 2317 15385 2329 15419
rect 2363 15416 2375 15419
rect 3234 15416 3240 15428
rect 2363 15388 3240 15416
rect 2363 15385 2375 15388
rect 2317 15379 2375 15385
rect 3234 15376 3240 15388
rect 3292 15376 3298 15428
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 9030 15416 9036 15428
rect 5408 15388 9036 15416
rect 5408 15376 5414 15388
rect 9030 15376 9036 15388
rect 9088 15376 9094 15428
rect 11698 15416 11704 15428
rect 11546 15388 11704 15416
rect 11698 15376 11704 15388
rect 11756 15376 11762 15428
rect 11977 15419 12035 15425
rect 11977 15385 11989 15419
rect 12023 15416 12035 15419
rect 12066 15416 12072 15428
rect 12023 15388 12072 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 16666 15376 16672 15428
rect 16724 15376 16730 15428
rect 2682 15348 2688 15360
rect 2643 15320 2688 15348
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 4246 15144 4252 15156
rect 2547 15116 4252 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 5537 15147 5595 15153
rect 5537 15144 5549 15147
rect 5408 15116 5549 15144
rect 5408 15104 5414 15116
rect 5537 15113 5549 15116
rect 5583 15113 5595 15147
rect 6546 15144 6552 15156
rect 5537 15107 5595 15113
rect 5828 15116 6552 15144
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 5828 15085 5856 15116
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 7742 15104 7748 15156
rect 7800 15144 7806 15156
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 7800 15116 8953 15144
rect 7800 15104 7806 15116
rect 8941 15113 8953 15116
rect 8987 15113 8999 15147
rect 8941 15107 8999 15113
rect 5813 15079 5871 15085
rect 5813 15076 5825 15079
rect 5776 15048 5825 15076
rect 5776 15036 5782 15048
rect 5813 15045 5825 15048
rect 5859 15045 5871 15079
rect 5813 15039 5871 15045
rect 6454 15036 6460 15088
rect 6512 15076 6518 15088
rect 7469 15079 7527 15085
rect 7469 15076 7481 15079
rect 6512 15048 7481 15076
rect 6512 15036 6518 15048
rect 7469 15045 7481 15048
rect 7515 15045 7527 15079
rect 9030 15076 9036 15088
rect 8694 15048 9036 15076
rect 7469 15039 7527 15045
rect 9030 15036 9036 15048
rect 9088 15036 9094 15088
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 14977 1915 15011
rect 1857 14971 1915 14977
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 2682 15008 2688 15020
rect 2363 14980 2688 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 1872 14940 1900 14971
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7193 15011 7251 15017
rect 7193 15008 7205 15011
rect 6972 14980 7205 15008
rect 6972 14968 6978 14980
rect 7193 14977 7205 14980
rect 7239 14977 7251 15011
rect 20162 15008 20168 15020
rect 20123 14980 20168 15008
rect 7193 14971 7251 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 57517 15011 57575 15017
rect 57517 14977 57529 15011
rect 57563 15008 57575 15011
rect 58342 15008 58348 15020
rect 57563 14980 58348 15008
rect 57563 14977 57575 14980
rect 57517 14971 57575 14977
rect 58342 14968 58348 14980
rect 58400 14968 58406 15020
rect 3053 14943 3111 14949
rect 3053 14940 3065 14943
rect 1872 14912 3065 14940
rect 3053 14909 3065 14912
rect 3099 14940 3111 14943
rect 8938 14940 8944 14952
rect 3099 14912 8944 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 8938 14900 8944 14912
rect 8996 14900 9002 14952
rect 20257 14943 20315 14949
rect 20257 14940 20269 14943
rect 19352 14912 20269 14940
rect 1670 14872 1676 14884
rect 1631 14844 1676 14872
rect 1670 14832 1676 14844
rect 1728 14832 1734 14884
rect 19352 14816 19380 14912
rect 20257 14909 20269 14912
rect 20303 14909 20315 14943
rect 20438 14940 20444 14952
rect 20399 14912 20444 14940
rect 20257 14903 20315 14909
rect 20438 14900 20444 14912
rect 20496 14900 20502 14952
rect 6546 14764 6552 14816
rect 6604 14804 6610 14816
rect 11054 14804 11060 14816
rect 6604 14776 11060 14804
rect 6604 14764 6610 14776
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 19334 14804 19340 14816
rect 19295 14776 19340 14804
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19797 14807 19855 14813
rect 19797 14773 19809 14807
rect 19843 14804 19855 14807
rect 20070 14804 20076 14816
rect 19843 14776 20076 14804
rect 19843 14773 19855 14776
rect 19797 14767 19855 14773
rect 20070 14764 20076 14776
rect 20128 14764 20134 14816
rect 57330 14764 57336 14816
rect 57388 14804 57394 14816
rect 58161 14807 58219 14813
rect 58161 14804 58173 14807
rect 57388 14776 58173 14804
rect 57388 14764 57394 14776
rect 58161 14773 58173 14776
rect 58207 14773 58219 14807
rect 58161 14767 58219 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 13262 14600 13268 14612
rect 10520 14572 13268 14600
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14464 2191 14467
rect 2958 14464 2964 14476
rect 2179 14436 2964 14464
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 10520 14473 10548 14572
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 22094 14600 22100 14612
rect 13872 14572 22100 14600
rect 13872 14560 13878 14572
rect 22094 14560 22100 14572
rect 22152 14560 22158 14612
rect 19426 14492 19432 14544
rect 19484 14532 19490 14544
rect 22281 14535 22339 14541
rect 22281 14532 22293 14535
rect 19484 14504 22293 14532
rect 19484 14492 19490 14504
rect 22281 14501 22293 14504
rect 22327 14501 22339 14535
rect 22281 14495 22339 14501
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14433 10563 14467
rect 10505 14427 10563 14433
rect 12158 14424 12164 14476
rect 12216 14464 12222 14476
rect 12253 14467 12311 14473
rect 12253 14464 12265 14467
rect 12216 14436 12265 14464
rect 12216 14424 12222 14436
rect 12253 14433 12265 14436
rect 12299 14433 12311 14467
rect 12526 14464 12532 14476
rect 12487 14436 12532 14464
rect 12253 14427 12311 14433
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 15749 14467 15807 14473
rect 15749 14464 15761 14467
rect 15436 14436 15761 14464
rect 15436 14424 15442 14436
rect 15749 14433 15761 14436
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 17773 14467 17831 14473
rect 16071 14436 17540 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 17512 14396 17540 14436
rect 17773 14433 17785 14467
rect 17819 14464 17831 14467
rect 18782 14464 18788 14476
rect 17819 14436 18788 14464
rect 17819 14433 17831 14436
rect 17773 14427 17831 14433
rect 18782 14424 18788 14436
rect 18840 14424 18846 14476
rect 20346 14424 20352 14476
rect 20404 14464 20410 14476
rect 20530 14464 20536 14476
rect 20404 14436 20536 14464
rect 20404 14424 20410 14436
rect 20530 14424 20536 14436
rect 20588 14464 20594 14476
rect 21085 14467 21143 14473
rect 21085 14464 21097 14467
rect 20588 14436 21097 14464
rect 20588 14424 20594 14436
rect 21085 14433 21097 14436
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 19978 14396 19984 14408
rect 17512 14368 19984 14396
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 22186 14356 22192 14408
rect 22244 14396 22250 14408
rect 22465 14399 22523 14405
rect 22465 14396 22477 14399
rect 22244 14368 22477 14396
rect 22244 14356 22250 14368
rect 22465 14365 22477 14368
rect 22511 14365 22523 14399
rect 22465 14359 22523 14365
rect 57701 14399 57759 14405
rect 57701 14365 57713 14399
rect 57747 14396 57759 14399
rect 58342 14396 58348 14408
rect 57747 14368 58348 14396
rect 57747 14365 57759 14368
rect 57701 14359 57759 14365
rect 58342 14356 58348 14368
rect 58400 14356 58406 14408
rect 1762 14288 1768 14340
rect 1820 14328 1826 14340
rect 2130 14328 2136 14340
rect 1820 14300 2136 14328
rect 1820 14288 1826 14300
rect 2130 14288 2136 14300
rect 2188 14328 2194 14340
rect 2317 14331 2375 14337
rect 2317 14328 2329 14331
rect 2188 14300 2329 14328
rect 2188 14288 2194 14300
rect 2317 14297 2329 14300
rect 2363 14328 2375 14331
rect 3145 14331 3203 14337
rect 3145 14328 3157 14331
rect 2363 14300 3157 14328
rect 2363 14297 2375 14300
rect 2317 14291 2375 14297
rect 3145 14297 3157 14300
rect 3191 14297 3203 14331
rect 3145 14291 3203 14297
rect 11698 14288 11704 14340
rect 11756 14288 11762 14340
rect 16666 14288 16672 14340
rect 16724 14288 16730 14340
rect 20349 14331 20407 14337
rect 20349 14328 20361 14331
rect 18800 14300 20361 14328
rect 18800 14272 18828 14300
rect 20349 14297 20361 14300
rect 20395 14297 20407 14331
rect 20349 14291 20407 14297
rect 2222 14260 2228 14272
rect 2183 14232 2228 14260
rect 2222 14220 2228 14232
rect 2280 14220 2286 14272
rect 2682 14260 2688 14272
rect 2643 14232 2688 14260
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 18782 14260 18788 14272
rect 18743 14232 18788 14260
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 19889 14263 19947 14269
rect 19889 14229 19901 14263
rect 19935 14260 19947 14263
rect 19978 14260 19984 14272
rect 19935 14232 19984 14260
rect 19935 14229 19947 14232
rect 19889 14223 19947 14229
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 20257 14263 20315 14269
rect 20257 14229 20269 14263
rect 20303 14260 20315 14263
rect 20530 14260 20536 14272
rect 20303 14232 20536 14260
rect 20303 14229 20315 14232
rect 20257 14223 20315 14229
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 57974 14220 57980 14272
rect 58032 14260 58038 14272
rect 58161 14263 58219 14269
rect 58161 14260 58173 14263
rect 58032 14232 58173 14260
rect 58032 14220 58038 14232
rect 58161 14229 58173 14232
rect 58207 14229 58219 14263
rect 58161 14223 58219 14229
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 1670 14056 1676 14068
rect 1631 14028 1676 14056
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 3878 14056 3884 14068
rect 2547 14028 3884 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 11054 14056 11060 14068
rect 11015 14028 11060 14056
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 13814 14056 13820 14068
rect 13775 14028 13820 14056
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 13924 14028 16574 14056
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13889 1915 13923
rect 1857 13883 1915 13889
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13920 2375 13923
rect 2682 13920 2688 13932
rect 2363 13892 2688 13920
rect 2363 13889 2375 13892
rect 2317 13883 2375 13889
rect 1872 13852 1900 13883
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 11072 13920 11100 14016
rect 11698 13988 11704 14000
rect 11659 13960 11704 13988
rect 11698 13948 11704 13960
rect 11756 13988 11762 14000
rect 13924 13988 13952 14028
rect 14936 13988 14964 14028
rect 11756 13960 13952 13988
rect 14858 13960 14964 13988
rect 11756 13948 11762 13960
rect 15378 13948 15384 14000
rect 15436 13988 15442 14000
rect 16546 13988 16574 14028
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 19705 14059 19763 14065
rect 19705 14056 19717 14059
rect 18104 14028 19717 14056
rect 18104 14016 18110 14028
rect 19705 14025 19717 14028
rect 19751 14025 19763 14059
rect 22186 14056 22192 14068
rect 22147 14028 22192 14056
rect 19705 14019 19763 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 16666 13988 16672 14000
rect 15436 13960 15608 13988
rect 16546 13960 16672 13988
rect 15436 13948 15442 13960
rect 12066 13920 12072 13932
rect 11072 13892 12072 13920
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 15580 13929 15608 13960
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 56686 13948 56692 14000
rect 56744 13988 56750 14000
rect 56781 13991 56839 13997
rect 56781 13988 56793 13991
rect 56744 13960 56793 13988
rect 56744 13948 56750 13960
rect 56781 13957 56793 13960
rect 56827 13988 56839 13991
rect 56870 13988 56876 14000
rect 56827 13960 56876 13988
rect 56827 13957 56839 13960
rect 56781 13951 56839 13957
rect 56870 13948 56876 13960
rect 56928 13988 56934 14000
rect 57698 13988 57704 14000
rect 56928 13960 57704 13988
rect 56928 13948 56934 13960
rect 57698 13948 57704 13960
rect 57756 13988 57762 14000
rect 58253 13991 58311 13997
rect 58253 13988 58265 13991
rect 57756 13960 58265 13988
rect 57756 13948 57762 13960
rect 58253 13957 58265 13960
rect 58299 13957 58311 13991
rect 58253 13951 58311 13957
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20070 13920 20076 13932
rect 19935 13892 20076 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20530 13880 20536 13932
rect 20588 13920 20594 13932
rect 22278 13920 22284 13932
rect 20588 13892 22284 13920
rect 20588 13880 20594 13892
rect 22278 13880 22284 13892
rect 22336 13920 22342 13932
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 22336 13892 22569 13920
rect 22336 13880 22342 13892
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 56505 13923 56563 13929
rect 56505 13920 56517 13923
rect 22557 13883 22615 13889
rect 56060 13892 56517 13920
rect 56060 13864 56088 13892
rect 56505 13889 56517 13892
rect 56551 13889 56563 13923
rect 56505 13883 56563 13889
rect 2406 13852 2412 13864
rect 1872 13824 2412 13852
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 2958 13852 2964 13864
rect 2919 13824 2964 13852
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 11698 13852 11704 13864
rect 6328 13824 11704 13852
rect 6328 13812 6334 13824
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15335 13824 15516 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15488 13784 15516 13824
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 22649 13855 22707 13861
rect 22649 13852 22661 13855
rect 22152 13824 22661 13852
rect 22152 13812 22158 13824
rect 22649 13821 22661 13824
rect 22695 13821 22707 13855
rect 22649 13815 22707 13821
rect 22833 13855 22891 13861
rect 22833 13821 22845 13855
rect 22879 13821 22891 13855
rect 56042 13852 56048 13864
rect 56003 13824 56048 13852
rect 22833 13815 22891 13821
rect 19426 13784 19432 13796
rect 15488 13756 19432 13784
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 22848 13784 22876 13815
rect 56042 13812 56048 13824
rect 56100 13812 56106 13864
rect 23474 13784 23480 13796
rect 22848 13756 23480 13784
rect 23474 13744 23480 13756
rect 23532 13744 23538 13796
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 22554 13716 22560 13728
rect 11756 13688 22560 13716
rect 11756 13676 11762 13688
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 3602 13472 3608 13524
rect 3660 13512 3666 13524
rect 16206 13512 16212 13524
rect 3660 13484 13676 13512
rect 16167 13484 16212 13512
rect 3660 13472 3666 13484
rect 2222 13404 2228 13456
rect 2280 13444 2286 13456
rect 4341 13447 4399 13453
rect 4341 13444 4353 13447
rect 2280 13416 4353 13444
rect 2280 13404 2286 13416
rect 4341 13413 4353 13416
rect 4387 13413 4399 13447
rect 13648 13444 13676 13484
rect 16206 13472 16212 13484
rect 16264 13512 16270 13524
rect 19334 13512 19340 13524
rect 16264 13484 19340 13512
rect 16264 13472 16270 13484
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 22094 13512 22100 13524
rect 22055 13484 22100 13512
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 22554 13512 22560 13524
rect 22515 13484 22560 13512
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 16666 13444 16672 13456
rect 13648 13416 16672 13444
rect 4341 13407 4399 13413
rect 16666 13404 16672 13416
rect 16724 13404 16730 13456
rect 58066 13444 58072 13456
rect 57624 13416 58072 13444
rect 3878 13336 3884 13388
rect 3936 13376 3942 13388
rect 5813 13379 5871 13385
rect 5813 13376 5825 13379
rect 3936 13348 5825 13376
rect 3936 13336 3942 13348
rect 5813 13345 5825 13348
rect 5859 13345 5871 13379
rect 11698 13376 11704 13388
rect 11659 13348 11704 13376
rect 5813 13339 5871 13345
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13376 17739 13379
rect 18046 13376 18052 13388
rect 17727 13348 18052 13376
rect 17727 13345 17739 13348
rect 17681 13339 17739 13345
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 57146 13376 57152 13388
rect 57107 13348 57152 13376
rect 57146 13336 57152 13348
rect 57204 13336 57210 13388
rect 57330 13385 57336 13388
rect 57308 13379 57336 13385
rect 57308 13345 57320 13379
rect 57308 13339 57336 13345
rect 57330 13336 57336 13339
rect 57388 13336 57394 13388
rect 57425 13379 57483 13385
rect 57425 13345 57437 13379
rect 57471 13376 57483 13379
rect 57624 13376 57652 13416
rect 58066 13404 58072 13416
rect 58124 13404 58130 13456
rect 57471 13348 57652 13376
rect 57471 13345 57483 13348
rect 57425 13339 57483 13345
rect 57698 13336 57704 13388
rect 57756 13376 57762 13388
rect 58161 13379 58219 13385
rect 57756 13348 57801 13376
rect 57756 13336 57762 13348
rect 58161 13345 58173 13379
rect 58207 13376 58219 13379
rect 58526 13376 58532 13388
rect 58207 13348 58532 13376
rect 58207 13345 58219 13348
rect 58161 13339 58219 13345
rect 58526 13336 58532 13348
rect 58584 13336 58590 13388
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13308 1915 13311
rect 2038 13308 2044 13320
rect 1903 13280 2044 13308
rect 1903 13277 1915 13280
rect 1857 13271 1915 13277
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 6914 13308 6920 13320
rect 6135 13280 6920 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 6914 13268 6920 13280
rect 6972 13268 6978 13320
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13308 13783 13311
rect 13814 13308 13820 13320
rect 13771 13280 13820 13308
rect 13771 13277 13783 13280
rect 13725 13271 13783 13277
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13277 18015 13311
rect 17957 13271 18015 13277
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 19978 13308 19984 13320
rect 19935 13280 19984 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 2372 13212 2544 13240
rect 2372 13200 2378 13212
rect 1670 13172 1676 13184
rect 1631 13144 1676 13172
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 2406 13172 2412 13184
rect 2367 13144 2412 13172
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 2516 13172 2544 13212
rect 5166 13200 5172 13252
rect 5224 13200 5230 13252
rect 12158 13200 12164 13252
rect 12216 13240 12222 13252
rect 13446 13240 13452 13252
rect 12216 13212 12282 13240
rect 13407 13212 13452 13240
rect 12216 13200 12222 13212
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 16666 13200 16672 13252
rect 16724 13200 16730 13252
rect 17770 13200 17776 13252
rect 17828 13240 17834 13252
rect 17972 13240 18000 13271
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 58250 13268 58256 13320
rect 58308 13308 58314 13320
rect 58345 13311 58403 13317
rect 58345 13308 58357 13311
rect 58308 13280 58357 13308
rect 58308 13268 58314 13280
rect 58345 13277 58357 13280
rect 58391 13277 58403 13311
rect 58345 13271 58403 13277
rect 17828 13212 18000 13240
rect 17828 13200 17834 13212
rect 11054 13172 11060 13184
rect 2516 13144 11060 13172
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 17954 13132 17960 13184
rect 18012 13172 18018 13184
rect 19705 13175 19763 13181
rect 19705 13172 19717 13175
rect 18012 13144 19717 13172
rect 18012 13132 18018 13144
rect 19705 13141 19717 13144
rect 19751 13141 19763 13175
rect 19705 13135 19763 13141
rect 56134 13132 56140 13184
rect 56192 13172 56198 13184
rect 56505 13175 56563 13181
rect 56505 13172 56517 13175
rect 56192 13144 56517 13172
rect 56192 13132 56198 13144
rect 56505 13141 56517 13144
rect 56551 13141 56563 13175
rect 56505 13135 56563 13141
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 3602 12968 3608 12980
rect 2746 12940 3608 12968
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 2746 12832 2774 12940
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 9861 12971 9919 12977
rect 9861 12937 9873 12971
rect 9907 12968 9919 12971
rect 9950 12968 9956 12980
rect 9907 12940 9956 12968
rect 9907 12937 9919 12940
rect 9861 12931 9919 12937
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 13446 12928 13452 12980
rect 13504 12968 13510 12980
rect 22462 12968 22468 12980
rect 13504 12940 22468 12968
rect 13504 12928 13510 12940
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 22554 12928 22560 12980
rect 22612 12968 22618 12980
rect 22925 12971 22983 12977
rect 22925 12968 22937 12971
rect 22612 12940 22937 12968
rect 22612 12928 22618 12940
rect 22925 12937 22937 12940
rect 22971 12937 22983 12971
rect 22925 12931 22983 12937
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 23661 12971 23719 12977
rect 23661 12968 23673 12971
rect 23532 12940 23673 12968
rect 23532 12928 23538 12940
rect 23661 12937 23673 12940
rect 23707 12937 23719 12971
rect 23661 12931 23719 12937
rect 57146 12928 57152 12980
rect 57204 12968 57210 12980
rect 57425 12971 57483 12977
rect 57425 12968 57437 12971
rect 57204 12940 57437 12968
rect 57204 12928 57210 12940
rect 57425 12937 57437 12940
rect 57471 12937 57483 12971
rect 57425 12931 57483 12937
rect 3050 12900 3056 12912
rect 2963 12872 3056 12900
rect 3050 12860 3056 12872
rect 3108 12900 3114 12912
rect 5442 12900 5448 12912
rect 3108 12872 5448 12900
rect 3108 12860 3114 12872
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 8389 12903 8447 12909
rect 8389 12869 8401 12903
rect 8435 12900 8447 12903
rect 8478 12900 8484 12912
rect 8435 12872 8484 12900
rect 8435 12869 8447 12872
rect 8389 12863 8447 12869
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 9030 12860 9036 12912
rect 9088 12860 9094 12912
rect 11146 12832 11152 12844
rect 1903 12804 2774 12832
rect 11059 12804 11152 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 11146 12792 11152 12804
rect 11204 12832 11210 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11204 12804 11713 12832
rect 11204 12792 11210 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 20165 12835 20223 12841
rect 20165 12832 20177 12835
rect 19484 12804 20177 12832
rect 19484 12792 19490 12804
rect 20165 12801 20177 12804
rect 20211 12832 20223 12835
rect 20622 12832 20628 12844
rect 20211 12804 20628 12832
rect 20211 12801 20223 12804
rect 20165 12795 20223 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 22738 12792 22744 12844
rect 22796 12832 22802 12844
rect 22833 12835 22891 12841
rect 22833 12832 22845 12835
rect 22796 12804 22845 12832
rect 22796 12792 22802 12804
rect 22833 12801 22845 12804
rect 22879 12801 22891 12835
rect 22833 12795 22891 12801
rect 57698 12792 57704 12844
rect 57756 12832 57762 12844
rect 58342 12832 58348 12844
rect 57756 12804 58348 12832
rect 57756 12792 57762 12804
rect 58342 12792 58348 12804
rect 58400 12792 58406 12844
rect 2038 12724 2044 12776
rect 2096 12764 2102 12776
rect 2317 12767 2375 12773
rect 2317 12764 2329 12767
rect 2096 12736 2329 12764
rect 2096 12724 2102 12736
rect 2317 12733 2329 12736
rect 2363 12764 2375 12767
rect 4798 12764 4804 12776
rect 2363 12736 4804 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 8110 12764 8116 12776
rect 8071 12736 8116 12764
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 16574 12764 16580 12776
rect 8220 12736 16580 12764
rect 2406 12656 2412 12708
rect 2464 12696 2470 12708
rect 8220 12696 8248 12736
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 20257 12767 20315 12773
rect 20257 12764 20269 12767
rect 18708 12736 20269 12764
rect 2464 12668 8248 12696
rect 2464 12656 2470 12668
rect 11054 12656 11060 12708
rect 11112 12696 11118 12708
rect 11974 12696 11980 12708
rect 11112 12668 11980 12696
rect 11112 12656 11118 12668
rect 11974 12656 11980 12668
rect 12032 12696 12038 12708
rect 12032 12668 16574 12696
rect 12032 12656 12038 12668
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 2314 12588 2320 12640
rect 2372 12628 2378 12640
rect 3050 12628 3056 12640
rect 2372 12600 3056 12628
rect 2372 12588 2378 12600
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 12986 12628 12992 12640
rect 12947 12600 12992 12628
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 16546 12628 16574 12668
rect 18708 12637 18736 12736
rect 20257 12733 20269 12736
rect 20303 12733 20315 12767
rect 20438 12764 20444 12776
rect 20399 12736 20444 12764
rect 20257 12727 20315 12733
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 23109 12767 23167 12773
rect 23109 12733 23121 12767
rect 23155 12764 23167 12767
rect 23474 12764 23480 12776
rect 23155 12736 23480 12764
rect 23155 12733 23167 12736
rect 23109 12727 23167 12733
rect 23474 12724 23480 12736
rect 23532 12724 23538 12776
rect 18693 12631 18751 12637
rect 18693 12628 18705 12631
rect 16546 12600 18705 12628
rect 18693 12597 18705 12600
rect 18739 12597 18751 12631
rect 18693 12591 18751 12597
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 19426 12628 19432 12640
rect 19383 12600 19432 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 19426 12588 19432 12600
rect 19484 12588 19490 12640
rect 19794 12628 19800 12640
rect 19755 12600 19800 12628
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 22465 12631 22523 12637
rect 22465 12597 22477 12631
rect 22511 12628 22523 12631
rect 22646 12628 22652 12640
rect 22511 12600 22652 12628
rect 22511 12597 22523 12600
rect 22465 12591 22523 12597
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 58158 12628 58164 12640
rect 58119 12600 58164 12628
rect 58158 12588 58164 12600
rect 58216 12588 58222 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 3329 12427 3387 12433
rect 3329 12393 3341 12427
rect 3375 12424 3387 12427
rect 7573 12427 7631 12433
rect 7573 12424 7585 12427
rect 3375 12396 7585 12424
rect 3375 12393 3387 12396
rect 3329 12387 3387 12393
rect 7573 12393 7585 12396
rect 7619 12393 7631 12427
rect 7573 12387 7631 12393
rect 14918 12384 14924 12436
rect 14976 12424 14982 12436
rect 18782 12424 18788 12436
rect 14976 12396 18788 12424
rect 14976 12384 14982 12396
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 22462 12424 22468 12436
rect 22423 12396 22468 12424
rect 22462 12384 22468 12396
rect 22520 12384 22526 12436
rect 57698 12424 57704 12436
rect 57659 12396 57704 12424
rect 57698 12384 57704 12396
rect 57756 12384 57762 12436
rect 6089 12359 6147 12365
rect 6089 12356 6101 12359
rect 2056 12328 6101 12356
rect 1854 12180 1860 12232
rect 1912 12220 1918 12232
rect 2056 12220 2084 12328
rect 6089 12325 6101 12328
rect 6135 12325 6147 12359
rect 6089 12319 6147 12325
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2958 12288 2964 12300
rect 2179 12260 2964 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2958 12248 2964 12260
rect 3016 12288 3022 12300
rect 3973 12291 4031 12297
rect 3973 12288 3985 12291
rect 3016 12260 3985 12288
rect 3016 12248 3022 12260
rect 3973 12257 3985 12260
rect 4019 12257 4031 12291
rect 3973 12251 4031 12257
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 14936 12297 14964 12384
rect 14921 12291 14979 12297
rect 6972 12260 7880 12288
rect 6972 12248 6978 12260
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 1912 12192 2237 12220
rect 1912 12180 1918 12192
rect 2225 12189 2237 12192
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2314 12180 2320 12232
rect 2372 12220 2378 12232
rect 7852 12229 7880 12260
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12288 16727 12291
rect 17954 12288 17960 12300
rect 16715 12260 17960 12288
rect 16715 12257 16727 12260
rect 16669 12251 16727 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 3145 12223 3203 12229
rect 3145 12220 3157 12223
rect 2372 12192 2417 12220
rect 2700 12192 3157 12220
rect 2372 12180 2378 12192
rect 2700 12093 2728 12192
rect 3145 12189 3157 12192
rect 3191 12189 3203 12223
rect 3145 12183 3203 12189
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12220 7895 12223
rect 8110 12220 8116 12232
rect 7883 12192 8116 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 8110 12180 8116 12192
rect 8168 12220 8174 12232
rect 8294 12220 8300 12232
rect 8168 12192 8300 12220
rect 8168 12180 8174 12192
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 16945 12223 17003 12229
rect 16945 12189 16957 12223
rect 16991 12220 17003 12223
rect 17770 12220 17776 12232
rect 16991 12192 17776 12220
rect 16991 12189 17003 12192
rect 16945 12183 17003 12189
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 5408 12124 6394 12152
rect 5408 12112 5414 12124
rect 16206 12112 16212 12164
rect 16264 12112 16270 12164
rect 16758 12112 16764 12164
rect 16816 12152 16822 12164
rect 16960 12152 16988 12183
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 19794 12220 19800 12232
rect 19755 12192 19800 12220
rect 19794 12180 19800 12192
rect 19852 12180 19858 12232
rect 22646 12220 22652 12232
rect 22607 12192 22652 12220
rect 22646 12180 22652 12192
rect 22704 12180 22710 12232
rect 57149 12223 57207 12229
rect 57149 12189 57161 12223
rect 57195 12220 57207 12223
rect 58342 12220 58348 12232
rect 57195 12192 58348 12220
rect 57195 12189 57207 12192
rect 57149 12183 57207 12189
rect 58342 12180 58348 12192
rect 58400 12180 58406 12232
rect 16816 12124 16988 12152
rect 16816 12112 16822 12124
rect 2685 12087 2743 12093
rect 2685 12053 2697 12087
rect 2731 12053 2743 12087
rect 2685 12047 2743 12053
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 13354 12084 13360 12096
rect 10836 12056 13360 12084
rect 10836 12044 10842 12056
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 13504 12056 19625 12084
rect 13504 12044 13510 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 57606 12044 57612 12096
rect 57664 12084 57670 12096
rect 58161 12087 58219 12093
rect 58161 12084 58173 12087
rect 57664 12056 58173 12084
rect 57664 12044 57670 12056
rect 58161 12053 58173 12056
rect 58207 12053 58219 12087
rect 58161 12047 58219 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 2590 11880 2596 11892
rect 2363 11852 2596 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 11974 11880 11980 11892
rect 11935 11852 11980 11880
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 12216 11852 13124 11880
rect 12216 11840 12222 11852
rect 2409 11815 2467 11821
rect 2409 11781 2421 11815
rect 2455 11812 2467 11815
rect 3142 11812 3148 11824
rect 2455 11784 3148 11812
rect 2455 11781 2467 11784
rect 2409 11775 2467 11781
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 5350 11812 5356 11824
rect 5198 11784 5356 11812
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 9674 11772 9680 11824
rect 9732 11772 9738 11824
rect 10778 11812 10784 11824
rect 10739 11784 10784 11812
rect 10778 11772 10784 11784
rect 10836 11772 10842 11824
rect 13096 11812 13124 11852
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 19337 11883 19395 11889
rect 19337 11880 19349 11883
rect 13412 11852 19349 11880
rect 13412 11840 13418 11852
rect 19337 11849 19349 11852
rect 19383 11880 19395 11883
rect 20257 11883 20315 11889
rect 20257 11880 20269 11883
rect 19383 11852 20269 11880
rect 19383 11849 19395 11852
rect 19337 11843 19395 11849
rect 20257 11849 20269 11852
rect 20303 11849 20315 11883
rect 20257 11843 20315 11849
rect 56318 11840 56324 11892
rect 56376 11880 56382 11892
rect 57146 11880 57152 11892
rect 56376 11852 57152 11880
rect 56376 11840 56382 11852
rect 57146 11840 57152 11852
rect 57204 11840 57210 11892
rect 16666 11812 16672 11824
rect 13018 11784 16672 11812
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11744 5963 11747
rect 6914 11744 6920 11756
rect 5951 11716 6920 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11676 2283 11679
rect 2958 11676 2964 11688
rect 2271 11648 2964 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 2777 11611 2835 11617
rect 2777 11577 2789 11611
rect 2823 11608 2835 11611
rect 3252 11608 3280 11707
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 16206 11704 16212 11756
rect 16264 11744 16270 11756
rect 18138 11744 18144 11756
rect 16264 11716 18144 11744
rect 16264 11704 16270 11716
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 20070 11704 20076 11756
rect 20128 11744 20134 11756
rect 20165 11747 20223 11753
rect 20165 11744 20177 11747
rect 20128 11716 20177 11744
rect 20128 11704 20134 11716
rect 20165 11713 20177 11716
rect 20211 11713 20223 11747
rect 20165 11707 20223 11713
rect 22738 11704 22744 11756
rect 22796 11744 22802 11756
rect 22833 11747 22891 11753
rect 22833 11744 22845 11747
rect 22796 11716 22845 11744
rect 22796 11704 22802 11716
rect 22833 11713 22845 11716
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 56318 11704 56324 11756
rect 56376 11744 56382 11756
rect 56594 11744 56600 11756
rect 56376 11716 56421 11744
rect 56555 11716 56600 11744
rect 56376 11704 56382 11716
rect 56594 11704 56600 11716
rect 56652 11704 56658 11756
rect 57974 11744 57980 11756
rect 57256 11716 57980 11744
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 3436 11648 5641 11676
rect 3436 11617 3464 11648
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 5629 11639 5687 11645
rect 8294 11636 8300 11688
rect 8352 11676 8358 11688
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8352 11648 8769 11676
rect 8352 11636 8358 11648
rect 8757 11645 8769 11648
rect 8803 11645 8815 11679
rect 9030 11676 9036 11688
rect 8991 11648 9036 11676
rect 8757 11639 8815 11645
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 13446 11676 13452 11688
rect 13407 11648 13452 11676
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 13814 11676 13820 11688
rect 13771 11648 13820 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 20346 11636 20352 11688
rect 20404 11676 20410 11688
rect 22925 11679 22983 11685
rect 22925 11676 22937 11679
rect 20404 11648 20449 11676
rect 22066 11648 22937 11676
rect 20404 11636 20410 11648
rect 2823 11580 3280 11608
rect 3421 11611 3479 11617
rect 2823 11577 2835 11580
rect 2777 11571 2835 11577
rect 3421 11577 3433 11611
rect 3467 11577 3479 11611
rect 3421 11571 3479 11577
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 2648 11512 4169 11540
rect 2648 11500 2654 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 19797 11543 19855 11549
rect 19797 11509 19809 11543
rect 19843 11540 19855 11543
rect 19886 11540 19892 11552
rect 19843 11512 19892 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 21358 11540 21364 11552
rect 21319 11512 21364 11540
rect 21358 11500 21364 11512
rect 21416 11540 21422 11552
rect 22066 11540 22094 11648
rect 22925 11645 22937 11648
rect 22971 11645 22983 11679
rect 22925 11639 22983 11645
rect 23106 11636 23112 11688
rect 23164 11676 23170 11688
rect 23661 11679 23719 11685
rect 23661 11676 23673 11679
rect 23164 11648 23673 11676
rect 23164 11636 23170 11648
rect 23661 11645 23673 11648
rect 23707 11645 23719 11679
rect 23661 11639 23719 11645
rect 56480 11679 56538 11685
rect 56480 11645 56492 11679
rect 56526 11676 56538 11679
rect 57256 11676 57284 11716
rect 57974 11704 57980 11716
rect 58032 11704 58038 11756
rect 58342 11744 58348 11756
rect 58303 11716 58348 11744
rect 58342 11704 58348 11716
rect 58400 11704 58406 11756
rect 56526 11648 57284 11676
rect 57333 11679 57391 11685
rect 56526 11645 56538 11648
rect 56480 11639 56538 11645
rect 57333 11645 57345 11679
rect 57379 11645 57391 11679
rect 57333 11639 57391 11645
rect 57517 11679 57575 11685
rect 57517 11645 57529 11679
rect 57563 11676 57575 11679
rect 58066 11676 58072 11688
rect 57563 11648 58072 11676
rect 57563 11645 57575 11648
rect 57517 11639 57575 11645
rect 56870 11608 56876 11620
rect 56831 11580 56876 11608
rect 56870 11568 56876 11580
rect 56928 11568 56934 11620
rect 57348 11608 57376 11639
rect 58066 11636 58072 11648
rect 58124 11636 58130 11688
rect 57974 11608 57980 11620
rect 57348 11580 57980 11608
rect 57974 11568 57980 11580
rect 58032 11568 58038 11620
rect 21416 11512 22094 11540
rect 22465 11543 22523 11549
rect 21416 11500 21422 11512
rect 22465 11509 22477 11543
rect 22511 11540 22523 11543
rect 22554 11540 22560 11552
rect 22511 11512 22560 11540
rect 22511 11509 22523 11512
rect 22465 11503 22523 11509
rect 22554 11500 22560 11512
rect 22612 11500 22618 11552
rect 55306 11500 55312 11552
rect 55364 11540 55370 11552
rect 55677 11543 55735 11549
rect 55677 11540 55689 11543
rect 55364 11512 55689 11540
rect 55364 11500 55370 11512
rect 55677 11509 55689 11512
rect 55723 11509 55735 11543
rect 55677 11503 55735 11509
rect 55766 11500 55772 11552
rect 55824 11540 55830 11552
rect 58161 11543 58219 11549
rect 58161 11540 58173 11543
rect 55824 11512 58173 11540
rect 55824 11500 55830 11512
rect 58161 11509 58173 11512
rect 58207 11509 58219 11543
rect 58161 11503 58219 11509
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2593 11339 2651 11345
rect 2593 11305 2605 11339
rect 2639 11336 2651 11339
rect 2958 11336 2964 11348
rect 2639 11308 2964 11336
rect 2639 11305 2651 11308
rect 2593 11299 2651 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 9088 11308 19717 11336
rect 9088 11296 9094 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 20625 11339 20683 11345
rect 20625 11336 20637 11339
rect 20404 11308 20637 11336
rect 20404 11296 20410 11308
rect 20625 11305 20637 11308
rect 20671 11305 20683 11339
rect 57146 11336 57152 11348
rect 57107 11308 57152 11336
rect 20625 11299 20683 11305
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 2590 11132 2596 11144
rect 1903 11104 2596 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 2590 11092 2596 11104
rect 2648 11092 2654 11144
rect 3142 11132 3148 11144
rect 3103 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 19886 11132 19892 11144
rect 19847 11104 19892 11132
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20640 11132 20668 11299
rect 57146 11296 57152 11308
rect 57204 11296 57210 11348
rect 20714 11228 20720 11280
rect 20772 11268 20778 11280
rect 22373 11271 22431 11277
rect 22373 11268 22385 11271
rect 20772 11240 22385 11268
rect 20772 11228 20778 11240
rect 22373 11237 22385 11240
rect 22419 11237 22431 11271
rect 22373 11231 22431 11237
rect 56686 11228 56692 11280
rect 56744 11268 56750 11280
rect 58161 11271 58219 11277
rect 58161 11268 58173 11271
rect 56744 11240 58173 11268
rect 56744 11228 56750 11240
rect 58161 11237 58173 11240
rect 58207 11237 58219 11271
rect 58161 11231 58219 11237
rect 22186 11200 22192 11212
rect 22066 11172 22192 11200
rect 22066 11132 22094 11172
rect 22186 11160 22192 11172
rect 22244 11200 22250 11212
rect 23106 11200 23112 11212
rect 22244 11172 23112 11200
rect 22244 11160 22250 11172
rect 23106 11160 23112 11172
rect 23164 11160 23170 11212
rect 56870 11160 56876 11212
rect 56928 11200 56934 11212
rect 57609 11203 57667 11209
rect 57609 11200 57621 11203
rect 56928 11172 57621 11200
rect 56928 11160 56934 11172
rect 57609 11169 57621 11172
rect 57655 11169 57667 11203
rect 57609 11163 57667 11169
rect 22554 11132 22560 11144
rect 20640 11104 22094 11132
rect 22515 11104 22560 11132
rect 22554 11092 22560 11104
rect 22612 11092 22618 11144
rect 58345 11135 58403 11141
rect 58345 11101 58357 11135
rect 58391 11132 58403 11135
rect 58434 11132 58440 11144
rect 58391 11104 58440 11132
rect 58391 11101 58403 11104
rect 58345 11095 58403 11101
rect 58434 11092 58440 11104
rect 58492 11092 58498 11144
rect 2976 11036 3188 11064
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 2976 10996 3004 11036
rect 1544 10968 3004 10996
rect 3160 10996 3188 11036
rect 18874 10996 18880 11008
rect 3160 10968 18880 10996
rect 1544 10956 1550 10968
rect 18874 10956 18880 10968
rect 18932 10996 18938 11008
rect 21358 10996 21364 11008
rect 18932 10968 21364 10996
rect 18932 10956 18938 10968
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 20714 10792 20720 10804
rect 17144 10764 20720 10792
rect 9582 10724 9588 10736
rect 9495 10696 9588 10724
rect 9582 10684 9588 10696
rect 9640 10724 9646 10736
rect 12986 10724 12992 10736
rect 9640 10696 12992 10724
rect 9640 10684 9646 10696
rect 12986 10684 12992 10696
rect 13044 10684 13050 10736
rect 17144 10733 17172 10764
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 57514 10792 57520 10804
rect 57475 10764 57520 10792
rect 57514 10752 57520 10764
rect 57572 10752 57578 10804
rect 58342 10792 58348 10804
rect 58303 10764 58348 10792
rect 58342 10752 58348 10764
rect 58400 10752 58406 10804
rect 17129 10727 17187 10733
rect 17129 10693 17141 10727
rect 17175 10693 17187 10727
rect 17129 10687 17187 10693
rect 18138 10684 18144 10736
rect 18196 10684 18202 10736
rect 18874 10724 18880 10736
rect 18835 10696 18880 10724
rect 18874 10684 18880 10696
rect 18932 10684 18938 10736
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 1872 10588 1900 10619
rect 20070 10616 20076 10668
rect 20128 10656 20134 10668
rect 20257 10659 20315 10665
rect 20257 10656 20269 10659
rect 20128 10628 20269 10656
rect 20128 10616 20134 10628
rect 20257 10625 20269 10628
rect 20303 10625 20315 10659
rect 55306 10656 55312 10668
rect 55267 10628 55312 10656
rect 20257 10619 20315 10625
rect 55306 10616 55312 10628
rect 55364 10616 55370 10668
rect 2406 10588 2412 10600
rect 1872 10560 2412 10588
rect 2406 10548 2412 10560
rect 2464 10588 2470 10600
rect 10134 10588 10140 10600
rect 2464 10560 10140 10588
rect 2464 10548 2470 10560
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14737 10591 14795 10597
rect 14737 10588 14749 10591
rect 13872 10560 14749 10588
rect 13872 10548 13878 10560
rect 14737 10557 14749 10560
rect 14783 10588 14795 10591
rect 16758 10588 16764 10600
rect 14783 10560 16764 10588
rect 14783 10557 14795 10560
rect 14737 10551 14795 10557
rect 16758 10548 16764 10560
rect 16816 10588 16822 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16816 10560 16865 10588
rect 16816 10548 16822 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 20349 10591 20407 10597
rect 20349 10588 20361 10591
rect 16853 10551 16911 10557
rect 19352 10560 20361 10588
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 2590 10452 2596 10464
rect 2455 10424 2596 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2590 10412 2596 10424
rect 2648 10412 2654 10464
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 19352 10461 19380 10560
rect 20349 10557 20361 10560
rect 20395 10557 20407 10591
rect 20349 10551 20407 10557
rect 20438 10548 20444 10600
rect 20496 10588 20502 10600
rect 23382 10588 23388 10600
rect 20496 10560 23388 10588
rect 20496 10548 20502 10560
rect 23382 10548 23388 10560
rect 23440 10548 23446 10600
rect 19337 10455 19395 10461
rect 19337 10452 19349 10455
rect 16356 10424 19349 10452
rect 16356 10412 16362 10424
rect 19337 10421 19349 10424
rect 19383 10421 19395 10455
rect 19886 10452 19892 10464
rect 19847 10424 19892 10452
rect 19337 10415 19395 10421
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 51718 10412 51724 10464
rect 51776 10452 51782 10464
rect 55125 10455 55183 10461
rect 55125 10452 55137 10455
rect 51776 10424 55137 10452
rect 51776 10412 51782 10424
rect 55125 10421 55137 10424
rect 55171 10421 55183 10455
rect 55125 10415 55183 10421
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 12066 10248 12072 10260
rect 12027 10220 12072 10248
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 16298 10248 16304 10260
rect 16259 10220 16304 10248
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 57974 10140 57980 10192
rect 58032 10180 58038 10192
rect 58342 10180 58348 10192
rect 58032 10152 58348 10180
rect 58032 10140 58038 10152
rect 58342 10140 58348 10152
rect 58400 10140 58406 10192
rect 56876 10124 56928 10130
rect 16758 10072 16764 10124
rect 16816 10112 16822 10124
rect 18049 10115 18107 10121
rect 18049 10112 18061 10115
rect 16816 10084 18061 10112
rect 16816 10072 16822 10084
rect 18049 10081 18061 10084
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 23201 10115 23259 10121
rect 23201 10081 23213 10115
rect 23247 10112 23259 10115
rect 23382 10112 23388 10124
rect 23247 10084 23388 10112
rect 23247 10081 23259 10084
rect 23201 10075 23259 10081
rect 23382 10072 23388 10084
rect 23440 10072 23446 10124
rect 56876 10066 56928 10072
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 9490 10044 9496 10056
rect 1903 10016 9496 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 16666 10004 16672 10056
rect 16724 10004 16730 10056
rect 19886 10044 19892 10056
rect 19847 10016 19892 10044
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 57149 10047 57207 10053
rect 57149 10013 57161 10047
rect 57195 10044 57207 10047
rect 57974 10044 57980 10056
rect 57195 10016 57980 10044
rect 57195 10013 57207 10016
rect 57149 10007 57207 10013
rect 57974 10004 57980 10016
rect 58032 10004 58038 10056
rect 17773 9979 17831 9985
rect 17773 9945 17785 9979
rect 17819 9976 17831 9979
rect 17819 9948 19748 9976
rect 17819 9945 17831 9948
rect 17773 9939 17831 9945
rect 1670 9908 1676 9920
rect 1631 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 19720 9917 19748 9948
rect 22094 9936 22100 9988
rect 22152 9976 22158 9988
rect 23017 9979 23075 9985
rect 23017 9976 23029 9979
rect 22152 9948 23029 9976
rect 22152 9936 22158 9948
rect 23017 9945 23029 9948
rect 23063 9945 23075 9979
rect 23017 9939 23075 9945
rect 57054 9936 57060 9988
rect 57112 9976 57118 9988
rect 57517 9979 57575 9985
rect 57517 9976 57529 9979
rect 57112 9948 57529 9976
rect 57112 9936 57118 9948
rect 57517 9945 57529 9948
rect 57563 9945 57575 9979
rect 57517 9939 57575 9945
rect 57609 9979 57667 9985
rect 57609 9945 57621 9979
rect 57655 9945 57667 9979
rect 57609 9939 57667 9945
rect 57885 9979 57943 9985
rect 57885 9945 57897 9979
rect 57931 9976 57943 9979
rect 58158 9976 58164 9988
rect 57931 9948 58164 9976
rect 57931 9945 57943 9948
rect 57885 9939 57943 9945
rect 2961 9911 3019 9917
rect 2961 9908 2973 9911
rect 2832 9880 2973 9908
rect 2832 9868 2838 9880
rect 2961 9877 2973 9880
rect 3007 9877 3019 9911
rect 2961 9871 3019 9877
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9877 19763 9911
rect 19705 9871 19763 9877
rect 22557 9911 22615 9917
rect 22557 9877 22569 9911
rect 22603 9908 22615 9911
rect 22646 9908 22652 9920
rect 22603 9880 22652 9908
rect 22603 9877 22615 9880
rect 22557 9871 22615 9877
rect 22646 9868 22652 9880
rect 22704 9868 22710 9920
rect 22738 9868 22744 9920
rect 22796 9908 22802 9920
rect 22925 9911 22983 9917
rect 22925 9908 22937 9911
rect 22796 9880 22937 9908
rect 22796 9868 22802 9880
rect 22925 9877 22937 9880
rect 22971 9877 22983 9911
rect 22925 9871 22983 9877
rect 50154 9868 50160 9920
rect 50212 9908 50218 9920
rect 56597 9911 56655 9917
rect 56597 9908 56609 9911
rect 50212 9880 56609 9908
rect 50212 9868 50218 9880
rect 56597 9877 56609 9880
rect 56643 9877 56655 9911
rect 56597 9871 56655 9877
rect 56781 9911 56839 9917
rect 56781 9877 56793 9911
rect 56827 9908 56839 9911
rect 57330 9908 57336 9920
rect 56827 9880 57336 9908
rect 56827 9877 56839 9880
rect 56781 9871 56839 9877
rect 57330 9868 57336 9880
rect 57388 9868 57394 9920
rect 57422 9868 57428 9920
rect 57480 9908 57486 9920
rect 57624 9908 57652 9939
rect 58158 9936 58164 9948
rect 58216 9936 58222 9988
rect 57480 9880 57652 9908
rect 57480 9868 57486 9880
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 2501 9707 2559 9713
rect 2501 9673 2513 9707
rect 2547 9704 2559 9707
rect 2547 9676 2912 9704
rect 2547 9673 2559 9676
rect 2501 9667 2559 9673
rect 2774 9636 2780 9648
rect 2240 9608 2780 9636
rect 2240 9509 2268 9608
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 2884 9636 2912 9676
rect 40862 9664 40868 9716
rect 40920 9704 40926 9716
rect 50154 9704 50160 9716
rect 40920 9676 50160 9704
rect 40920 9664 40926 9676
rect 50154 9664 50160 9676
rect 50212 9664 50218 9716
rect 3786 9636 3792 9648
rect 2884 9608 3792 9636
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 55398 9596 55404 9648
rect 55456 9636 55462 9648
rect 55677 9639 55735 9645
rect 55677 9636 55689 9639
rect 55456 9608 55689 9636
rect 55456 9596 55462 9608
rect 55677 9605 55689 9608
rect 55723 9636 55735 9639
rect 56226 9636 56232 9648
rect 55723 9608 56232 9636
rect 55723 9605 55735 9608
rect 55677 9599 55735 9605
rect 56226 9596 56232 9608
rect 56284 9596 56290 9648
rect 56597 9639 56655 9645
rect 56597 9605 56609 9639
rect 56643 9636 56655 9639
rect 57054 9636 57060 9648
rect 56643 9608 57060 9636
rect 56643 9605 56655 9608
rect 56597 9599 56655 9605
rect 57054 9596 57060 9608
rect 57112 9596 57118 9648
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 2884 9540 3341 9568
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9469 2283 9503
rect 2406 9500 2412 9512
rect 2367 9472 2412 9500
rect 2225 9463 2283 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 2884 9441 2912 9540
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 6687 9540 7389 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7377 9537 7389 9540
rect 7423 9568 7435 9571
rect 11054 9568 11060 9580
rect 7423 9540 11060 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 11054 9528 11060 9540
rect 11112 9568 11118 9580
rect 12066 9568 12072 9580
rect 11112 9540 12072 9568
rect 11112 9528 11118 9540
rect 12066 9528 12072 9540
rect 12124 9568 12130 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 12124 9540 12173 9568
rect 12124 9528 12130 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 22646 9568 22652 9580
rect 22607 9540 22652 9568
rect 12161 9531 12219 9537
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 56870 9528 56876 9580
rect 56928 9568 56934 9580
rect 57425 9571 57483 9577
rect 57425 9568 57437 9571
rect 56928 9540 57437 9568
rect 56928 9528 56934 9540
rect 57425 9537 57437 9540
rect 57471 9537 57483 9571
rect 57425 9531 57483 9537
rect 57790 9528 57796 9580
rect 57848 9568 57854 9580
rect 58161 9571 58219 9577
rect 58161 9568 58173 9571
rect 57848 9540 58173 9568
rect 57848 9528 57854 9540
rect 58161 9537 58173 9540
rect 58207 9537 58219 9571
rect 58161 9531 58219 9537
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 9766 9500 9772 9512
rect 3476 9472 9772 9500
rect 3476 9460 3482 9472
rect 9766 9460 9772 9472
rect 9824 9500 9830 9512
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9824 9472 10057 9500
rect 9824 9460 9830 9472
rect 10045 9469 10057 9472
rect 10091 9500 10103 9503
rect 19426 9500 19432 9512
rect 10091 9472 19432 9500
rect 10091 9469 10103 9472
rect 10045 9463 10103 9469
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 2869 9435 2927 9441
rect 2869 9401 2881 9435
rect 2915 9401 2927 9435
rect 2869 9395 2927 9401
rect 5350 9392 5356 9444
rect 5408 9432 5414 9444
rect 6825 9435 6883 9441
rect 6825 9432 6837 9435
rect 5408 9404 6837 9432
rect 5408 9392 5414 9404
rect 6825 9401 6837 9404
rect 6871 9432 6883 9435
rect 8754 9432 8760 9444
rect 6871 9404 8760 9432
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 12158 9392 12164 9444
rect 12216 9432 12222 9444
rect 12345 9435 12403 9441
rect 12345 9432 12357 9435
rect 12216 9404 12357 9432
rect 12216 9392 12222 9404
rect 12345 9401 12357 9404
rect 12391 9432 12403 9435
rect 14826 9432 14832 9444
rect 12391 9404 14832 9432
rect 12391 9401 12403 9404
rect 12345 9395 12403 9401
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 14918 9392 14924 9444
rect 14976 9432 14982 9444
rect 22094 9432 22100 9444
rect 14976 9404 22100 9432
rect 14976 9392 14982 9404
rect 22094 9392 22100 9404
rect 22152 9392 22158 9444
rect 58250 9392 58256 9444
rect 58308 9432 58314 9444
rect 58345 9435 58403 9441
rect 58345 9432 58357 9435
rect 58308 9404 58357 9432
rect 58308 9392 58314 9404
rect 58345 9401 58357 9404
rect 58391 9401 58403 9435
rect 58345 9395 58403 9401
rect 3510 9364 3516 9376
rect 3471 9336 3516 9364
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 3973 9367 4031 9373
rect 3973 9364 3985 9367
rect 3844 9336 3985 9364
rect 3844 9324 3850 9336
rect 3973 9333 3985 9336
rect 4019 9333 4031 9367
rect 3973 9327 4031 9333
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 19518 9364 19524 9376
rect 13780 9336 19524 9364
rect 13780 9324 13786 9336
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19610 9324 19616 9376
rect 19668 9364 19674 9376
rect 22465 9367 22523 9373
rect 22465 9364 22477 9367
rect 19668 9336 22477 9364
rect 19668 9324 19674 9336
rect 22465 9333 22477 9336
rect 22511 9333 22523 9367
rect 22465 9327 22523 9333
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 4893 9163 4951 9169
rect 4893 9160 4905 9163
rect 2464 9132 4905 9160
rect 2464 9120 2470 9132
rect 4893 9129 4905 9132
rect 4939 9129 4951 9163
rect 4893 9123 4951 9129
rect 14461 9163 14519 9169
rect 14461 9129 14473 9163
rect 14507 9160 14519 9163
rect 14918 9160 14924 9172
rect 14507 9132 14924 9160
rect 14507 9129 14519 9132
rect 14461 9123 14519 9129
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15951 9163 16009 9169
rect 15951 9129 15963 9163
rect 15997 9160 16009 9163
rect 19610 9160 19616 9172
rect 15997 9132 19616 9160
rect 15997 9129 16009 9132
rect 15951 9123 16009 9129
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 20993 9163 21051 9169
rect 20993 9129 21005 9163
rect 21039 9160 21051 9163
rect 23474 9160 23480 9172
rect 21039 9132 23480 9160
rect 21039 9129 21051 9132
rect 20993 9123 21051 9129
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 9024 2467 9027
rect 2774 9024 2780 9036
rect 2455 8996 2780 9024
rect 2455 8993 2467 8996
rect 2409 8987 2467 8993
rect 2774 8984 2780 8996
rect 2832 9024 2838 9036
rect 3418 9024 3424 9036
rect 2832 8996 3424 9024
rect 2832 8984 2838 8996
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 6365 9027 6423 9033
rect 6365 9024 6377 9027
rect 3568 8996 6377 9024
rect 3568 8984 3574 8996
rect 6365 8993 6377 8996
rect 6411 8993 6423 9027
rect 6365 8987 6423 8993
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9585 9027 9643 9033
rect 9585 9024 9597 9027
rect 9548 8996 9597 9024
rect 9548 8984 9554 8996
rect 9585 8993 9597 8996
rect 9631 8993 9643 9027
rect 9766 9024 9772 9036
rect 9727 8996 9772 9024
rect 9585 8987 9643 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 10965 9027 11023 9033
rect 10965 8993 10977 9027
rect 11011 9024 11023 9027
rect 11238 9024 11244 9036
rect 11011 8996 11244 9024
rect 11011 8993 11023 8996
rect 10965 8987 11023 8993
rect 11238 8984 11244 8996
rect 11296 9024 11302 9036
rect 13722 9024 13728 9036
rect 11296 8996 13728 9024
rect 11296 8984 11302 8996
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 16209 9027 16267 9033
rect 16209 9024 16221 9027
rect 13832 8996 16221 9024
rect 13832 8968 13860 8996
rect 16209 8993 16221 8996
rect 16255 8993 16267 9027
rect 16209 8987 16267 8993
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 19576 8996 20177 9024
rect 19576 8984 19582 8996
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 9024 20407 9027
rect 21008 9024 21036 9123
rect 23474 9120 23480 9132
rect 23532 9120 23538 9172
rect 57149 9163 57207 9169
rect 57149 9129 57161 9163
rect 57195 9160 57207 9163
rect 57790 9160 57796 9172
rect 57195 9132 57796 9160
rect 57195 9129 57207 9132
rect 57149 9123 57207 9129
rect 57790 9120 57796 9132
rect 57848 9120 57854 9172
rect 58066 9120 58072 9172
rect 58124 9160 58130 9172
rect 58161 9163 58219 9169
rect 58161 9160 58173 9163
rect 58124 9132 58173 9160
rect 58124 9120 58130 9132
rect 58161 9129 58173 9132
rect 58207 9129 58219 9163
rect 58161 9123 58219 9129
rect 57054 9052 57060 9104
rect 57112 9092 57118 9104
rect 57609 9095 57667 9101
rect 57609 9092 57621 9095
rect 57112 9064 57621 9092
rect 57112 9052 57118 9064
rect 57609 9061 57621 9064
rect 57655 9061 57667 9095
rect 57609 9055 57667 9061
rect 20395 8996 21036 9024
rect 23109 9027 23167 9033
rect 20395 8993 20407 8996
rect 20349 8987 20407 8993
rect 23109 8993 23121 9027
rect 23155 9024 23167 9027
rect 23382 9024 23388 9036
rect 23155 8996 23388 9024
rect 23155 8993 23167 8996
rect 23109 8987 23167 8993
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 57624 9024 57652 9055
rect 57790 9024 57796 9036
rect 57624 8996 57796 9024
rect 57790 8984 57796 8996
rect 57848 8984 57854 9036
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 3142 8956 3148 8968
rect 2639 8928 3148 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 3142 8916 3148 8928
rect 3200 8956 3206 8968
rect 6641 8959 6699 8965
rect 3200 8928 3740 8956
rect 3200 8916 3206 8928
rect 3712 8832 3740 8928
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7374 8956 7380 8968
rect 6687 8928 7380 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 12989 8959 13047 8965
rect 8619 8928 9168 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 5350 8848 5356 8900
rect 5408 8848 5414 8900
rect 2498 8820 2504 8832
rect 2459 8792 2504 8820
rect 2498 8780 2504 8792
rect 2556 8780 2562 8832
rect 2958 8820 2964 8832
rect 2919 8792 2964 8820
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 3973 8823 4031 8829
rect 3973 8820 3985 8823
rect 3752 8792 3985 8820
rect 3752 8780 3758 8792
rect 3973 8789 3985 8792
rect 4019 8789 4031 8823
rect 3973 8783 4031 8789
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 9140 8829 9168 8928
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13814 8956 13820 8968
rect 13035 8928 13820 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 14826 8916 14832 8968
rect 14884 8916 14890 8968
rect 22462 8916 22468 8968
rect 22520 8956 22526 8968
rect 22833 8959 22891 8965
rect 22833 8956 22845 8959
rect 22520 8928 22845 8956
rect 22520 8916 22526 8928
rect 22833 8925 22845 8928
rect 22879 8925 22891 8959
rect 58342 8956 58348 8968
rect 58303 8928 58348 8956
rect 22833 8919 22891 8925
rect 58342 8916 58348 8928
rect 58400 8916 58406 8968
rect 9493 8891 9551 8897
rect 9493 8857 9505 8891
rect 9539 8888 9551 8891
rect 10318 8888 10324 8900
rect 9539 8860 10324 8888
rect 9539 8857 9551 8860
rect 9493 8851 9551 8857
rect 10318 8848 10324 8860
rect 10376 8888 10382 8900
rect 10376 8860 10456 8888
rect 10376 8848 10382 8860
rect 10428 8829 10456 8860
rect 12158 8848 12164 8900
rect 12216 8848 12222 8900
rect 12713 8891 12771 8897
rect 12713 8857 12725 8891
rect 12759 8888 12771 8891
rect 14642 8888 14648 8900
rect 12759 8860 14648 8888
rect 12759 8857 12771 8860
rect 12713 8851 12771 8857
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 22925 8891 22983 8897
rect 22925 8888 22937 8891
rect 22066 8860 22937 8888
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8352 8792 8401 8820
rect 8352 8780 8358 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 10413 8823 10471 8829
rect 10413 8789 10425 8823
rect 10459 8820 10471 8823
rect 10502 8820 10508 8832
rect 10459 8792 10508 8820
rect 10459 8789 10471 8792
rect 10413 8783 10471 8789
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 19705 8823 19763 8829
rect 19705 8789 19717 8823
rect 19751 8820 19763 8823
rect 19978 8820 19984 8832
rect 19751 8792 19984 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20070 8780 20076 8832
rect 20128 8820 20134 8832
rect 21910 8820 21916 8832
rect 20128 8792 20173 8820
rect 21871 8792 21916 8820
rect 20128 8780 20134 8792
rect 21910 8780 21916 8792
rect 21968 8820 21974 8832
rect 22066 8820 22094 8860
rect 22925 8857 22937 8860
rect 22971 8857 22983 8891
rect 22925 8851 22983 8857
rect 21968 8792 22094 8820
rect 22465 8823 22523 8829
rect 21968 8780 21974 8792
rect 22465 8789 22477 8823
rect 22511 8820 22523 8823
rect 22554 8820 22560 8832
rect 22511 8792 22560 8820
rect 22511 8789 22523 8792
rect 22465 8783 22523 8789
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 11701 8619 11759 8625
rect 11701 8616 11713 8619
rect 2648 8588 11713 8616
rect 2648 8576 2654 8588
rect 11701 8585 11713 8588
rect 11747 8585 11759 8619
rect 11701 8579 11759 8585
rect 18693 8619 18751 8625
rect 18693 8585 18705 8619
rect 18739 8585 18751 8619
rect 18693 8579 18751 8585
rect 3329 8551 3387 8557
rect 3329 8517 3341 8551
rect 3375 8548 3387 8551
rect 3418 8548 3424 8560
rect 3375 8520 3424 8548
rect 3375 8517 3387 8520
rect 3329 8511 3387 8517
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 8294 8548 8300 8560
rect 8255 8520 8300 8548
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 8754 8508 8760 8560
rect 8812 8508 8818 8560
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2406 8480 2412 8492
rect 1903 8452 2412 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8480 2651 8483
rect 2958 8480 2964 8492
rect 2639 8452 2964 8480
rect 2639 8449 2651 8452
rect 2593 8443 2651 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7432 8384 8033 8412
rect 7432 8372 7438 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 9548 8384 9781 8412
rect 9548 8372 9554 8384
rect 9769 8381 9781 8384
rect 9815 8381 9827 8415
rect 11716 8412 11744 8579
rect 12894 8548 12900 8560
rect 12742 8520 12900 8548
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 13173 8551 13231 8557
rect 13173 8517 13185 8551
rect 13219 8548 13231 8551
rect 18708 8548 18736 8579
rect 18782 8576 18788 8628
rect 18840 8616 18846 8628
rect 19242 8616 19248 8628
rect 18840 8588 19248 8616
rect 18840 8576 18846 8588
rect 19242 8576 19248 8588
rect 19300 8616 19306 8628
rect 19705 8619 19763 8625
rect 19705 8616 19717 8619
rect 19300 8588 19717 8616
rect 19300 8576 19306 8588
rect 19705 8585 19717 8588
rect 19751 8585 19763 8619
rect 19705 8579 19763 8585
rect 57517 8619 57575 8625
rect 57517 8585 57529 8619
rect 57563 8616 57575 8619
rect 58342 8616 58348 8628
rect 57563 8588 58348 8616
rect 57563 8585 57575 8588
rect 57517 8579 57575 8585
rect 58342 8576 58348 8588
rect 58400 8576 58406 8628
rect 19797 8551 19855 8557
rect 19797 8548 19809 8551
rect 13219 8520 18736 8548
rect 18800 8520 19809 8548
rect 13219 8517 13231 8520
rect 13173 8511 13231 8517
rect 13449 8415 13507 8421
rect 11716 8384 13400 8412
rect 9769 8375 9827 8381
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 6638 8344 6644 8356
rect 2823 8316 6644 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 13372 8344 13400 8384
rect 13449 8381 13461 8415
rect 13495 8412 13507 8415
rect 13814 8412 13820 8424
rect 13495 8384 13820 8412
rect 13495 8381 13507 8384
rect 13449 8375 13507 8381
rect 13814 8372 13820 8384
rect 13872 8412 13878 8424
rect 14366 8412 14372 8424
rect 13872 8384 14372 8412
rect 13872 8372 13878 8384
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 18800 8412 18828 8520
rect 19797 8517 19809 8520
rect 19843 8517 19855 8551
rect 19797 8511 19855 8517
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 22554 8480 22560 8492
rect 18923 8452 19380 8480
rect 22515 8452 22560 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 18156 8384 18828 8412
rect 18156 8353 18184 8384
rect 19352 8353 19380 8452
rect 22554 8440 22560 8452
rect 22612 8440 22618 8492
rect 56965 8483 57023 8489
rect 56965 8449 56977 8483
rect 57011 8480 57023 8483
rect 58342 8480 58348 8492
rect 57011 8452 58348 8480
rect 57011 8449 57023 8452
rect 56965 8443 57023 8449
rect 58342 8440 58348 8452
rect 58400 8440 58406 8492
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 19889 8415 19947 8421
rect 19889 8412 19901 8415
rect 19484 8384 19901 8412
rect 19484 8372 19490 8384
rect 19889 8381 19901 8384
rect 19935 8412 19947 8415
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 19935 8384 20545 8412
rect 19935 8381 19947 8384
rect 19889 8375 19947 8381
rect 20533 8381 20545 8384
rect 20579 8412 20591 8415
rect 20622 8412 20628 8424
rect 20579 8384 20628 8412
rect 20579 8381 20591 8384
rect 20533 8375 20591 8381
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 18141 8347 18199 8353
rect 18141 8344 18153 8347
rect 13372 8316 18153 8344
rect 18141 8313 18153 8316
rect 18187 8313 18199 8347
rect 18141 8307 18199 8313
rect 19337 8347 19395 8353
rect 19337 8313 19349 8347
rect 19383 8313 19395 8347
rect 19337 8307 19395 8313
rect 21726 8304 21732 8356
rect 21784 8344 21790 8356
rect 22373 8347 22431 8353
rect 22373 8344 22385 8347
rect 21784 8316 22385 8344
rect 21784 8304 21790 8316
rect 22373 8313 22385 8316
rect 22419 8313 22431 8347
rect 22373 8307 22431 8313
rect 57974 8304 57980 8356
rect 58032 8344 58038 8356
rect 58161 8347 58219 8353
rect 58161 8344 58173 8347
rect 58032 8316 58173 8344
rect 58032 8304 58038 8316
rect 58161 8313 58173 8316
rect 58207 8313 58219 8347
rect 58161 8307 58219 8313
rect 57422 8236 57428 8288
rect 57480 8276 57486 8288
rect 57698 8276 57704 8288
rect 57480 8248 57704 8276
rect 57480 8236 57486 8248
rect 57698 8236 57704 8248
rect 57756 8236 57762 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1670 8072 1676 8084
rect 1631 8044 1676 8072
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 3142 8072 3148 8084
rect 3055 8044 3148 8072
rect 3142 8032 3148 8044
rect 3200 8072 3206 8084
rect 3418 8072 3424 8084
rect 3200 8044 3424 8072
rect 3200 8032 3206 8044
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 19521 8075 19579 8081
rect 19521 8072 19533 8075
rect 14700 8044 19533 8072
rect 14700 8032 14706 8044
rect 19521 8041 19533 8044
rect 19567 8041 19579 8075
rect 19521 8035 19579 8041
rect 23385 8075 23443 8081
rect 23385 8041 23397 8075
rect 23431 8072 23443 8075
rect 23474 8072 23480 8084
rect 23431 8044 23480 8072
rect 23431 8041 23443 8044
rect 23385 8035 23443 8041
rect 18598 7964 18604 8016
rect 18656 8004 18662 8016
rect 21910 8004 21916 8016
rect 18656 7976 21916 8004
rect 18656 7964 18662 7976
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 2498 7936 2504 7948
rect 1872 7908 2504 7936
rect 1872 7877 1900 7908
rect 2498 7896 2504 7908
rect 2556 7936 2562 7948
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 2556 7908 5181 7936
rect 2556 7896 2562 7908
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 6638 7936 6644 7948
rect 6599 7908 6644 7936
rect 5169 7899 5227 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 22741 7939 22799 7945
rect 22741 7905 22753 7939
rect 22787 7936 22799 7939
rect 23400 7936 23428 8035
rect 23474 8032 23480 8044
rect 23532 8032 23538 8084
rect 58710 8072 58716 8084
rect 57256 8044 58716 8072
rect 56870 7964 56876 8016
rect 56928 8004 56934 8016
rect 57146 8004 57152 8016
rect 56928 7976 57152 8004
rect 56928 7964 56934 7976
rect 57146 7964 57152 7976
rect 57204 7964 57210 8016
rect 22787 7908 23428 7936
rect 57256 7936 57284 8044
rect 58710 8032 58716 8044
rect 58768 8032 58774 8084
rect 57606 7945 57612 7948
rect 57425 7939 57483 7945
rect 57425 7936 57437 7939
rect 57256 7908 57437 7936
rect 22787 7905 22799 7908
rect 22741 7899 22799 7905
rect 57425 7905 57437 7908
rect 57471 7905 57483 7939
rect 57425 7899 57483 7905
rect 57563 7939 57612 7945
rect 57563 7905 57575 7939
rect 57609 7905 57612 7939
rect 57563 7899 57612 7905
rect 57606 7896 57612 7899
rect 57664 7896 57670 7948
rect 57698 7896 57704 7948
rect 57756 7936 57762 7948
rect 57756 7908 57801 7936
rect 57756 7896 57762 7908
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2774 7868 2780 7880
rect 2639 7840 2780 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7374 7868 7380 7880
rect 6963 7840 7380 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 19978 7868 19984 7880
rect 19751 7840 19984 7868
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 56505 7871 56563 7877
rect 56505 7837 56517 7871
rect 56551 7868 56563 7871
rect 56594 7868 56600 7880
rect 56551 7840 56600 7868
rect 56551 7837 56563 7840
rect 56505 7831 56563 7837
rect 56594 7828 56600 7840
rect 56652 7828 56658 7880
rect 56689 7871 56747 7877
rect 56689 7837 56701 7871
rect 56735 7868 56747 7871
rect 56870 7868 56876 7880
rect 56735 7840 56876 7868
rect 56735 7837 56747 7840
rect 56689 7831 56747 7837
rect 56870 7828 56876 7840
rect 56928 7828 56934 7880
rect 6638 7800 6644 7812
rect 6210 7772 6644 7800
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 22557 7803 22615 7809
rect 22557 7800 22569 7803
rect 21560 7772 22569 7800
rect 21560 7744 21588 7772
rect 22557 7769 22569 7772
rect 22603 7769 22615 7803
rect 22557 7763 22615 7769
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 18782 7732 18788 7744
rect 18743 7704 18788 7732
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 21542 7732 21548 7744
rect 21503 7704 21548 7732
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 22094 7692 22100 7744
rect 22152 7732 22158 7744
rect 22462 7732 22468 7744
rect 22152 7704 22197 7732
rect 22423 7704 22468 7732
rect 22152 7692 22158 7704
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 58345 7735 58403 7741
rect 58345 7701 58357 7735
rect 58391 7732 58403 7735
rect 58434 7732 58440 7744
rect 58391 7704 58440 7732
rect 58391 7701 58403 7704
rect 58345 7695 58403 7701
rect 58434 7692 58440 7704
rect 58492 7692 58498 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7497 2927 7531
rect 3970 7528 3976 7540
rect 3931 7500 3976 7528
rect 2869 7491 2927 7497
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 2240 7364 2513 7392
rect 2240 7188 2268 7364
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2884 7392 2912 7491
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 18598 7528 18604 7540
rect 18559 7500 18604 7528
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 56594 7488 56600 7540
rect 56652 7528 56658 7540
rect 58161 7531 58219 7537
rect 58161 7528 58173 7531
rect 56652 7500 58173 7528
rect 56652 7488 56658 7500
rect 58161 7497 58173 7500
rect 58207 7497 58219 7531
rect 58161 7491 58219 7497
rect 9582 7460 9588 7472
rect 9543 7432 9588 7460
rect 9582 7420 9588 7432
rect 9640 7460 9646 7472
rect 12989 7463 13047 7469
rect 12989 7460 13001 7463
rect 9640 7432 13001 7460
rect 9640 7420 9646 7432
rect 12989 7429 13001 7432
rect 13035 7429 13047 7463
rect 12989 7423 13047 7429
rect 18138 7420 18144 7472
rect 18196 7420 18202 7472
rect 56962 7460 56968 7472
rect 56875 7432 56968 7460
rect 56962 7420 56968 7432
rect 57020 7460 57026 7472
rect 57698 7460 57704 7472
rect 57020 7432 57704 7460
rect 57020 7420 57026 7432
rect 57698 7420 57704 7432
rect 57756 7420 57762 7472
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 2884 7364 3341 7392
rect 2501 7355 2559 7361
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7392 22155 7395
rect 22830 7392 22836 7404
rect 22143 7364 22836 7392
rect 22143 7361 22155 7364
rect 22097 7355 22155 7361
rect 22830 7352 22836 7364
rect 22888 7392 22894 7404
rect 23109 7395 23167 7401
rect 23109 7392 23121 7395
rect 22888 7364 23121 7392
rect 22888 7352 22894 7364
rect 23109 7361 23121 7364
rect 23155 7361 23167 7395
rect 23753 7395 23811 7401
rect 23753 7392 23765 7395
rect 23109 7355 23167 7361
rect 23492 7364 23765 7392
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7293 2375 7327
rect 2317 7287 2375 7293
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7324 2467 7327
rect 2774 7324 2780 7336
rect 2455 7296 2780 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 2332 7256 2360 7287
rect 2774 7284 2780 7296
rect 2832 7324 2838 7336
rect 4062 7324 4068 7336
rect 2832 7296 4068 7324
rect 2832 7284 2838 7296
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7432 7296 7849 7324
rect 7432 7284 7438 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 14366 7284 14372 7336
rect 14424 7324 14430 7336
rect 14737 7327 14795 7333
rect 14737 7324 14749 7327
rect 14424 7296 14749 7324
rect 14424 7284 14430 7296
rect 14737 7293 14749 7296
rect 14783 7324 14795 7327
rect 16850 7324 16856 7336
rect 14783 7296 16856 7324
rect 14783 7293 14795 7296
rect 14737 7287 14795 7293
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7324 17187 7327
rect 21726 7324 21732 7336
rect 17175 7296 21732 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 21726 7284 21732 7296
rect 21784 7284 21790 7336
rect 23382 7324 23388 7336
rect 23343 7296 23388 7324
rect 23382 7284 23388 7296
rect 23440 7284 23446 7336
rect 2866 7256 2872 7268
rect 2332 7228 2872 7256
rect 2866 7216 2872 7228
rect 2924 7256 2930 7268
rect 3142 7256 3148 7268
rect 2924 7228 3148 7256
rect 2924 7216 2930 7228
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 3970 7256 3976 7268
rect 3344 7228 3976 7256
rect 3344 7188 3372 7228
rect 3970 7216 3976 7228
rect 4028 7216 4034 7268
rect 23492 7256 23520 7364
rect 23753 7361 23765 7364
rect 23799 7361 23811 7395
rect 23753 7355 23811 7361
rect 56413 7395 56471 7401
rect 56413 7361 56425 7395
rect 56459 7392 56471 7395
rect 58342 7392 58348 7404
rect 56459 7364 58348 7392
rect 56459 7361 56471 7364
rect 56413 7355 56471 7361
rect 58342 7352 58348 7364
rect 58400 7352 58406 7404
rect 57146 7284 57152 7336
rect 57204 7324 57210 7336
rect 57425 7327 57483 7333
rect 57425 7324 57437 7327
rect 57204 7296 57437 7324
rect 57204 7284 57210 7296
rect 57425 7293 57437 7296
rect 57471 7293 57483 7327
rect 57425 7287 57483 7293
rect 23124 7228 23520 7256
rect 23124 7200 23152 7228
rect 3510 7188 3516 7200
rect 2240 7160 3372 7188
rect 3471 7160 3516 7188
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 19150 7188 19156 7200
rect 19111 7160 19156 7188
rect 19150 7148 19156 7160
rect 19208 7148 19214 7200
rect 22649 7191 22707 7197
rect 22649 7157 22661 7191
rect 22695 7188 22707 7191
rect 23106 7188 23112 7200
rect 22695 7160 23112 7188
rect 22695 7157 22707 7160
rect 22649 7151 22707 7157
rect 23106 7148 23112 7160
rect 23164 7148 23170 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 3510 6944 3516 6996
rect 3568 6984 3574 6996
rect 5549 6987 5607 6993
rect 5549 6984 5561 6987
rect 3568 6956 5561 6984
rect 3568 6944 3574 6956
rect 5549 6953 5561 6956
rect 5595 6953 5607 6987
rect 23474 6984 23480 6996
rect 23435 6956 23480 6984
rect 5549 6947 5607 6953
rect 23474 6944 23480 6956
rect 23532 6944 23538 6996
rect 56318 6944 56324 6996
rect 56376 6984 56382 6996
rect 56962 6984 56968 6996
rect 56376 6956 56968 6984
rect 56376 6944 56382 6956
rect 56962 6944 56968 6956
rect 57020 6944 57026 6996
rect 4062 6916 4068 6928
rect 4023 6888 4068 6916
rect 4062 6876 4068 6888
rect 4120 6876 4126 6928
rect 56873 6919 56931 6925
rect 56873 6885 56885 6919
rect 56919 6916 56931 6919
rect 57146 6916 57152 6928
rect 56919 6888 57152 6916
rect 56919 6885 56931 6888
rect 56873 6879 56931 6885
rect 57146 6876 57152 6888
rect 57204 6916 57210 6928
rect 57330 6916 57336 6928
rect 57204 6888 57336 6916
rect 57204 6876 57210 6888
rect 57330 6876 57336 6888
rect 57388 6876 57394 6928
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 2866 6848 2872 6860
rect 2271 6820 2872 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 3234 6848 3240 6860
rect 3195 6820 3240 6848
rect 3234 6808 3240 6820
rect 3292 6808 3298 6860
rect 10134 6808 10140 6860
rect 10192 6848 10198 6860
rect 19150 6848 19156 6860
rect 10192 6820 19156 6848
rect 10192 6808 10198 6820
rect 19150 6808 19156 6820
rect 19208 6848 19214 6860
rect 19889 6851 19947 6857
rect 19889 6848 19901 6851
rect 19208 6820 19901 6848
rect 19208 6808 19214 6820
rect 19889 6817 19901 6820
rect 19935 6817 19947 6851
rect 19889 6811 19947 6817
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6848 20131 6851
rect 20622 6848 20628 6860
rect 20119 6820 20628 6848
rect 20119 6817 20131 6820
rect 20073 6811 20131 6817
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 22005 6851 22063 6857
rect 22005 6817 22017 6851
rect 22051 6848 22063 6851
rect 22186 6848 22192 6860
rect 22051 6820 22192 6848
rect 22051 6817 22063 6820
rect 22005 6811 22063 6817
rect 22186 6808 22192 6820
rect 22244 6808 22250 6860
rect 56318 6848 56324 6860
rect 56279 6820 56324 6848
rect 56318 6808 56324 6820
rect 56376 6808 56382 6860
rect 56597 6851 56655 6857
rect 56597 6817 56609 6851
rect 56643 6848 56655 6851
rect 56778 6848 56784 6860
rect 56643 6820 56784 6848
rect 56643 6817 56655 6820
rect 56597 6811 56655 6817
rect 56778 6808 56784 6820
rect 56836 6808 56842 6860
rect 2409 6715 2467 6721
rect 2409 6681 2421 6715
rect 2455 6712 2467 6715
rect 3252 6712 3280 6808
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 4062 6780 4068 6792
rect 3752 6752 4068 6780
rect 3752 6740 3758 6752
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 7374 6780 7380 6792
rect 5859 6752 7380 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15930 6780 15936 6792
rect 15528 6752 15936 6780
rect 15528 6740 15534 6752
rect 15930 6740 15936 6752
rect 15988 6780 15994 6792
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 15988 6752 18797 6780
rect 15988 6740 15994 6752
rect 18785 6749 18797 6752
rect 18831 6780 18843 6783
rect 19797 6783 19855 6789
rect 19797 6780 19809 6783
rect 18831 6752 19809 6780
rect 18831 6749 18843 6752
rect 18785 6743 18843 6749
rect 19797 6749 19809 6752
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6780 21419 6783
rect 22094 6780 22100 6792
rect 21407 6752 22100 6780
rect 21407 6749 21419 6752
rect 21361 6743 21419 6749
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 22830 6740 22836 6792
rect 22888 6780 22894 6792
rect 23017 6783 23075 6789
rect 23017 6780 23029 6783
rect 22888 6752 23029 6780
rect 22888 6740 22894 6752
rect 23017 6749 23029 6752
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 23106 6740 23112 6792
rect 23164 6780 23170 6792
rect 23937 6783 23995 6789
rect 23937 6780 23949 6783
rect 23164 6752 23949 6780
rect 23164 6740 23170 6752
rect 23937 6749 23949 6752
rect 23983 6780 23995 6783
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 23983 6752 24593 6780
rect 23983 6749 23995 6752
rect 23937 6743 23995 6749
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 56410 6740 56416 6792
rect 56468 6789 56474 6792
rect 56468 6783 56517 6789
rect 56468 6749 56471 6783
rect 56505 6749 56517 6783
rect 56468 6743 56517 6749
rect 56468 6740 56474 6743
rect 57146 6740 57152 6792
rect 57204 6780 57210 6792
rect 57333 6783 57391 6789
rect 57333 6780 57345 6783
rect 57204 6752 57345 6780
rect 57204 6740 57210 6752
rect 57333 6749 57345 6752
rect 57379 6749 57391 6783
rect 57333 6743 57391 6749
rect 57517 6783 57575 6789
rect 57517 6749 57529 6783
rect 57563 6749 57575 6783
rect 58342 6780 58348 6792
rect 58303 6752 58348 6780
rect 57517 6743 57575 6749
rect 3510 6712 3516 6724
rect 2455 6684 3516 6712
rect 2455 6681 2467 6684
rect 2409 6675 2467 6681
rect 3510 6672 3516 6684
rect 3568 6672 3574 6724
rect 6638 6712 6644 6724
rect 5106 6684 6644 6712
rect 6638 6672 6644 6684
rect 6696 6672 6702 6724
rect 13906 6672 13912 6724
rect 13964 6712 13970 6724
rect 21542 6712 21548 6724
rect 13964 6684 21548 6712
rect 13964 6672 13970 6684
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 22189 6715 22247 6721
rect 22189 6681 22201 6715
rect 22235 6712 22247 6715
rect 22462 6712 22468 6724
rect 22235 6684 22468 6712
rect 22235 6681 22247 6684
rect 22189 6675 22247 6681
rect 22462 6672 22468 6684
rect 22520 6672 22526 6724
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2556 6616 2789 6644
rect 2556 6604 2562 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 2777 6607 2835 6613
rect 15102 6604 15108 6656
rect 15160 6644 15166 6656
rect 18138 6644 18144 6656
rect 15160 6616 18144 6644
rect 15160 6604 15166 6616
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 19426 6644 19432 6656
rect 19387 6616 19432 6644
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 21174 6644 21180 6656
rect 21135 6616 21180 6644
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 22554 6644 22560 6656
rect 22152 6616 22197 6644
rect 22515 6616 22560 6644
rect 22152 6604 22158 6616
rect 22554 6604 22560 6616
rect 22612 6604 22618 6656
rect 55582 6604 55588 6656
rect 55640 6644 55646 6656
rect 55677 6647 55735 6653
rect 55677 6644 55689 6647
rect 55640 6616 55689 6644
rect 55640 6604 55646 6616
rect 55677 6613 55689 6616
rect 55723 6613 55735 6647
rect 55677 6607 55735 6613
rect 55766 6604 55772 6656
rect 55824 6644 55830 6656
rect 56410 6644 56416 6656
rect 55824 6616 56416 6644
rect 55824 6604 55830 6616
rect 56410 6604 56416 6616
rect 56468 6604 56474 6656
rect 57532 6644 57560 6743
rect 58342 6740 58348 6752
rect 58400 6740 58406 6792
rect 58161 6647 58219 6653
rect 58161 6644 58173 6647
rect 57532 6616 58173 6644
rect 58161 6613 58173 6616
rect 58207 6613 58219 6647
rect 58161 6607 58219 6613
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2866 6400 2872 6452
rect 2924 6440 2930 6452
rect 3145 6443 3203 6449
rect 3145 6440 3157 6443
rect 2924 6412 3157 6440
rect 2924 6400 2930 6412
rect 3145 6409 3157 6412
rect 3191 6409 3203 6443
rect 21361 6443 21419 6449
rect 21361 6440 21373 6443
rect 3145 6403 3203 6409
rect 7852 6412 21373 6440
rect 7466 6332 7472 6384
rect 7524 6372 7530 6384
rect 7852 6381 7880 6412
rect 21361 6409 21373 6412
rect 21407 6440 21419 6443
rect 22094 6440 22100 6452
rect 21407 6412 22100 6440
rect 21407 6409 21419 6412
rect 21361 6403 21419 6409
rect 22094 6400 22100 6412
rect 22152 6400 22158 6452
rect 56962 6440 56968 6452
rect 56923 6412 56968 6440
rect 56962 6400 56968 6412
rect 57020 6400 57026 6452
rect 57330 6400 57336 6452
rect 57388 6440 57394 6452
rect 57425 6443 57483 6449
rect 57425 6440 57437 6443
rect 57388 6412 57437 6440
rect 57388 6400 57394 6412
rect 57425 6409 57437 6412
rect 57471 6409 57483 6443
rect 57425 6403 57483 6409
rect 58342 6400 58348 6452
rect 58400 6400 58406 6452
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 7524 6344 7849 6372
rect 7524 6332 7530 6344
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 9674 6372 9680 6384
rect 9154 6344 9680 6372
rect 7837 6335 7895 6341
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 13817 6375 13875 6381
rect 13817 6341 13829 6375
rect 13863 6372 13875 6375
rect 13906 6372 13912 6384
rect 13863 6344 13912 6372
rect 13863 6341 13875 6344
rect 13817 6335 13875 6341
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 15102 6332 15108 6384
rect 15160 6332 15166 6384
rect 15565 6375 15623 6381
rect 15565 6341 15577 6375
rect 15611 6372 15623 6375
rect 21174 6372 21180 6384
rect 15611 6344 21180 6372
rect 15611 6341 15623 6344
rect 15565 6335 15623 6341
rect 21174 6332 21180 6344
rect 21232 6332 21238 6384
rect 56413 6375 56471 6381
rect 56413 6341 56425 6375
rect 56459 6372 56471 6375
rect 58360 6372 58388 6400
rect 56459 6344 58388 6372
rect 56459 6341 56471 6344
rect 56413 6335 56471 6341
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2314 6304 2320 6316
rect 1903 6276 2320 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 2498 6304 2504 6316
rect 2459 6276 2504 6304
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 19426 6304 19432 6316
rect 19387 6276 19432 6304
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19794 6264 19800 6316
rect 19852 6304 19858 6316
rect 20073 6307 20131 6313
rect 20073 6304 20085 6307
rect 19852 6276 20085 6304
rect 19852 6264 19858 6276
rect 20073 6273 20085 6276
rect 20119 6273 20131 6307
rect 22554 6304 22560 6316
rect 22515 6276 22560 6304
rect 20073 6267 20131 6273
rect 22554 6264 22560 6276
rect 22612 6264 22618 6316
rect 22830 6264 22836 6316
rect 22888 6304 22894 6316
rect 23017 6307 23075 6313
rect 23017 6304 23029 6307
rect 22888 6276 23029 6304
rect 22888 6264 22894 6276
rect 23017 6273 23029 6276
rect 23063 6273 23075 6307
rect 23017 6267 23075 6273
rect 23106 6264 23112 6316
rect 23164 6304 23170 6316
rect 23569 6307 23627 6313
rect 23569 6304 23581 6307
rect 23164 6276 23581 6304
rect 23164 6264 23170 6276
rect 23569 6273 23581 6276
rect 23615 6304 23627 6307
rect 24213 6307 24271 6313
rect 24213 6304 24225 6307
rect 23615 6276 24225 6304
rect 23615 6273 23627 6276
rect 23569 6267 23627 6273
rect 24213 6273 24225 6276
rect 24259 6273 24271 6307
rect 24213 6267 24271 6273
rect 55861 6307 55919 6313
rect 55861 6273 55873 6307
rect 55907 6304 55919 6307
rect 58342 6304 58348 6316
rect 55907 6276 58348 6304
rect 55907 6273 55919 6276
rect 55861 6267 55919 6273
rect 58342 6264 58348 6276
rect 58400 6264 58406 6316
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 9548 6208 9597 6236
rect 9548 6196 9554 6208
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9585 6199 9643 6205
rect 9784 6208 9873 6236
rect 2682 6100 2688 6112
rect 2643 6072 2688 6100
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 9784 6100 9812 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16850 6236 16856 6248
rect 15887 6208 16856 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16850 6196 16856 6208
rect 16908 6236 16914 6248
rect 18598 6236 18604 6248
rect 16908 6208 18604 6236
rect 16908 6196 16914 6208
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 16942 6128 16948 6180
rect 17000 6168 17006 6180
rect 22373 6171 22431 6177
rect 22373 6168 22385 6171
rect 17000 6140 22385 6168
rect 17000 6128 17006 6140
rect 22373 6137 22385 6140
rect 22419 6137 22431 6171
rect 22373 6131 22431 6137
rect 44818 6128 44824 6180
rect 44876 6168 44882 6180
rect 53098 6168 53104 6180
rect 44876 6140 53104 6168
rect 44876 6128 44882 6140
rect 53098 6128 53104 6140
rect 53156 6128 53162 6180
rect 56778 6128 56784 6180
rect 56836 6168 56842 6180
rect 57330 6168 57336 6180
rect 56836 6140 57336 6168
rect 56836 6128 56842 6140
rect 57330 6128 57336 6140
rect 57388 6128 57394 6180
rect 9640 6072 9812 6100
rect 9640 6060 9646 6072
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 11664 6072 19257 6100
rect 11664 6060 11670 6072
rect 19245 6069 19257 6072
rect 19291 6069 19303 6103
rect 19245 6063 19303 6069
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19889 6103 19947 6109
rect 19889 6100 19901 6103
rect 19392 6072 19901 6100
rect 19392 6060 19398 6072
rect 19889 6069 19901 6072
rect 19935 6069 19947 6103
rect 19889 6063 19947 6069
rect 22186 6060 22192 6112
rect 22244 6100 22250 6112
rect 22646 6100 22652 6112
rect 22244 6072 22652 6100
rect 22244 6060 22250 6072
rect 22646 6060 22652 6072
rect 22704 6100 22710 6112
rect 23109 6103 23167 6109
rect 23109 6100 23121 6103
rect 22704 6072 23121 6100
rect 22704 6060 22710 6072
rect 23109 6069 23121 6072
rect 23155 6069 23167 6103
rect 23109 6063 23167 6069
rect 57054 6060 57060 6112
rect 57112 6100 57118 6112
rect 58161 6103 58219 6109
rect 58161 6100 58173 6103
rect 57112 6072 58173 6100
rect 57112 6060 57118 6072
rect 58161 6069 58173 6072
rect 58207 6069 58219 6103
rect 58161 6063 58219 6069
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1670 5896 1676 5908
rect 1631 5868 1676 5896
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 2740 5868 5764 5896
rect 2740 5856 2746 5868
rect 2314 5788 2320 5840
rect 2372 5828 2378 5840
rect 5629 5831 5687 5837
rect 5629 5828 5641 5831
rect 2372 5800 5641 5828
rect 2372 5788 2378 5800
rect 5629 5797 5641 5800
rect 5675 5797 5687 5831
rect 5629 5791 5687 5797
rect 5736 5760 5764 5868
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 16942 5896 16948 5908
rect 9548 5868 16948 5896
rect 9548 5856 9554 5868
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 19794 5896 19800 5908
rect 19755 5868 19800 5896
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 22646 5896 22652 5908
rect 22607 5868 22652 5896
rect 22646 5856 22652 5868
rect 22704 5856 22710 5908
rect 56686 5856 56692 5908
rect 56744 5896 56750 5908
rect 57606 5896 57612 5908
rect 56744 5868 57612 5896
rect 56744 5856 56750 5868
rect 57606 5856 57612 5868
rect 57664 5856 57670 5908
rect 10134 5828 10140 5840
rect 10095 5800 10140 5828
rect 10134 5788 10140 5800
rect 10192 5788 10198 5840
rect 16574 5788 16580 5840
rect 16632 5828 16638 5840
rect 16761 5831 16819 5837
rect 16761 5828 16773 5831
rect 16632 5800 16773 5828
rect 16632 5788 16638 5800
rect 16761 5797 16773 5800
rect 16807 5797 16819 5831
rect 16761 5791 16819 5797
rect 56778 5788 56784 5840
rect 56836 5828 56842 5840
rect 57149 5831 57207 5837
rect 57149 5828 57161 5831
rect 56836 5800 57161 5828
rect 56836 5788 56842 5800
rect 57149 5797 57161 5800
rect 57195 5828 57207 5831
rect 57238 5828 57244 5840
rect 57195 5800 57244 5828
rect 57195 5797 57207 5800
rect 57149 5791 57207 5797
rect 57238 5788 57244 5800
rect 57296 5788 57302 5840
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 5736 5732 7113 5760
rect 7101 5729 7113 5732
rect 7147 5729 7159 5763
rect 7374 5760 7380 5772
rect 7287 5732 7380 5760
rect 7101 5723 7159 5729
rect 7374 5720 7380 5732
rect 7432 5760 7438 5772
rect 9582 5760 9588 5772
rect 7432 5732 9588 5760
rect 7432 5720 7438 5732
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 11606 5760 11612 5772
rect 11567 5732 11612 5760
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 20438 5760 20444 5772
rect 20399 5732 20444 5760
rect 20438 5720 20444 5732
rect 20496 5720 20502 5772
rect 56505 5763 56563 5769
rect 56505 5729 56517 5763
rect 56551 5760 56563 5763
rect 57054 5760 57060 5772
rect 56551 5732 57060 5760
rect 56551 5729 56563 5732
rect 56505 5723 56563 5729
rect 57054 5720 57060 5732
rect 57112 5720 57118 5772
rect 57422 5760 57428 5772
rect 57383 5732 57428 5760
rect 57422 5720 57428 5732
rect 57480 5720 57486 5772
rect 57606 5769 57612 5772
rect 57563 5763 57612 5769
rect 57563 5729 57575 5763
rect 57609 5729 57612 5763
rect 57563 5723 57612 5729
rect 57606 5720 57612 5723
rect 57664 5720 57670 5772
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2590 5692 2596 5704
rect 1903 5664 2596 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 14366 5692 14372 5704
rect 11931 5664 14372 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 18598 5692 18604 5704
rect 18555 5664 18604 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 20162 5692 20168 5704
rect 19484 5664 20168 5692
rect 19484 5652 19490 5664
rect 20162 5652 20168 5664
rect 20220 5652 20226 5704
rect 56686 5692 56692 5704
rect 56647 5664 56692 5692
rect 56686 5652 56692 5664
rect 56744 5652 56750 5704
rect 57698 5692 57704 5704
rect 57659 5664 57704 5692
rect 57698 5652 57704 5664
rect 57756 5652 57762 5704
rect 6638 5584 6644 5636
rect 6696 5624 6702 5636
rect 9674 5624 9680 5636
rect 6696 5596 9680 5624
rect 6696 5584 6702 5596
rect 9674 5584 9680 5596
rect 9732 5624 9738 5636
rect 10318 5624 10324 5636
rect 9732 5596 10324 5624
rect 9732 5584 9738 5596
rect 10318 5584 10324 5596
rect 10376 5624 10382 5636
rect 18230 5624 18236 5636
rect 10376 5596 10442 5624
rect 17802 5596 17908 5624
rect 18191 5596 18236 5624
rect 10376 5584 10382 5596
rect 17586 5516 17592 5568
rect 17644 5556 17650 5568
rect 17880 5556 17908 5596
rect 18230 5584 18236 5596
rect 18288 5584 18294 5636
rect 18138 5556 18144 5568
rect 17644 5528 18144 5556
rect 17644 5516 17650 5528
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 20254 5516 20260 5568
rect 20312 5556 20318 5568
rect 20993 5559 21051 5565
rect 20993 5556 21005 5559
rect 20312 5528 21005 5556
rect 20312 5516 20318 5528
rect 20993 5525 21005 5528
rect 21039 5525 21051 5559
rect 20993 5519 21051 5525
rect 22830 5516 22836 5568
rect 22888 5556 22894 5568
rect 23201 5559 23259 5565
rect 23201 5556 23213 5559
rect 22888 5528 23213 5556
rect 22888 5516 22894 5528
rect 23201 5525 23213 5528
rect 23247 5525 23259 5559
rect 23201 5519 23259 5525
rect 56962 5516 56968 5568
rect 57020 5556 57026 5568
rect 57698 5556 57704 5568
rect 57020 5528 57704 5556
rect 57020 5516 57026 5528
rect 57698 5516 57704 5528
rect 57756 5516 57762 5568
rect 58250 5516 58256 5568
rect 58308 5556 58314 5568
rect 58345 5559 58403 5565
rect 58345 5556 58357 5559
rect 58308 5528 58357 5556
rect 58308 5516 58314 5528
rect 58345 5525 58357 5528
rect 58391 5525 58403 5559
rect 58345 5519 58403 5525
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 4798 5312 4804 5364
rect 4856 5352 4862 5364
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 4856 5324 11897 5352
rect 4856 5312 4862 5324
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 13630 5352 13636 5364
rect 11885 5315 11943 5321
rect 13280 5324 13636 5352
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 2682 5216 2688 5228
rect 1903 5188 2688 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 1670 5080 1676 5092
rect 1631 5052 1676 5080
rect 1670 5040 1676 5052
rect 1728 5040 1734 5092
rect 11900 5012 11928 5315
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 13280 5284 13308 5324
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 18230 5312 18236 5364
rect 18288 5352 18294 5364
rect 19245 5355 19303 5361
rect 19245 5352 19257 5355
rect 18288 5324 19257 5352
rect 18288 5312 18294 5324
rect 19245 5321 19257 5324
rect 19291 5321 19303 5355
rect 19245 5315 19303 5321
rect 20257 5355 20315 5361
rect 20257 5321 20269 5355
rect 20303 5352 20315 5355
rect 20346 5352 20352 5364
rect 20303 5324 20352 5352
rect 20303 5321 20315 5324
rect 20257 5315 20315 5321
rect 20346 5312 20352 5324
rect 20404 5352 20410 5364
rect 20530 5352 20536 5364
rect 20404 5324 20536 5352
rect 20404 5312 20410 5324
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 56962 5352 56968 5364
rect 56923 5324 56968 5352
rect 56962 5312 56968 5324
rect 57020 5312 57026 5364
rect 57238 5312 57244 5364
rect 57296 5352 57302 5364
rect 57425 5355 57483 5361
rect 57425 5352 57437 5355
rect 57296 5324 57437 5352
rect 57296 5312 57302 5324
rect 57425 5321 57437 5324
rect 57471 5321 57483 5355
rect 57425 5315 57483 5321
rect 58161 5355 58219 5361
rect 58161 5321 58173 5355
rect 58207 5352 58219 5355
rect 58526 5352 58532 5364
rect 58207 5324 58532 5352
rect 58207 5321 58219 5324
rect 58161 5315 58219 5321
rect 58526 5312 58532 5324
rect 58584 5312 58590 5364
rect 12952 5256 13308 5284
rect 13357 5287 13415 5293
rect 12952 5244 12958 5256
rect 13357 5253 13369 5287
rect 13403 5284 13415 5287
rect 19334 5284 19340 5296
rect 13403 5256 19340 5284
rect 13403 5253 13415 5256
rect 13357 5247 13415 5253
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 14366 5216 14372 5228
rect 13679 5188 14372 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 19429 5219 19487 5225
rect 19429 5185 19441 5219
rect 19475 5216 19487 5219
rect 56413 5219 56471 5225
rect 19475 5188 19932 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 19904 5089 19932 5188
rect 56413 5185 56425 5219
rect 56459 5216 56471 5219
rect 58342 5216 58348 5228
rect 56459 5188 58348 5216
rect 56459 5185 56471 5188
rect 56413 5179 56471 5185
rect 58342 5176 58348 5188
rect 58400 5176 58406 5228
rect 20162 5108 20168 5160
rect 20220 5148 20226 5160
rect 20349 5151 20407 5157
rect 20349 5148 20361 5151
rect 20220 5120 20361 5148
rect 20220 5108 20226 5120
rect 20349 5117 20361 5120
rect 20395 5117 20407 5151
rect 20349 5111 20407 5117
rect 20438 5108 20444 5160
rect 20496 5148 20502 5160
rect 20496 5120 20541 5148
rect 20496 5108 20502 5120
rect 19889 5083 19947 5089
rect 19889 5049 19901 5083
rect 19935 5049 19947 5083
rect 19889 5043 19947 5049
rect 20254 5012 20260 5024
rect 11900 4984 20260 5012
rect 20254 4972 20260 4984
rect 20312 4972 20318 5024
rect 22741 5015 22799 5021
rect 22741 4981 22753 5015
rect 22787 5012 22799 5015
rect 22830 5012 22836 5024
rect 22787 4984 22836 5012
rect 22787 4981 22799 4984
rect 22741 4975 22799 4981
rect 22830 4972 22836 4984
rect 22888 4972 22894 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 3053 4811 3111 4817
rect 3053 4808 3065 4811
rect 2924 4780 3065 4808
rect 2924 4768 2930 4780
rect 3053 4777 3065 4780
rect 3099 4808 3111 4811
rect 3970 4808 3976 4820
rect 3099 4780 3976 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 16574 4768 16580 4820
rect 16632 4808 16638 4820
rect 19705 4811 19763 4817
rect 19705 4808 19717 4811
rect 16632 4780 19717 4808
rect 16632 4768 16638 4780
rect 19705 4777 19717 4780
rect 19751 4808 19763 4811
rect 20162 4808 20168 4820
rect 19751 4780 20168 4808
rect 19751 4777 19763 4780
rect 19705 4771 19763 4777
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 56502 4808 56508 4820
rect 56463 4780 56508 4808
rect 56502 4768 56508 4780
rect 56560 4768 56566 4820
rect 57514 4808 57520 4820
rect 57475 4780 57520 4808
rect 57514 4768 57520 4780
rect 57572 4768 57578 4820
rect 58158 4808 58164 4820
rect 58119 4780 58164 4808
rect 58158 4768 58164 4780
rect 58216 4768 58222 4820
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 2498 4604 2504 4616
rect 1903 4576 2504 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 57057 4607 57115 4613
rect 57057 4573 57069 4607
rect 57103 4604 57115 4607
rect 57698 4604 57704 4616
rect 57103 4576 57704 4604
rect 57103 4573 57115 4576
rect 57057 4567 57115 4573
rect 57698 4564 57704 4576
rect 57756 4564 57762 4616
rect 58342 4604 58348 4616
rect 58303 4576 58348 4604
rect 58342 4564 58348 4576
rect 58400 4564 58406 4616
rect 55953 4539 56011 4545
rect 55953 4505 55965 4539
rect 55999 4536 56011 4539
rect 58360 4536 58388 4564
rect 55999 4508 58388 4536
rect 55999 4505 56011 4508
rect 55953 4499 56011 4505
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4428 1734 4480
rect 20162 4428 20168 4480
rect 20220 4468 20226 4480
rect 20257 4471 20315 4477
rect 20257 4468 20269 4471
rect 20220 4440 20269 4468
rect 20220 4428 20226 4440
rect 20257 4437 20269 4440
rect 20303 4437 20315 4471
rect 20257 4431 20315 4437
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21358 4468 21364 4480
rect 21131 4440 21364 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21358 4428 21364 4440
rect 21416 4428 21422 4480
rect 22741 4471 22799 4477
rect 22741 4437 22753 4471
rect 22787 4468 22799 4471
rect 23014 4468 23020 4480
rect 22787 4440 23020 4468
rect 22787 4437 22799 4440
rect 22741 4431 22799 4437
rect 23014 4428 23020 4440
rect 23072 4428 23078 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2593 4267 2651 4273
rect 2593 4264 2605 4267
rect 2464 4236 2605 4264
rect 2464 4224 2470 4236
rect 2593 4233 2605 4236
rect 2639 4233 2651 4267
rect 2593 4227 2651 4233
rect 2961 4267 3019 4273
rect 2961 4233 2973 4267
rect 3007 4233 3019 4267
rect 19242 4264 19248 4276
rect 19203 4236 19248 4264
rect 2961 4227 3019 4233
rect 2608 4128 2636 4227
rect 2976 4128 3004 4227
rect 19242 4224 19248 4236
rect 19300 4264 19306 4276
rect 20073 4267 20131 4273
rect 20073 4264 20085 4267
rect 19300 4236 20085 4264
rect 19300 4224 19306 4236
rect 20073 4233 20085 4236
rect 20119 4233 20131 4267
rect 23198 4264 23204 4276
rect 20073 4227 20131 4233
rect 21376 4236 23204 4264
rect 3326 4156 3332 4208
rect 3384 4196 3390 4208
rect 3384 4168 3556 4196
rect 3384 4156 3390 4168
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 2608 4100 2912 4128
rect 2976 4100 3433 4128
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 2682 4060 2688 4072
rect 2547 4032 2688 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 2424 3992 2452 4023
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 2884 4060 2912 4100
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 3528 4128 3556 4168
rect 4632 4168 6684 4196
rect 4632 4128 4660 4168
rect 3528 4100 4660 4128
rect 3421 4091 3479 4097
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 4764 4100 6561 4128
rect 4764 4088 4770 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6656 4128 6684 4168
rect 6656 4100 8064 4128
rect 6549 4091 6607 4097
rect 4157 4063 4215 4069
rect 4157 4060 4169 4063
rect 2884 4032 4169 4060
rect 4157 4029 4169 4032
rect 4203 4060 4215 4063
rect 7926 4060 7932 4072
rect 4203 4032 7932 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8036 4060 8064 4100
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 19426 4128 19432 4140
rect 9916 4100 19432 4128
rect 9916 4088 9922 4100
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 21376 4137 21404 4236
rect 23198 4224 23204 4236
rect 23256 4224 23262 4276
rect 22462 4156 22468 4208
rect 22520 4196 22526 4208
rect 22925 4199 22983 4205
rect 22925 4196 22937 4199
rect 22520 4168 22937 4196
rect 22520 4156 22526 4168
rect 22925 4165 22937 4168
rect 22971 4165 22983 4199
rect 22925 4159 22983 4165
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 19576 4100 20177 4128
rect 19576 4088 19582 4100
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 21361 4131 21419 4137
rect 21361 4128 21373 4131
rect 20165 4091 20223 4097
rect 20364 4100 21373 4128
rect 20364 4072 20392 4100
rect 21361 4097 21373 4100
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 24118 4088 24124 4140
rect 24176 4128 24182 4140
rect 30006 4128 30012 4140
rect 24176 4100 30012 4128
rect 24176 4088 24182 4100
rect 30006 4088 30012 4100
rect 30064 4088 30070 4140
rect 55674 4088 55680 4140
rect 55732 4128 55738 4140
rect 55769 4131 55827 4137
rect 55769 4128 55781 4131
rect 55732 4100 55781 4128
rect 55732 4088 55738 4100
rect 55769 4097 55781 4100
rect 55815 4097 55827 4131
rect 55769 4091 55827 4097
rect 56873 4131 56931 4137
rect 56873 4097 56885 4131
rect 56919 4128 56931 4131
rect 57517 4131 57575 4137
rect 57517 4128 57529 4131
rect 56919 4100 57529 4128
rect 56919 4097 56931 4100
rect 56873 4091 56931 4097
rect 57517 4097 57529 4100
rect 57563 4128 57575 4131
rect 57790 4128 57796 4140
rect 57563 4100 57796 4128
rect 57563 4097 57575 4100
rect 57517 4091 57575 4097
rect 57790 4088 57796 4100
rect 57848 4088 57854 4140
rect 58253 4131 58311 4137
rect 58253 4097 58265 4131
rect 58299 4097 58311 4131
rect 58253 4091 58311 4097
rect 16390 4060 16396 4072
rect 8036 4032 16396 4060
rect 16390 4020 16396 4032
rect 16448 4060 16454 4072
rect 16448 4032 20300 4060
rect 16448 4020 16454 4032
rect 2866 3992 2872 4004
rect 2424 3964 2872 3992
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3418 3952 3424 4004
rect 3476 3992 3482 4004
rect 11146 3992 11152 4004
rect 3476 3964 11152 3992
rect 3476 3952 3482 3964
rect 11146 3952 11152 3964
rect 11204 3952 11210 4004
rect 16758 3952 16764 4004
rect 16816 3992 16822 4004
rect 18141 3995 18199 4001
rect 16816 3964 18092 3992
rect 16816 3952 16822 3964
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 2406 3924 2412 3936
rect 1811 3896 2412 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 3602 3924 3608 3936
rect 3563 3896 3608 3924
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 4028 3896 4629 3924
rect 4028 3884 4034 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 7282 3924 7288 3936
rect 6779 3896 7288 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 7282 3884 7288 3896
rect 7340 3924 7346 3936
rect 11054 3924 11060 3936
rect 7340 3896 11060 3924
rect 7340 3884 7346 3896
rect 11054 3884 11060 3896
rect 11112 3924 11118 3936
rect 11974 3924 11980 3936
rect 11112 3896 11980 3924
rect 11112 3884 11118 3896
rect 11974 3884 11980 3896
rect 12032 3884 12038 3936
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 17770 3924 17776 3936
rect 17635 3896 17776 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18064 3924 18092 3964
rect 18141 3961 18153 3995
rect 18187 3992 18199 3995
rect 20070 3992 20076 4004
rect 18187 3964 20076 3992
rect 18187 3961 18199 3964
rect 18141 3955 18199 3961
rect 20070 3952 20076 3964
rect 20128 3952 20134 4004
rect 20272 3992 20300 4032
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 20404 4032 20497 4060
rect 20404 4020 20410 4032
rect 20622 4020 20628 4072
rect 20680 4060 20686 4072
rect 21085 4063 21143 4069
rect 21085 4060 21097 4063
rect 20680 4032 21097 4060
rect 20680 4020 20686 4032
rect 21085 4029 21097 4032
rect 21131 4029 21143 4063
rect 21085 4023 21143 4029
rect 23017 4063 23075 4069
rect 23017 4029 23029 4063
rect 23063 4029 23075 4063
rect 23198 4060 23204 4072
rect 23159 4032 23204 4060
rect 23017 4023 23075 4029
rect 22005 3995 22063 4001
rect 22005 3992 22017 3995
rect 20272 3964 22017 3992
rect 22005 3961 22017 3964
rect 22051 3992 22063 3995
rect 23032 3992 23060 4023
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 23750 4020 23756 4072
rect 23808 4060 23814 4072
rect 28902 4060 28908 4072
rect 23808 4032 28908 4060
rect 23808 4020 23814 4032
rect 28902 4020 28908 4032
rect 28960 4020 28966 4072
rect 56134 4020 56140 4072
rect 56192 4060 56198 4072
rect 58268 4060 58296 4091
rect 56192 4032 58296 4060
rect 56192 4020 56198 4032
rect 22051 3964 23060 3992
rect 22051 3961 22063 3964
rect 22005 3955 22063 3961
rect 53374 3952 53380 4004
rect 53432 3992 53438 4004
rect 57333 3995 57391 4001
rect 57333 3992 57345 3995
rect 53432 3964 57345 3992
rect 53432 3952 53438 3964
rect 57333 3961 57345 3964
rect 57379 3961 57391 3995
rect 57333 3955 57391 3961
rect 18601 3927 18659 3933
rect 18601 3924 18613 3927
rect 18064 3896 18613 3924
rect 18601 3893 18613 3896
rect 18647 3924 18659 3927
rect 19518 3924 19524 3936
rect 18647 3896 19524 3924
rect 18647 3893 18659 3896
rect 18601 3887 18659 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19702 3924 19708 3936
rect 19663 3896 19708 3924
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 22094 3884 22100 3936
rect 22152 3924 22158 3936
rect 22557 3927 22615 3933
rect 22557 3924 22569 3927
rect 22152 3896 22569 3924
rect 22152 3884 22158 3896
rect 22557 3893 22569 3896
rect 22603 3893 22615 3927
rect 22557 3887 22615 3893
rect 55309 3927 55367 3933
rect 55309 3893 55321 3927
rect 55355 3924 55367 3927
rect 56502 3924 56508 3936
rect 55355 3896 56508 3924
rect 55355 3893 55367 3896
rect 55309 3887 55367 3893
rect 56502 3884 56508 3896
rect 56560 3884 56566 3936
rect 58069 3927 58127 3933
rect 58069 3893 58081 3927
rect 58115 3924 58127 3927
rect 58158 3924 58164 3936
rect 58115 3896 58164 3924
rect 58115 3893 58127 3896
rect 58069 3887 58127 3893
rect 58158 3884 58164 3896
rect 58216 3884 58222 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 2746 3692 4997 3720
rect 2498 3612 2504 3664
rect 2556 3652 2562 3664
rect 2746 3652 2774 3692
rect 4985 3689 4997 3692
rect 5031 3689 5043 3723
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 4985 3683 5043 3689
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 8938 3680 8944 3732
rect 8996 3720 9002 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 8996 3692 11345 3720
rect 8996 3680 9002 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 11333 3683 11391 3689
rect 2556 3624 2774 3652
rect 4157 3655 4215 3661
rect 2556 3612 2562 3624
rect 4157 3621 4169 3655
rect 4203 3621 4215 3655
rect 4157 3615 4215 3621
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 2866 3584 2872 3596
rect 2455 3556 2872 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 4172 3584 4200 3615
rect 6457 3587 6515 3593
rect 6457 3584 6469 3587
rect 4172 3556 6469 3584
rect 6457 3553 6469 3556
rect 6503 3553 6515 3587
rect 9858 3584 9864 3596
rect 9819 3556 9864 3584
rect 6457 3547 6515 3553
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 11348 3584 11376 3683
rect 11974 3680 11980 3732
rect 12032 3720 12038 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 12032 3692 13645 3720
rect 12032 3680 12038 3692
rect 13633 3689 13645 3692
rect 13679 3720 13691 3723
rect 14274 3720 14280 3732
rect 13679 3692 14280 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 16390 3720 16396 3732
rect 16351 3692 16396 3720
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 40862 3720 40868 3732
rect 16500 3692 21496 3720
rect 40823 3692 40868 3720
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 16500 3652 16528 3692
rect 13780 3624 16528 3652
rect 13780 3612 13786 3624
rect 20073 3587 20131 3593
rect 11348 3556 19840 3584
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 2590 3516 2596 3528
rect 2547 3488 2596 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3516 6791 3519
rect 6914 3516 6920 3528
rect 6779 3488 6920 3516
rect 6779 3485 6791 3488
rect 6733 3479 6791 3485
rect 6914 3476 6920 3488
rect 6972 3516 6978 3528
rect 9582 3516 9588 3528
rect 6972 3488 9588 3516
rect 6972 3476 6978 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14332 3488 14381 3516
rect 14332 3476 14338 3488
rect 14369 3485 14381 3488
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3516 14795 3519
rect 18141 3519 18199 3525
rect 14783 3488 15516 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 1578 3408 1584 3460
rect 1636 3448 1642 3460
rect 5074 3448 5080 3460
rect 1636 3420 5080 3448
rect 1636 3408 1642 3420
rect 5074 3408 5080 3420
rect 5132 3408 5138 3460
rect 6546 3448 6552 3460
rect 6026 3420 6552 3448
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 6822 3408 6828 3460
rect 6880 3448 6886 3460
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 6880 3420 7757 3448
rect 6880 3408 6886 3420
rect 7745 3417 7757 3420
rect 7791 3417 7803 3451
rect 7745 3411 7803 3417
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 10318 3448 10324 3460
rect 9088 3420 10324 3448
rect 9088 3408 9094 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 14752 3448 14780 3479
rect 13688 3420 14780 3448
rect 13688 3408 13694 3420
rect 1765 3383 1823 3389
rect 1765 3349 1777 3383
rect 1811 3380 1823 3383
rect 1946 3380 1952 3392
rect 1811 3352 1952 3380
rect 1811 3349 1823 3352
rect 1765 3343 1823 3349
rect 1946 3340 1952 3352
rect 2004 3380 2010 3392
rect 2222 3380 2228 3392
rect 2004 3352 2228 3380
rect 2004 3340 2010 3352
rect 2222 3340 2228 3352
rect 2280 3380 2286 3392
rect 2593 3383 2651 3389
rect 2593 3380 2605 3383
rect 2280 3352 2605 3380
rect 2280 3340 2286 3352
rect 2593 3349 2605 3352
rect 2639 3349 2651 3383
rect 2958 3380 2964 3392
rect 2919 3352 2964 3380
rect 2593 3343 2651 3349
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 7006 3380 7012 3392
rect 4488 3352 7012 3380
rect 4488 3340 4494 3352
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 8570 3380 8576 3392
rect 8531 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 14734 3340 14740 3392
rect 14792 3380 14798 3392
rect 15197 3383 15255 3389
rect 15197 3380 15209 3383
rect 14792 3352 15209 3380
rect 14792 3340 14798 3352
rect 15197 3349 15209 3352
rect 15243 3349 15255 3383
rect 15488 3380 15516 3488
rect 18141 3485 18153 3519
rect 18187 3516 18199 3519
rect 18598 3516 18604 3528
rect 18187 3488 18604 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3516 18935 3519
rect 19702 3516 19708 3528
rect 18923 3488 19708 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 19702 3476 19708 3488
rect 19760 3476 19766 3528
rect 19812 3516 19840 3556
rect 20073 3553 20085 3587
rect 20119 3584 20131 3587
rect 20346 3584 20352 3596
rect 20119 3556 20352 3584
rect 20119 3553 20131 3556
rect 20073 3547 20131 3553
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 21468 3593 21496 3692
rect 40862 3680 40868 3692
rect 40920 3680 40926 3732
rect 48685 3723 48743 3729
rect 48685 3689 48697 3723
rect 48731 3720 48743 3723
rect 55950 3720 55956 3732
rect 48731 3692 55956 3720
rect 48731 3689 48743 3692
rect 48685 3683 48743 3689
rect 21453 3587 21511 3593
rect 21453 3553 21465 3587
rect 21499 3584 21511 3587
rect 23017 3587 23075 3593
rect 23017 3584 23029 3587
rect 21499 3556 23029 3584
rect 21499 3553 21511 3556
rect 21453 3547 21511 3553
rect 23017 3553 23029 3556
rect 23063 3553 23075 3587
rect 23017 3547 23075 3553
rect 23198 3544 23204 3596
rect 23256 3584 23262 3596
rect 23753 3587 23811 3593
rect 23753 3584 23765 3587
rect 23256 3556 23765 3584
rect 23256 3544 23262 3556
rect 23753 3553 23765 3556
rect 23799 3553 23811 3587
rect 23753 3547 23811 3553
rect 20162 3516 20168 3528
rect 19812 3488 20168 3516
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 40405 3519 40463 3525
rect 22152 3488 22197 3516
rect 22152 3476 22158 3488
rect 40405 3485 40417 3519
rect 40451 3516 40463 3519
rect 40862 3516 40868 3528
rect 40451 3488 40868 3516
rect 40451 3485 40463 3488
rect 40405 3479 40463 3485
rect 40862 3476 40868 3488
rect 40920 3476 40926 3528
rect 48133 3519 48191 3525
rect 48133 3485 48145 3519
rect 48179 3516 48191 3519
rect 48700 3516 48728 3683
rect 55950 3680 55956 3692
rect 56008 3680 56014 3732
rect 53742 3612 53748 3664
rect 53800 3652 53806 3664
rect 57330 3652 57336 3664
rect 53800 3624 57336 3652
rect 53800 3612 53806 3624
rect 57330 3612 57336 3624
rect 57388 3612 57394 3664
rect 54021 3587 54079 3593
rect 54021 3553 54033 3587
rect 54067 3584 54079 3587
rect 55306 3584 55312 3596
rect 54067 3556 55312 3584
rect 54067 3553 54079 3556
rect 54021 3547 54079 3553
rect 55306 3544 55312 3556
rect 55364 3544 55370 3596
rect 55582 3544 55588 3596
rect 55640 3584 55646 3596
rect 55640 3556 56364 3584
rect 55640 3544 55646 3556
rect 54662 3516 54668 3528
rect 48179 3488 48728 3516
rect 54623 3488 54668 3516
rect 48179 3485 48191 3488
rect 48133 3479 48191 3485
rect 54662 3476 54668 3488
rect 54720 3476 54726 3528
rect 55674 3516 55680 3528
rect 55635 3488 55680 3516
rect 55674 3476 55680 3488
rect 55732 3476 55738 3528
rect 56336 3525 56364 3556
rect 56321 3519 56379 3525
rect 56321 3485 56333 3519
rect 56367 3485 56379 3519
rect 56321 3479 56379 3485
rect 56594 3476 56600 3528
rect 56652 3516 56658 3528
rect 56965 3519 57023 3525
rect 56965 3516 56977 3519
rect 56652 3488 56977 3516
rect 56652 3476 56658 3488
rect 56965 3485 56977 3488
rect 57011 3485 57023 3519
rect 57422 3516 57428 3528
rect 57383 3488 57428 3516
rect 56965 3479 57023 3485
rect 57422 3476 57428 3488
rect 57480 3476 57486 3528
rect 58250 3516 58256 3528
rect 58211 3488 58256 3516
rect 58250 3476 58256 3488
rect 58308 3476 58314 3528
rect 17586 3448 17592 3460
rect 17434 3420 17592 3448
rect 17512 3380 17540 3420
rect 17586 3408 17592 3420
rect 17644 3408 17650 3460
rect 17865 3451 17923 3457
rect 17865 3417 17877 3451
rect 17911 3448 17923 3451
rect 17911 3420 21956 3448
rect 17911 3417 17923 3420
rect 17865 3411 17923 3417
rect 15488 3352 17540 3380
rect 15197 3343 15255 3349
rect 18322 3340 18328 3392
rect 18380 3380 18386 3392
rect 18693 3383 18751 3389
rect 18693 3380 18705 3383
rect 18380 3352 18705 3380
rect 18380 3340 18386 3352
rect 18693 3349 18705 3352
rect 18739 3349 18751 3383
rect 18693 3343 18751 3349
rect 19978 3340 19984 3392
rect 20036 3380 20042 3392
rect 20257 3383 20315 3389
rect 20257 3380 20269 3383
rect 20036 3352 20269 3380
rect 20036 3340 20042 3352
rect 20257 3349 20269 3352
rect 20303 3380 20315 3383
rect 20438 3380 20444 3392
rect 20303 3352 20444 3380
rect 20303 3349 20315 3352
rect 20257 3343 20315 3349
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 20530 3340 20536 3392
rect 20588 3380 20594 3392
rect 21928 3389 21956 3420
rect 23198 3408 23204 3460
rect 23256 3448 23262 3460
rect 23937 3451 23995 3457
rect 23937 3448 23949 3451
rect 23256 3420 23949 3448
rect 23256 3408 23262 3420
rect 23937 3417 23949 3420
rect 23983 3417 23995 3451
rect 23937 3411 23995 3417
rect 20625 3383 20683 3389
rect 20625 3380 20637 3383
rect 20588 3352 20637 3380
rect 20588 3340 20594 3352
rect 20625 3349 20637 3352
rect 20671 3349 20683 3383
rect 20625 3343 20683 3349
rect 21913 3383 21971 3389
rect 21913 3349 21925 3383
rect 21959 3349 21971 3383
rect 21913 3343 21971 3349
rect 22370 3340 22376 3392
rect 22428 3380 22434 3392
rect 22557 3383 22615 3389
rect 22557 3380 22569 3383
rect 22428 3352 22569 3380
rect 22428 3340 22434 3352
rect 22557 3349 22569 3352
rect 22603 3349 22615 3383
rect 22557 3343 22615 3349
rect 22738 3340 22744 3392
rect 22796 3380 22802 3392
rect 22925 3383 22983 3389
rect 22925 3380 22937 3383
rect 22796 3352 22937 3380
rect 22796 3340 22802 3352
rect 22925 3349 22937 3352
rect 22971 3349 22983 3383
rect 22925 3343 22983 3349
rect 40221 3383 40279 3389
rect 40221 3349 40233 3383
rect 40267 3380 40279 3383
rect 40310 3380 40316 3392
rect 40267 3352 40316 3380
rect 40267 3349 40279 3352
rect 40221 3343 40279 3349
rect 40310 3340 40316 3352
rect 40368 3340 40374 3392
rect 47949 3383 48007 3389
rect 47949 3349 47961 3383
rect 47995 3380 48007 3383
rect 48038 3380 48044 3392
rect 47995 3352 48044 3380
rect 47995 3349 48007 3352
rect 47949 3343 48007 3349
rect 48038 3340 48044 3352
rect 48096 3340 48102 3392
rect 54478 3380 54484 3392
rect 54439 3352 54484 3380
rect 54478 3340 54484 3352
rect 54536 3340 54542 3392
rect 55490 3380 55496 3392
rect 55451 3352 55496 3380
rect 55490 3340 55496 3352
rect 55548 3340 55554 3392
rect 56134 3380 56140 3392
rect 56095 3352 56140 3380
rect 56134 3340 56140 3352
rect 56192 3340 56198 3392
rect 56778 3380 56784 3392
rect 56739 3352 56784 3380
rect 56778 3340 56784 3352
rect 56836 3340 56842 3392
rect 57609 3383 57667 3389
rect 57609 3349 57621 3383
rect 57655 3380 57667 3383
rect 57974 3380 57980 3392
rect 57655 3352 57980 3380
rect 57655 3349 57667 3352
rect 57609 3343 57667 3349
rect 57974 3340 57980 3352
rect 58032 3340 58038 3392
rect 58066 3340 58072 3392
rect 58124 3380 58130 3392
rect 58124 3352 58169 3380
rect 58124 3340 58130 3352
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1762 3176 1768 3188
rect 1723 3148 1768 3176
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 2590 3136 2596 3188
rect 2648 3136 2654 3188
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3970 3176 3976 3188
rect 3007 3148 3976 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 12621 3179 12679 3185
rect 12621 3176 12633 3179
rect 5132 3148 12633 3176
rect 5132 3136 5138 3148
rect 12621 3145 12633 3148
rect 12667 3176 12679 3179
rect 13722 3176 13728 3188
rect 12667 3148 13728 3176
rect 12667 3145 12679 3148
rect 12621 3139 12679 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 14108 3148 22201 3176
rect 1780 3040 1808 3136
rect 2608 3108 2636 3136
rect 4430 3108 4436 3120
rect 2608 3080 4436 3108
rect 4430 3068 4436 3080
rect 4488 3068 4494 3120
rect 6638 3108 6644 3120
rect 5290 3080 6644 3108
rect 6638 3068 6644 3080
rect 6696 3108 6702 3120
rect 6733 3111 6791 3117
rect 6733 3108 6745 3111
rect 6696 3080 6745 3108
rect 6696 3068 6702 3080
rect 6733 3077 6745 3080
rect 6779 3077 6791 3111
rect 6733 3071 6791 3077
rect 9030 3068 9036 3120
rect 9088 3068 9094 3120
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 9640 3080 9812 3108
rect 9640 3068 9646 3080
rect 2590 3040 2596 3052
rect 1780 3012 2596 3040
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 2958 3000 2964 3052
rect 3016 3040 3022 3052
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 3016 3012 3433 3040
rect 3016 3000 3022 3012
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3602 3000 3608 3052
rect 3660 3040 3666 3052
rect 5997 3043 6055 3049
rect 3660 3012 4568 3040
rect 3660 3000 3666 3012
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2941 2467 2975
rect 2409 2935 2467 2941
rect 2424 2904 2452 2935
rect 2682 2932 2688 2984
rect 2740 2972 2746 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 2740 2944 4261 2972
rect 2740 2932 2746 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4540 2972 4568 3012
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 6914 3040 6920 3052
rect 6043 3012 6920 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7282 3040 7288 3052
rect 7055 3012 7288 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 9784 3049 9812 3080
rect 13630 3068 13636 3120
rect 13688 3068 13694 3120
rect 14108 3117 14136 3148
rect 22189 3145 22201 3148
rect 22235 3145 22247 3179
rect 23198 3176 23204 3188
rect 23159 3148 23204 3176
rect 22189 3139 22247 3145
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 27246 3176 27252 3188
rect 27207 3148 27252 3176
rect 27246 3136 27252 3148
rect 27304 3136 27310 3188
rect 28813 3179 28871 3185
rect 28813 3145 28825 3179
rect 28859 3176 28871 3179
rect 28902 3176 28908 3188
rect 28859 3148 28908 3176
rect 28859 3145 28871 3148
rect 28813 3139 28871 3145
rect 28902 3136 28908 3148
rect 28960 3136 28966 3188
rect 29917 3179 29975 3185
rect 29917 3145 29929 3179
rect 29963 3176 29975 3179
rect 30006 3176 30012 3188
rect 29963 3148 30012 3176
rect 29963 3145 29975 3148
rect 29917 3139 29975 3145
rect 30006 3136 30012 3148
rect 30064 3136 30070 3188
rect 30926 3176 30932 3188
rect 30887 3148 30932 3176
rect 30926 3136 30932 3148
rect 30984 3136 30990 3188
rect 33229 3179 33287 3185
rect 33229 3145 33241 3179
rect 33275 3176 33287 3179
rect 33318 3176 33324 3188
rect 33275 3148 33324 3176
rect 33275 3145 33287 3148
rect 33229 3139 33287 3145
rect 33318 3136 33324 3148
rect 33376 3136 33382 3188
rect 43622 3136 43628 3188
rect 43680 3176 43686 3188
rect 43809 3179 43867 3185
rect 43809 3176 43821 3179
rect 43680 3148 43821 3176
rect 43680 3136 43686 3148
rect 43809 3145 43821 3148
rect 43855 3176 43867 3179
rect 44358 3176 44364 3188
rect 43855 3148 44364 3176
rect 43855 3145 43867 3148
rect 43809 3139 43867 3145
rect 44358 3136 44364 3148
rect 44416 3136 44422 3188
rect 44818 3176 44824 3188
rect 44779 3148 44824 3176
rect 44818 3136 44824 3148
rect 44876 3136 44882 3188
rect 45830 3176 45836 3188
rect 45791 3148 45836 3176
rect 45830 3136 45836 3148
rect 45888 3136 45894 3188
rect 51442 3176 51448 3188
rect 51403 3148 51448 3176
rect 51442 3136 51448 3148
rect 51500 3136 51506 3188
rect 53742 3176 53748 3188
rect 53703 3148 53748 3176
rect 53742 3136 53748 3148
rect 53800 3136 53806 3188
rect 54662 3136 54668 3188
rect 54720 3176 54726 3188
rect 54757 3179 54815 3185
rect 54757 3176 54769 3179
rect 54720 3148 54769 3176
rect 54720 3136 54726 3148
rect 54757 3145 54769 3148
rect 54803 3145 54815 3179
rect 56686 3176 56692 3188
rect 56647 3148 56692 3176
rect 54757 3139 54815 3145
rect 56686 3136 56692 3148
rect 56744 3136 56750 3188
rect 14093 3111 14151 3117
rect 14093 3077 14105 3111
rect 14139 3077 14151 3111
rect 14093 3071 14151 3077
rect 17586 3068 17592 3120
rect 17644 3068 17650 3120
rect 18322 3108 18328 3120
rect 18283 3080 18328 3108
rect 18322 3068 18328 3080
rect 18380 3068 18386 3120
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 14424 3012 14469 3040
rect 14424 3000 14430 3012
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 19334 3040 19340 3052
rect 18656 3012 18701 3040
rect 19295 3012 19340 3040
rect 18656 3000 18662 3012
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 20530 3040 20536 3052
rect 20491 3012 20536 3040
rect 20530 3000 20536 3012
rect 20588 3000 20594 3052
rect 21082 3000 21088 3052
rect 21140 3040 21146 3052
rect 21358 3040 21364 3052
rect 21140 3012 21364 3040
rect 21140 3000 21146 3012
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 22370 3040 22376 3052
rect 22331 3012 22376 3040
rect 22370 3000 22376 3012
rect 22428 3000 22434 3052
rect 22830 3040 22836 3052
rect 22791 3012 22836 3040
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 23014 3040 23020 3052
rect 22975 3012 23020 3040
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 27264 3040 27292 3136
rect 30282 3068 30288 3120
rect 30340 3108 30346 3120
rect 32306 3108 32312 3120
rect 30340 3080 32312 3108
rect 30340 3068 30346 3080
rect 32306 3068 32312 3080
rect 32364 3068 32370 3120
rect 37734 3068 37740 3120
rect 37792 3108 37798 3120
rect 37921 3111 37979 3117
rect 37921 3108 37933 3111
rect 37792 3080 37933 3108
rect 37792 3068 37798 3080
rect 37921 3077 37933 3080
rect 37967 3108 37979 3111
rect 58066 3108 58072 3120
rect 37967 3080 58072 3108
rect 37967 3077 37979 3080
rect 37921 3071 37979 3077
rect 58066 3068 58072 3080
rect 58124 3068 58130 3120
rect 27801 3043 27859 3049
rect 27801 3040 27813 3043
rect 27264 3012 27813 3040
rect 27801 3009 27813 3012
rect 27847 3009 27859 3043
rect 27801 3003 27859 3009
rect 54297 3043 54355 3049
rect 54297 3009 54309 3043
rect 54343 3040 54355 3043
rect 55950 3040 55956 3052
rect 54343 3012 55956 3040
rect 54343 3009 54355 3012
rect 54297 3003 54355 3009
rect 55950 3000 55956 3012
rect 56008 3000 56014 3052
rect 56042 3000 56048 3052
rect 56100 3040 56106 3052
rect 56100 3012 56145 3040
rect 56100 3000 56106 3012
rect 56502 3000 56508 3052
rect 56560 3040 56566 3052
rect 56873 3043 56931 3049
rect 56873 3040 56885 3043
rect 56560 3012 56885 3040
rect 56560 3000 56566 3012
rect 56873 3009 56885 3012
rect 56919 3009 56931 3043
rect 56873 3003 56931 3009
rect 57330 3000 57336 3052
rect 57388 3040 57394 3052
rect 57517 3043 57575 3049
rect 57517 3040 57529 3043
rect 57388 3012 57529 3040
rect 57388 3000 57394 3012
rect 57517 3009 57529 3012
rect 57563 3009 57575 3043
rect 57517 3003 57575 3009
rect 58253 3043 58311 3049
rect 58253 3009 58265 3043
rect 58299 3040 58311 3043
rect 58434 3040 58440 3052
rect 58299 3012 58440 3040
rect 58299 3009 58311 3012
rect 58253 3003 58311 3009
rect 58434 3000 58440 3012
rect 58492 3000 58498 3052
rect 5721 2975 5779 2981
rect 5721 2972 5733 2975
rect 4540 2944 5733 2972
rect 4249 2935 4307 2941
rect 5721 2941 5733 2944
rect 5767 2941 5779 2975
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 5721 2935 5779 2941
rect 6932 2944 9505 2972
rect 2866 2904 2872 2916
rect 2424 2876 2872 2904
rect 2866 2864 2872 2876
rect 2924 2864 2930 2916
rect 6932 2904 6960 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 16301 2975 16359 2981
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 18874 2972 18880 2984
rect 16347 2944 18880 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 18874 2932 18880 2944
rect 18932 2972 18938 2984
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 18932 2944 19073 2972
rect 18932 2932 18938 2944
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 38654 2972 38660 2984
rect 38567 2944 38660 2972
rect 19061 2935 19119 2941
rect 38654 2932 38660 2944
rect 38712 2972 38718 2984
rect 56134 2972 56140 2984
rect 38712 2944 56140 2972
rect 38712 2932 38718 2944
rect 56134 2932 56140 2944
rect 56192 2932 56198 2984
rect 6564 2876 6960 2904
rect 3605 2839 3663 2845
rect 3605 2805 3617 2839
rect 3651 2836 3663 2839
rect 6564 2836 6592 2876
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 8021 2907 8079 2913
rect 8021 2904 8033 2907
rect 7064 2876 8033 2904
rect 7064 2864 7070 2876
rect 8021 2873 8033 2876
rect 8067 2873 8079 2907
rect 8021 2867 8079 2873
rect 15749 2907 15807 2913
rect 15749 2873 15761 2907
rect 15795 2904 15807 2907
rect 16666 2904 16672 2916
rect 15795 2876 16672 2904
rect 15795 2873 15807 2876
rect 15749 2867 15807 2873
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 16758 2864 16764 2916
rect 16816 2904 16822 2916
rect 16853 2907 16911 2913
rect 16853 2904 16865 2907
rect 16816 2876 16865 2904
rect 16816 2864 16822 2876
rect 16853 2873 16865 2876
rect 16899 2873 16911 2907
rect 16853 2867 16911 2873
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 20349 2907 20407 2913
rect 20349 2904 20361 2907
rect 19484 2876 20361 2904
rect 19484 2864 19490 2876
rect 20349 2873 20361 2876
rect 20395 2873 20407 2907
rect 20349 2867 20407 2873
rect 20438 2864 20444 2916
rect 20496 2904 20502 2916
rect 21177 2907 21235 2913
rect 21177 2904 21189 2907
rect 20496 2876 21189 2904
rect 20496 2864 20502 2876
rect 21177 2873 21189 2876
rect 21223 2873 21235 2907
rect 21177 2867 21235 2873
rect 39206 2864 39212 2916
rect 39264 2904 39270 2916
rect 39393 2907 39451 2913
rect 39393 2904 39405 2907
rect 39264 2876 39405 2904
rect 39264 2864 39270 2876
rect 39393 2873 39405 2876
rect 39439 2904 39451 2907
rect 58069 2907 58127 2913
rect 58069 2904 58081 2907
rect 39439 2876 58081 2904
rect 39439 2873 39451 2876
rect 39393 2867 39451 2873
rect 58069 2873 58081 2876
rect 58115 2873 58127 2907
rect 58069 2867 58127 2873
rect 3651 2808 6592 2836
rect 7561 2839 7619 2845
rect 3651 2805 3663 2808
rect 3605 2799 3663 2805
rect 7561 2805 7573 2839
rect 7607 2836 7619 2839
rect 7834 2836 7840 2848
rect 7607 2808 7840 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 10042 2796 10048 2848
rect 10100 2836 10106 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 10100 2808 10241 2836
rect 10100 2796 10106 2808
rect 10229 2805 10241 2808
rect 10275 2805 10287 2839
rect 11146 2836 11152 2848
rect 11107 2808 11152 2836
rect 10229 2799 10287 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 12250 2836 12256 2848
rect 12115 2808 12256 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 15197 2839 15255 2845
rect 15197 2805 15209 2839
rect 15243 2836 15255 2839
rect 15562 2836 15568 2848
rect 15243 2808 15568 2836
rect 15243 2805 15255 2808
rect 15197 2799 15255 2805
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 23661 2839 23719 2845
rect 23661 2836 23673 2839
rect 23532 2808 23673 2836
rect 23532 2796 23538 2808
rect 23661 2805 23673 2808
rect 23707 2805 23719 2839
rect 24394 2836 24400 2848
rect 24355 2808 24400 2836
rect 23661 2799 23719 2805
rect 24394 2796 24400 2808
rect 24452 2796 24458 2848
rect 25498 2836 25504 2848
rect 25459 2808 25504 2836
rect 25498 2796 25504 2808
rect 25556 2796 25562 2848
rect 27706 2796 27712 2848
rect 27764 2836 27770 2848
rect 27985 2839 28043 2845
rect 27985 2836 27997 2839
rect 27764 2808 27997 2836
rect 27764 2796 27770 2808
rect 27985 2805 27997 2808
rect 28031 2805 28043 2839
rect 35986 2836 35992 2848
rect 35947 2808 35992 2836
rect 27985 2799 28043 2805
rect 35986 2796 35992 2808
rect 36044 2796 36050 2848
rect 50614 2796 50620 2848
rect 50672 2836 50678 2848
rect 50801 2839 50859 2845
rect 50801 2836 50813 2839
rect 50672 2808 50813 2836
rect 50672 2796 50678 2808
rect 50801 2805 50813 2808
rect 50847 2836 50859 2839
rect 54570 2836 54576 2848
rect 50847 2808 54576 2836
rect 50847 2805 50859 2808
rect 50801 2799 50859 2805
rect 54570 2796 54576 2808
rect 54628 2796 54634 2848
rect 55585 2839 55643 2845
rect 55585 2805 55597 2839
rect 55631 2836 55643 2839
rect 56042 2836 56048 2848
rect 55631 2808 56048 2836
rect 55631 2805 55643 2808
rect 55585 2799 55643 2805
rect 56042 2796 56048 2808
rect 56100 2796 56106 2848
rect 56229 2839 56287 2845
rect 56229 2805 56241 2839
rect 56275 2836 56287 2839
rect 57146 2836 57152 2848
rect 56275 2808 57152 2836
rect 56275 2805 56287 2808
rect 56229 2799 56287 2805
rect 57146 2796 57152 2808
rect 57204 2796 57210 2848
rect 57330 2836 57336 2848
rect 57291 2808 57336 2836
rect 57330 2796 57336 2808
rect 57388 2796 57394 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 2593 2635 2651 2641
rect 2593 2601 2605 2635
rect 2639 2632 2651 2635
rect 4706 2632 4712 2644
rect 2639 2604 4712 2632
rect 2639 2601 2651 2604
rect 2593 2595 2651 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 4798 2592 4804 2644
rect 4856 2632 4862 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 4856 2604 10977 2632
rect 4856 2592 4862 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 22462 2632 22468 2644
rect 22423 2604 22468 2632
rect 10965 2595 11023 2601
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 22738 2592 22744 2644
rect 22796 2632 22802 2644
rect 23385 2635 23443 2641
rect 23385 2632 23397 2635
rect 22796 2604 23397 2632
rect 22796 2592 22802 2604
rect 23385 2601 23397 2604
rect 23431 2601 23443 2635
rect 23385 2595 23443 2601
rect 24949 2635 25007 2641
rect 24949 2601 24961 2635
rect 24995 2632 25007 2635
rect 28626 2632 28632 2644
rect 24995 2604 28632 2632
rect 24995 2601 25007 2604
rect 24949 2595 25007 2601
rect 28626 2592 28632 2604
rect 28684 2592 28690 2644
rect 55674 2632 55680 2644
rect 42904 2604 55680 2632
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2774 2564 2780 2576
rect 1995 2536 2780 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 4062 2524 4068 2576
rect 4120 2564 4126 2576
rect 12529 2567 12587 2573
rect 12529 2564 12541 2567
rect 4120 2536 12541 2564
rect 4120 2524 4126 2536
rect 12529 2533 12541 2536
rect 12575 2533 12587 2567
rect 15930 2564 15936 2576
rect 15891 2536 15936 2564
rect 12529 2527 12587 2533
rect 15930 2524 15936 2536
rect 15988 2524 15994 2576
rect 17129 2567 17187 2573
rect 17129 2533 17141 2567
rect 17175 2564 17187 2567
rect 18782 2564 18788 2576
rect 17175 2536 18788 2564
rect 17175 2533 17187 2536
rect 17129 2527 17187 2533
rect 18782 2524 18788 2536
rect 18840 2524 18846 2576
rect 38378 2564 38384 2576
rect 26206 2536 38384 2564
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 2648 2468 6837 2496
rect 2648 2456 2654 2468
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 7926 2496 7932 2508
rect 7887 2468 7932 2496
rect 6825 2459 6883 2465
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 10502 2456 10508 2508
rect 10560 2496 10566 2508
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 10560 2468 14565 2496
rect 10560 2456 10566 2468
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 18141 2499 18199 2505
rect 18141 2465 18153 2499
rect 18187 2496 18199 2499
rect 19150 2496 19156 2508
rect 18187 2468 19156 2496
rect 18187 2465 18199 2468
rect 18141 2459 18199 2465
rect 19150 2456 19156 2468
rect 19208 2456 19214 2508
rect 20070 2496 20076 2508
rect 20031 2468 20076 2496
rect 20070 2456 20076 2468
rect 20128 2456 20134 2508
rect 20254 2456 20260 2508
rect 20312 2496 20318 2508
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 20312 2468 20361 2496
rect 20312 2456 20318 2468
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 20349 2459 20407 2465
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4522 2428 4528 2440
rect 3467 2400 4528 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4522 2388 4528 2400
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 5721 2431 5779 2437
rect 5721 2428 5733 2431
rect 5684 2400 5733 2428
rect 5684 2388 5690 2400
rect 5721 2397 5733 2400
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6972 2400 7021 2428
rect 6972 2388 6978 2400
rect 7009 2397 7021 2400
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 8938 2428 8944 2440
rect 8628 2400 8944 2428
rect 8628 2388 8634 2400
rect 8938 2388 8944 2400
rect 8996 2428 9002 2440
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 8996 2400 9229 2428
rect 8996 2388 9002 2400
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 17770 2388 17776 2440
rect 17828 2428 17834 2440
rect 17865 2431 17923 2437
rect 17865 2428 17877 2431
rect 17828 2400 17877 2428
rect 17828 2388 17834 2400
rect 17865 2397 17877 2400
rect 17911 2397 17923 2431
rect 17865 2391 17923 2397
rect 22281 2431 22339 2437
rect 22281 2397 22293 2431
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 4157 2363 4215 2369
rect 4157 2329 4169 2363
rect 4203 2360 4215 2363
rect 5644 2360 5672 2388
rect 4203 2332 5672 2360
rect 4203 2329 4215 2332
rect 4157 2323 4215 2329
rect 7834 2320 7840 2372
rect 7892 2360 7898 2372
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 7892 2332 8125 2360
rect 7892 2320 7898 2332
rect 8113 2329 8125 2332
rect 8159 2329 8171 2363
rect 8113 2323 8171 2329
rect 10042 2320 10048 2372
rect 10100 2360 10106 2372
rect 10321 2363 10379 2369
rect 10321 2360 10333 2363
rect 10100 2332 10333 2360
rect 10100 2320 10106 2332
rect 10321 2329 10333 2332
rect 10367 2329 10379 2363
rect 10321 2323 10379 2329
rect 11057 2363 11115 2369
rect 11057 2329 11069 2363
rect 11103 2360 11115 2363
rect 11146 2360 11152 2372
rect 11103 2332 11152 2360
rect 11103 2329 11115 2332
rect 11057 2323 11115 2329
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 11885 2363 11943 2369
rect 11885 2329 11897 2363
rect 11931 2360 11943 2363
rect 13354 2360 13360 2372
rect 11931 2332 13360 2360
rect 11931 2329 11943 2332
rect 11885 2323 11943 2329
rect 13354 2320 13360 2332
rect 13412 2360 13418 2372
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 13412 2332 13645 2360
rect 13412 2320 13418 2332
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 13633 2323 13691 2329
rect 14458 2320 14464 2372
rect 14516 2360 14522 2372
rect 14734 2360 14740 2372
rect 14516 2332 14740 2360
rect 14516 2320 14522 2332
rect 14734 2320 14740 2332
rect 14792 2320 14798 2372
rect 15562 2320 15568 2372
rect 15620 2360 15626 2372
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 15620 2332 15761 2360
rect 15620 2320 15626 2332
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 15749 2323 15807 2329
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 16945 2363 17003 2369
rect 16945 2360 16957 2363
rect 16724 2332 16957 2360
rect 16724 2320 16730 2332
rect 16945 2329 16957 2332
rect 16991 2329 17003 2363
rect 16945 2323 17003 2329
rect 19613 2363 19671 2369
rect 19613 2329 19625 2363
rect 19659 2360 19671 2363
rect 22186 2360 22192 2372
rect 19659 2332 22192 2360
rect 19659 2329 19671 2332
rect 19613 2323 19671 2329
rect 22186 2320 22192 2332
rect 22244 2360 22250 2372
rect 22296 2360 22324 2391
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23532 2400 23581 2428
rect 23532 2388 23538 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 26053 2431 26111 2437
rect 26053 2397 26065 2431
rect 26099 2428 26111 2431
rect 26206 2428 26234 2536
rect 38378 2524 38384 2536
rect 38436 2524 38442 2576
rect 27890 2496 27896 2508
rect 27851 2468 27896 2496
rect 27890 2456 27896 2468
rect 27948 2456 27954 2508
rect 35529 2499 35587 2505
rect 35529 2465 35541 2499
rect 35575 2496 35587 2499
rect 35575 2468 42840 2496
rect 35575 2465 35587 2468
rect 35529 2459 35587 2465
rect 28902 2428 28908 2440
rect 26099 2400 26234 2428
rect 28863 2400 28908 2428
rect 26099 2397 26111 2400
rect 26053 2391 26111 2397
rect 28902 2388 28908 2400
rect 28960 2388 28966 2440
rect 30006 2428 30012 2440
rect 29967 2400 30012 2428
rect 30006 2388 30012 2400
rect 30064 2388 30070 2440
rect 30926 2388 30932 2440
rect 30984 2428 30990 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 30984 2400 31125 2428
rect 30984 2388 30990 2400
rect 31113 2397 31125 2400
rect 31159 2397 31171 2431
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 31113 2391 31171 2397
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 33318 2428 33324 2440
rect 33279 2400 33324 2428
rect 33318 2388 33324 2400
rect 33376 2388 33382 2440
rect 34977 2431 35035 2437
rect 34977 2428 34989 2431
rect 34348 2400 34989 2428
rect 22244 2332 22324 2360
rect 22244 2320 22250 2332
rect 24394 2320 24400 2372
rect 24452 2360 24458 2372
rect 24673 2363 24731 2369
rect 24673 2360 24685 2363
rect 24452 2332 24685 2360
rect 24452 2320 24458 2332
rect 24673 2329 24685 2332
rect 24719 2329 24731 2363
rect 24673 2323 24731 2329
rect 25498 2320 25504 2372
rect 25556 2360 25562 2372
rect 25685 2363 25743 2369
rect 25685 2360 25697 2363
rect 25556 2332 25697 2360
rect 25556 2320 25562 2332
rect 25685 2329 25697 2332
rect 25731 2329 25743 2363
rect 25685 2323 25743 2329
rect 27157 2363 27215 2369
rect 27157 2329 27169 2363
rect 27203 2329 27215 2363
rect 27157 2323 27215 2329
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4614 2292 4620 2304
rect 3936 2264 4620 2292
rect 3936 2252 3942 2264
rect 4614 2252 4620 2264
rect 4672 2252 4678 2304
rect 4798 2292 4804 2304
rect 4759 2264 4804 2292
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 5902 2292 5908 2304
rect 5863 2264 5908 2292
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 10226 2292 10232 2304
rect 10187 2264 10232 2292
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 13538 2292 13544 2304
rect 13499 2264 13544 2292
rect 13538 2252 13544 2264
rect 13596 2252 13602 2304
rect 21358 2292 21364 2304
rect 21319 2264 21364 2292
rect 21358 2252 21364 2264
rect 21416 2292 21422 2304
rect 22830 2292 22836 2304
rect 21416 2264 22836 2292
rect 21416 2252 21422 2264
rect 22830 2252 22836 2264
rect 22888 2252 22894 2304
rect 26602 2292 26608 2304
rect 26563 2264 26608 2292
rect 26602 2252 26608 2264
rect 26660 2292 26666 2304
rect 27172 2292 27200 2323
rect 34348 2304 34376 2400
rect 34977 2397 34989 2400
rect 35023 2397 35035 2431
rect 34977 2391 35035 2397
rect 35986 2388 35992 2440
rect 36044 2428 36050 2440
rect 36081 2431 36139 2437
rect 36081 2428 36093 2431
rect 36044 2400 36093 2428
rect 36044 2388 36050 2400
rect 36081 2397 36093 2400
rect 36127 2397 36139 2431
rect 37734 2428 37740 2440
rect 37695 2400 37740 2428
rect 36081 2391 36139 2397
rect 37734 2388 37740 2400
rect 37792 2388 37798 2440
rect 38473 2431 38531 2437
rect 38473 2397 38485 2431
rect 38519 2428 38531 2431
rect 38654 2428 38660 2440
rect 38519 2400 38660 2428
rect 38519 2397 38531 2400
rect 38473 2391 38531 2397
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 39206 2428 39212 2440
rect 39167 2400 39212 2428
rect 39206 2388 39212 2400
rect 39264 2388 39270 2440
rect 40310 2428 40316 2440
rect 40271 2400 40316 2428
rect 40310 2388 40316 2400
rect 40368 2388 40374 2440
rect 41325 2431 41383 2437
rect 41325 2397 41337 2431
rect 41371 2428 41383 2431
rect 41371 2400 41920 2428
rect 41371 2397 41383 2400
rect 41325 2391 41383 2397
rect 36354 2360 36360 2372
rect 36315 2332 36360 2360
rect 36354 2320 36360 2332
rect 36412 2320 36418 2372
rect 41892 2304 41920 2400
rect 42812 2360 42840 2468
rect 42904 2437 42932 2604
rect 55674 2592 55680 2604
rect 55732 2592 55738 2644
rect 56689 2635 56747 2641
rect 56689 2601 56701 2635
rect 56735 2632 56747 2635
rect 57422 2632 57428 2644
rect 56735 2604 57428 2632
rect 56735 2601 56747 2604
rect 56689 2595 56747 2601
rect 57422 2592 57428 2604
rect 57480 2592 57486 2644
rect 57330 2564 57336 2576
rect 51184 2536 57336 2564
rect 47872 2468 51028 2496
rect 42889 2431 42947 2437
rect 42889 2397 42901 2431
rect 42935 2397 42947 2431
rect 43622 2428 43628 2440
rect 43583 2400 43628 2428
rect 42889 2391 42947 2397
rect 43622 2388 43628 2400
rect 43680 2388 43686 2440
rect 44637 2431 44695 2437
rect 44637 2397 44649 2431
rect 44683 2428 44695 2431
rect 44818 2428 44824 2440
rect 44683 2400 44824 2428
rect 44683 2397 44695 2400
rect 44637 2391 44695 2397
rect 44818 2388 44824 2400
rect 44876 2388 44882 2440
rect 45741 2431 45799 2437
rect 45741 2397 45753 2431
rect 45787 2428 45799 2431
rect 45830 2428 45836 2440
rect 45787 2400 45836 2428
rect 45787 2397 45799 2400
rect 45741 2391 45799 2397
rect 45830 2388 45836 2400
rect 45888 2388 45894 2440
rect 46857 2431 46915 2437
rect 46857 2397 46869 2431
rect 46903 2428 46915 2431
rect 47872 2428 47900 2468
rect 48038 2428 48044 2440
rect 46903 2400 47900 2428
rect 47999 2400 48044 2428
rect 46903 2397 46915 2400
rect 46857 2391 46915 2397
rect 48038 2388 48044 2400
rect 48096 2388 48102 2440
rect 49050 2428 49056 2440
rect 49011 2400 49056 2428
rect 49050 2388 49056 2400
rect 49108 2428 49114 2440
rect 49513 2431 49571 2437
rect 49513 2428 49525 2431
rect 49108 2400 49525 2428
rect 49108 2388 49114 2400
rect 49513 2397 49525 2400
rect 49559 2397 49571 2431
rect 50614 2428 50620 2440
rect 50575 2400 50620 2428
rect 49513 2391 49571 2397
rect 50614 2388 50620 2400
rect 50672 2388 50678 2440
rect 51000 2428 51028 2468
rect 51184 2428 51212 2536
rect 57330 2524 57336 2536
rect 57388 2524 57394 2576
rect 56778 2496 56784 2508
rect 55784 2468 56784 2496
rect 51000 2400 51212 2428
rect 51353 2431 51411 2437
rect 51353 2397 51365 2431
rect 51399 2428 51411 2431
rect 51442 2428 51448 2440
rect 51399 2400 51448 2428
rect 51399 2397 51411 2400
rect 51353 2391 51411 2397
rect 51442 2388 51448 2400
rect 51500 2388 51506 2440
rect 52365 2431 52423 2437
rect 52365 2397 52377 2431
rect 52411 2428 52423 2431
rect 53374 2428 53380 2440
rect 52411 2400 53380 2428
rect 52411 2397 52423 2400
rect 52365 2391 52423 2397
rect 53374 2388 53380 2400
rect 53432 2388 53438 2440
rect 53469 2431 53527 2437
rect 53469 2397 53481 2431
rect 53515 2428 53527 2431
rect 54478 2428 54484 2440
rect 53515 2400 54484 2428
rect 53515 2397 53527 2400
rect 53469 2391 53527 2397
rect 54478 2388 54484 2400
rect 54536 2388 54542 2440
rect 54573 2431 54631 2437
rect 54573 2397 54585 2431
rect 54619 2428 54631 2431
rect 55490 2428 55496 2440
rect 54619 2400 55496 2428
rect 54619 2397 54631 2400
rect 54573 2391 54631 2397
rect 55490 2388 55496 2400
rect 55548 2388 55554 2440
rect 55582 2388 55588 2440
rect 55640 2388 55646 2440
rect 55784 2437 55812 2468
rect 56778 2456 56784 2468
rect 56836 2456 56842 2508
rect 55769 2431 55827 2437
rect 55769 2397 55781 2431
rect 55815 2397 55827 2431
rect 55769 2391 55827 2397
rect 55950 2388 55956 2440
rect 56008 2428 56014 2440
rect 56410 2428 56416 2440
rect 56008 2400 56416 2428
rect 56008 2388 56014 2400
rect 56410 2388 56416 2400
rect 56468 2428 56474 2440
rect 56505 2431 56563 2437
rect 56505 2428 56517 2431
rect 56468 2400 56517 2428
rect 56468 2388 56474 2400
rect 56505 2397 56517 2400
rect 56551 2397 56563 2431
rect 57514 2428 57520 2440
rect 57475 2400 57520 2428
rect 56505 2391 56563 2397
rect 57514 2388 57520 2400
rect 57572 2388 57578 2440
rect 57974 2388 57980 2440
rect 58032 2428 58038 2440
rect 58069 2431 58127 2437
rect 58069 2428 58081 2431
rect 58032 2400 58081 2428
rect 58032 2388 58038 2400
rect 58069 2397 58081 2400
rect 58115 2397 58127 2431
rect 58069 2391 58127 2397
rect 55600 2360 55628 2388
rect 42812 2332 55628 2360
rect 55674 2320 55680 2372
rect 55732 2360 55738 2372
rect 58158 2360 58164 2372
rect 55732 2332 58164 2360
rect 55732 2320 55738 2332
rect 58158 2320 58164 2332
rect 58216 2320 58222 2372
rect 26660 2264 27200 2292
rect 26660 2252 26666 2264
rect 28810 2252 28816 2304
rect 28868 2292 28874 2304
rect 29089 2295 29147 2301
rect 29089 2292 29101 2295
rect 28868 2264 29101 2292
rect 28868 2252 28874 2264
rect 29089 2261 29101 2264
rect 29135 2261 29147 2295
rect 29089 2255 29147 2261
rect 29914 2252 29920 2304
rect 29972 2292 29978 2304
rect 30193 2295 30251 2301
rect 30193 2292 30205 2295
rect 29972 2264 30205 2292
rect 29972 2252 29978 2264
rect 30193 2261 30205 2264
rect 30239 2261 30251 2295
rect 30193 2255 30251 2261
rect 31018 2252 31024 2304
rect 31076 2292 31082 2304
rect 31297 2295 31355 2301
rect 31297 2292 31309 2295
rect 31076 2264 31309 2292
rect 31076 2252 31082 2264
rect 31297 2261 31309 2264
rect 31343 2261 31355 2295
rect 31297 2255 31355 2261
rect 32122 2252 32128 2304
rect 32180 2292 32186 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 32180 2264 32505 2292
rect 32180 2252 32186 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 33226 2252 33232 2304
rect 33284 2292 33290 2304
rect 33505 2295 33563 2301
rect 33505 2292 33517 2295
rect 33284 2264 33517 2292
rect 33284 2252 33290 2264
rect 33505 2261 33517 2264
rect 33551 2261 33563 2295
rect 34330 2292 34336 2304
rect 34291 2264 34336 2292
rect 33505 2255 33563 2261
rect 34330 2252 34336 2264
rect 34388 2252 34394 2304
rect 36538 2252 36544 2304
rect 36596 2292 36602 2304
rect 37553 2295 37611 2301
rect 37553 2292 37565 2295
rect 36596 2264 37565 2292
rect 36596 2252 36602 2264
rect 37553 2261 37565 2264
rect 37599 2261 37611 2295
rect 37553 2255 37611 2261
rect 37642 2252 37648 2304
rect 37700 2292 37706 2304
rect 38289 2295 38347 2301
rect 38289 2292 38301 2295
rect 37700 2264 38301 2292
rect 37700 2252 37706 2264
rect 38289 2261 38301 2264
rect 38335 2261 38347 2295
rect 38289 2255 38347 2261
rect 38746 2252 38752 2304
rect 38804 2292 38810 2304
rect 39025 2295 39083 2301
rect 39025 2292 39037 2295
rect 38804 2264 39037 2292
rect 38804 2252 38810 2264
rect 39025 2261 39037 2264
rect 39071 2261 39083 2295
rect 39025 2255 39083 2261
rect 39850 2252 39856 2304
rect 39908 2292 39914 2304
rect 40129 2295 40187 2301
rect 40129 2292 40141 2295
rect 39908 2264 40141 2292
rect 39908 2252 39914 2264
rect 40129 2261 40141 2264
rect 40175 2261 40187 2295
rect 40129 2255 40187 2261
rect 40954 2252 40960 2304
rect 41012 2292 41018 2304
rect 41141 2295 41199 2301
rect 41141 2292 41153 2295
rect 41012 2264 41153 2292
rect 41012 2252 41018 2264
rect 41141 2261 41153 2264
rect 41187 2261 41199 2295
rect 41874 2292 41880 2304
rect 41835 2264 41880 2292
rect 41141 2255 41199 2261
rect 41874 2252 41880 2264
rect 41932 2252 41938 2304
rect 42058 2252 42064 2304
rect 42116 2292 42122 2304
rect 42705 2295 42763 2301
rect 42705 2292 42717 2295
rect 42116 2264 42717 2292
rect 42116 2252 42122 2264
rect 42705 2261 42717 2264
rect 42751 2261 42763 2295
rect 42705 2255 42763 2261
rect 43162 2252 43168 2304
rect 43220 2292 43226 2304
rect 43441 2295 43499 2301
rect 43441 2292 43453 2295
rect 43220 2264 43453 2292
rect 43220 2252 43226 2264
rect 43441 2261 43453 2264
rect 43487 2261 43499 2295
rect 43441 2255 43499 2261
rect 44266 2252 44272 2304
rect 44324 2292 44330 2304
rect 44453 2295 44511 2301
rect 44453 2292 44465 2295
rect 44324 2264 44465 2292
rect 44324 2252 44330 2264
rect 44453 2261 44465 2264
rect 44499 2261 44511 2295
rect 44453 2255 44511 2261
rect 45370 2252 45376 2304
rect 45428 2292 45434 2304
rect 45557 2295 45615 2301
rect 45557 2292 45569 2295
rect 45428 2264 45569 2292
rect 45428 2252 45434 2264
rect 45557 2261 45569 2264
rect 45603 2261 45615 2295
rect 45557 2255 45615 2261
rect 46474 2252 46480 2304
rect 46532 2292 46538 2304
rect 46661 2295 46719 2301
rect 46661 2292 46673 2295
rect 46532 2264 46673 2292
rect 46532 2252 46538 2264
rect 46661 2261 46673 2264
rect 46707 2261 46719 2295
rect 46661 2255 46719 2261
rect 47578 2252 47584 2304
rect 47636 2292 47642 2304
rect 47857 2295 47915 2301
rect 47857 2292 47869 2295
rect 47636 2264 47869 2292
rect 47636 2252 47642 2264
rect 47857 2261 47869 2264
rect 47903 2261 47915 2295
rect 47857 2255 47915 2261
rect 48682 2252 48688 2304
rect 48740 2292 48746 2304
rect 48869 2295 48927 2301
rect 48869 2292 48881 2295
rect 48740 2264 48881 2292
rect 48740 2252 48746 2264
rect 48869 2261 48881 2264
rect 48915 2261 48927 2295
rect 48869 2255 48927 2261
rect 49786 2252 49792 2304
rect 49844 2292 49850 2304
rect 50433 2295 50491 2301
rect 50433 2292 50445 2295
rect 49844 2264 50445 2292
rect 49844 2252 49850 2264
rect 50433 2261 50445 2264
rect 50479 2261 50491 2295
rect 50433 2255 50491 2261
rect 50890 2252 50896 2304
rect 50948 2292 50954 2304
rect 51169 2295 51227 2301
rect 51169 2292 51181 2295
rect 50948 2264 51181 2292
rect 50948 2252 50954 2264
rect 51169 2261 51181 2264
rect 51215 2261 51227 2295
rect 51169 2255 51227 2261
rect 51994 2252 52000 2304
rect 52052 2292 52058 2304
rect 52181 2295 52239 2301
rect 52181 2292 52193 2295
rect 52052 2264 52193 2292
rect 52052 2252 52058 2264
rect 52181 2261 52193 2264
rect 52227 2261 52239 2295
rect 52181 2255 52239 2261
rect 53098 2252 53104 2304
rect 53156 2292 53162 2304
rect 53285 2295 53343 2301
rect 53285 2292 53297 2295
rect 53156 2264 53297 2292
rect 53156 2252 53162 2264
rect 53285 2261 53297 2264
rect 53331 2261 53343 2295
rect 53285 2255 53343 2261
rect 54202 2252 54208 2304
rect 54260 2292 54266 2304
rect 54389 2295 54447 2301
rect 54389 2292 54401 2295
rect 54260 2264 54401 2292
rect 54260 2252 54266 2264
rect 54389 2261 54401 2264
rect 54435 2261 54447 2295
rect 54389 2255 54447 2261
rect 55306 2252 55312 2304
rect 55364 2292 55370 2304
rect 55585 2295 55643 2301
rect 55585 2292 55597 2295
rect 55364 2264 55597 2292
rect 55364 2252 55370 2264
rect 55585 2261 55597 2264
rect 55631 2261 55643 2295
rect 55585 2255 55643 2261
rect 56870 2252 56876 2304
rect 56928 2292 56934 2304
rect 57333 2295 57391 2301
rect 57333 2292 57345 2295
rect 56928 2264 57345 2292
rect 56928 2252 56934 2264
rect 57333 2261 57345 2264
rect 57379 2261 57391 2295
rect 57333 2255 57391 2261
rect 57514 2252 57520 2304
rect 57572 2292 57578 2304
rect 58253 2295 58311 2301
rect 58253 2292 58265 2295
rect 57572 2264 58265 2292
rect 57572 2252 57578 2264
rect 58253 2261 58265 2264
rect 58299 2261 58311 2295
rect 58253 2255 58311 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 4798 2048 4804 2100
rect 4856 2088 4862 2100
rect 23014 2088 23020 2100
rect 4856 2060 23020 2088
rect 4856 2048 4862 2060
rect 23014 2048 23020 2060
rect 23072 2048 23078 2100
rect 36354 2048 36360 2100
rect 36412 2088 36418 2100
rect 55398 2088 55404 2100
rect 36412 2060 55404 2088
rect 36412 2048 36418 2060
rect 55398 2048 55404 2060
rect 55456 2048 55462 2100
rect 3786 1980 3792 2032
rect 3844 2020 3850 2032
rect 13538 2020 13544 2032
rect 3844 1992 13544 2020
rect 3844 1980 3850 1992
rect 13538 1980 13544 1992
rect 13596 1980 13602 2032
rect 41874 1980 41880 2032
rect 41932 2020 41938 2032
rect 51718 2020 51724 2032
rect 41932 1992 51724 2020
rect 41932 1980 41938 1992
rect 51718 1980 51724 1992
rect 51776 1980 51782 2032
rect 3510 1912 3516 1964
rect 3568 1952 3574 1964
rect 10226 1952 10232 1964
rect 3568 1924 10232 1952
rect 3568 1912 3574 1924
rect 10226 1912 10232 1924
rect 10284 1912 10290 1964
rect 5902 1844 5908 1896
rect 5960 1884 5966 1896
rect 21358 1884 21364 1896
rect 5960 1856 21364 1884
rect 5960 1844 5966 1856
rect 21358 1844 21364 1856
rect 21416 1844 21422 1896
rect 2222 1776 2228 1828
rect 2280 1816 2286 1828
rect 9306 1816 9312 1828
rect 2280 1788 9312 1816
rect 2280 1776 2286 1788
rect 9306 1776 9312 1788
rect 9364 1776 9370 1828
<< via1 >>
rect 2228 57808 2280 57860
rect 26240 57808 26292 57860
rect 21640 57740 21692 57792
rect 30288 57740 30340 57792
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 11428 57468 11480 57520
rect 13820 57468 13872 57520
rect 16212 57511 16264 57520
rect 1860 57400 1912 57452
rect 2228 57443 2280 57452
rect 2228 57409 2237 57443
rect 2237 57409 2271 57443
rect 2271 57409 2280 57443
rect 2228 57400 2280 57409
rect 3056 57400 3108 57452
rect 4252 57400 4304 57452
rect 4620 57400 4672 57452
rect 5540 57400 5592 57452
rect 6000 57443 6052 57452
rect 6000 57409 6009 57443
rect 6009 57409 6043 57443
rect 6043 57409 6052 57443
rect 6000 57400 6052 57409
rect 6644 57400 6696 57452
rect 7840 57400 7892 57452
rect 8484 57400 8536 57452
rect 9036 57400 9088 57452
rect 10232 57400 10284 57452
rect 12624 57400 12676 57452
rect 16212 57477 16221 57511
rect 16221 57477 16255 57511
rect 16255 57477 16264 57511
rect 22008 57536 22060 57588
rect 25780 57536 25832 57588
rect 26976 57536 27028 57588
rect 29368 57536 29420 57588
rect 34152 57536 34204 57588
rect 16212 57468 16264 57477
rect 15016 57400 15068 57452
rect 21916 57468 21968 57520
rect 17408 57400 17460 57452
rect 18604 57400 18656 57452
rect 19984 57400 20036 57452
rect 20996 57400 21048 57452
rect 22192 57400 22244 57452
rect 23388 57400 23440 57452
rect 24584 57400 24636 57452
rect 28172 57400 28224 57452
rect 30564 57400 30616 57452
rect 31760 57400 31812 57452
rect 32128 57400 32180 57452
rect 32956 57400 33008 57452
rect 45468 57536 45520 57588
rect 42892 57468 42944 57520
rect 50436 57536 50488 57588
rect 35348 57400 35400 57452
rect 36544 57400 36596 57452
rect 37740 57400 37792 57452
rect 38936 57400 38988 57452
rect 40132 57400 40184 57452
rect 41328 57400 41380 57452
rect 42800 57443 42852 57452
rect 42800 57409 42809 57443
rect 42809 57409 42843 57443
rect 42843 57409 42852 57443
rect 42800 57400 42852 57409
rect 43720 57400 43772 57452
rect 44916 57400 44968 57452
rect 46112 57400 46164 57452
rect 47308 57400 47360 57452
rect 48504 57400 48556 57452
rect 49700 57400 49752 57452
rect 50344 57400 50396 57452
rect 51080 57400 51132 57452
rect 52092 57400 52144 57452
rect 53288 57400 53340 57452
rect 54484 57400 54536 57452
rect 5724 57375 5776 57384
rect 5724 57341 5733 57375
rect 5733 57341 5767 57375
rect 5767 57341 5776 57375
rect 5724 57332 5776 57341
rect 8300 57375 8352 57384
rect 8300 57341 8309 57375
rect 8309 57341 8343 57375
rect 8343 57341 8352 57375
rect 8300 57332 8352 57341
rect 18972 57332 19024 57384
rect 3424 57239 3476 57248
rect 3424 57205 3433 57239
rect 3433 57205 3467 57239
rect 3467 57205 3476 57239
rect 3424 57196 3476 57205
rect 6920 57239 6972 57248
rect 6920 57205 6929 57239
rect 6929 57205 6963 57239
rect 6963 57205 6972 57239
rect 9312 57239 9364 57248
rect 6920 57196 6972 57205
rect 9312 57205 9321 57239
rect 9321 57205 9355 57239
rect 9355 57205 9364 57239
rect 9312 57196 9364 57205
rect 11888 57239 11940 57248
rect 11888 57205 11897 57239
rect 11897 57205 11931 57239
rect 11931 57205 11940 57239
rect 11888 57196 11940 57205
rect 12900 57239 12952 57248
rect 12900 57205 12909 57239
rect 12909 57205 12943 57239
rect 12943 57205 12952 57239
rect 12900 57196 12952 57205
rect 20812 57264 20864 57316
rect 28632 57332 28684 57384
rect 40040 57332 40092 57384
rect 25044 57264 25096 57316
rect 33140 57264 33192 57316
rect 37648 57264 37700 57316
rect 40500 57264 40552 57316
rect 44272 57332 44324 57384
rect 44180 57264 44232 57316
rect 55680 57400 55732 57452
rect 56876 57400 56928 57452
rect 58072 57400 58124 57452
rect 16304 57196 16356 57248
rect 17040 57239 17092 57248
rect 17040 57205 17049 57239
rect 17049 57205 17083 57239
rect 17083 57205 17092 57239
rect 17040 57196 17092 57205
rect 18880 57239 18932 57248
rect 18880 57205 18889 57239
rect 18889 57205 18923 57239
rect 18923 57205 18932 57239
rect 18880 57196 18932 57205
rect 22284 57196 22336 57248
rect 22468 57239 22520 57248
rect 22468 57205 22477 57239
rect 22477 57205 22511 57239
rect 22511 57205 22520 57239
rect 22468 57196 22520 57205
rect 24860 57239 24912 57248
rect 24860 57205 24869 57239
rect 24869 57205 24903 57239
rect 24903 57205 24912 57239
rect 24860 57196 24912 57205
rect 25136 57196 25188 57248
rect 27160 57239 27212 57248
rect 27160 57205 27169 57239
rect 27169 57205 27203 57239
rect 27203 57205 27212 57239
rect 27160 57196 27212 57205
rect 28540 57196 28592 57248
rect 29736 57239 29788 57248
rect 29736 57205 29745 57239
rect 29745 57205 29779 57239
rect 29779 57205 29788 57239
rect 29736 57196 29788 57205
rect 32496 57239 32548 57248
rect 32496 57205 32505 57239
rect 32505 57205 32539 57239
rect 32539 57205 32548 57239
rect 32496 57196 32548 57205
rect 33232 57239 33284 57248
rect 33232 57205 33241 57239
rect 33241 57205 33275 57239
rect 33275 57205 33284 57239
rect 33232 57196 33284 57205
rect 34796 57196 34848 57248
rect 35440 57196 35492 57248
rect 36544 57196 36596 57248
rect 37188 57196 37240 57248
rect 39028 57239 39080 57248
rect 39028 57205 39037 57239
rect 39037 57205 39071 57239
rect 39071 57205 39080 57239
rect 39028 57196 39080 57205
rect 41420 57239 41472 57248
rect 41420 57205 41429 57239
rect 41429 57205 41463 57239
rect 41463 57205 41472 57239
rect 41420 57196 41472 57205
rect 42800 57196 42852 57248
rect 46204 57239 46256 57248
rect 46204 57205 46213 57239
rect 46213 57205 46247 57239
rect 46247 57205 46256 57239
rect 46204 57196 46256 57205
rect 52184 57239 52236 57248
rect 52184 57205 52193 57239
rect 52193 57205 52227 57239
rect 52227 57205 52236 57239
rect 52184 57196 52236 57205
rect 53380 57239 53432 57248
rect 53380 57205 53389 57239
rect 53389 57205 53423 57239
rect 53423 57205 53432 57239
rect 53380 57196 53432 57205
rect 54576 57239 54628 57248
rect 54576 57205 54585 57239
rect 54585 57205 54619 57239
rect 54619 57205 54628 57239
rect 54576 57196 54628 57205
rect 54668 57196 54720 57248
rect 58164 57239 58216 57248
rect 58164 57205 58173 57239
rect 58173 57205 58207 57239
rect 58207 57205 58216 57239
rect 58164 57196 58216 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 1860 57035 1912 57044
rect 1860 57001 1869 57035
rect 1869 57001 1903 57035
rect 1903 57001 1912 57035
rect 1860 56992 1912 57001
rect 3056 57035 3108 57044
rect 3056 57001 3065 57035
rect 3065 57001 3099 57035
rect 3099 57001 3108 57035
rect 3056 56992 3108 57001
rect 4620 56992 4672 57044
rect 6000 57035 6052 57044
rect 6000 57001 6009 57035
rect 6009 57001 6043 57035
rect 6043 57001 6052 57035
rect 6000 56992 6052 57001
rect 6644 57035 6696 57044
rect 6644 57001 6653 57035
rect 6653 57001 6687 57035
rect 6687 57001 6696 57035
rect 6644 56992 6696 57001
rect 8484 57035 8536 57044
rect 8484 57001 8493 57035
rect 8493 57001 8527 57035
rect 8527 57001 8536 57035
rect 8484 56992 8536 57001
rect 9036 56992 9088 57044
rect 12624 57035 12676 57044
rect 12624 57001 12633 57035
rect 12633 57001 12667 57035
rect 12667 57001 12676 57035
rect 12624 56992 12676 57001
rect 15016 57035 15068 57044
rect 15016 57001 15025 57035
rect 15025 57001 15059 57035
rect 15059 57001 15068 57035
rect 15016 56992 15068 57001
rect 16304 56992 16356 57044
rect 9312 56924 9364 56976
rect 17868 56924 17920 56976
rect 19984 56992 20036 57044
rect 21640 57035 21692 57044
rect 21640 57001 21649 57035
rect 21649 57001 21683 57035
rect 21683 57001 21692 57035
rect 21640 56992 21692 57001
rect 22192 57035 22244 57044
rect 22192 57001 22201 57035
rect 22201 57001 22235 57035
rect 22235 57001 22244 57035
rect 22192 56992 22244 57001
rect 24584 57035 24636 57044
rect 24584 57001 24593 57035
rect 24593 57001 24627 57035
rect 24627 57001 24636 57035
rect 24584 56992 24636 57001
rect 26240 56992 26292 57044
rect 28172 57035 28224 57044
rect 28172 57001 28181 57035
rect 28181 57001 28215 57035
rect 28215 57001 28224 57035
rect 28172 56992 28224 57001
rect 32128 57035 32180 57044
rect 32128 57001 32137 57035
rect 32137 57001 32171 57035
rect 32171 57001 32180 57035
rect 32128 56992 32180 57001
rect 35348 57035 35400 57044
rect 35348 57001 35357 57035
rect 35357 57001 35391 57035
rect 35391 57001 35400 57035
rect 35348 56992 35400 57001
rect 36452 57035 36504 57044
rect 36452 57001 36461 57035
rect 36461 57001 36495 57035
rect 36495 57001 36504 57035
rect 36452 56992 36504 57001
rect 38936 56992 38988 57044
rect 41328 57035 41380 57044
rect 41328 57001 41337 57035
rect 41337 57001 41371 57035
rect 41371 57001 41380 57035
rect 41328 56992 41380 57001
rect 44916 56992 44968 57044
rect 47308 56992 47360 57044
rect 50344 57035 50396 57044
rect 50344 57001 50353 57035
rect 50353 57001 50387 57035
rect 50387 57001 50396 57035
rect 50344 56992 50396 57001
rect 52092 57035 52144 57044
rect 52092 57001 52101 57035
rect 52101 57001 52135 57035
rect 52135 57001 52144 57035
rect 52092 56992 52144 57001
rect 54484 57035 54536 57044
rect 54484 57001 54493 57035
rect 54493 57001 54527 57035
rect 54527 57001 54536 57035
rect 54484 56992 54536 57001
rect 56876 56992 56928 57044
rect 22100 56924 22152 56976
rect 22468 56924 22520 56976
rect 28908 56924 28960 56976
rect 42708 56924 42760 56976
rect 50436 56924 50488 56976
rect 11888 56856 11940 56908
rect 20444 56856 20496 56908
rect 22284 56856 22336 56908
rect 26424 56856 26476 56908
rect 29736 56899 29788 56908
rect 29736 56865 29745 56899
rect 29745 56865 29779 56899
rect 29779 56865 29788 56899
rect 29736 56856 29788 56865
rect 12900 56788 12952 56840
rect 20720 56788 20772 56840
rect 20812 56788 20864 56840
rect 28448 56788 28500 56840
rect 41420 56856 41472 56908
rect 39212 56831 39264 56840
rect 17408 56763 17460 56772
rect 17408 56729 17417 56763
rect 17417 56729 17451 56763
rect 17451 56729 17460 56763
rect 17408 56720 17460 56729
rect 21364 56720 21416 56772
rect 28264 56720 28316 56772
rect 38660 56720 38712 56772
rect 39212 56797 39221 56831
rect 39221 56797 39255 56831
rect 39255 56797 39264 56831
rect 39212 56788 39264 56797
rect 39304 56831 39356 56840
rect 39304 56797 39313 56831
rect 39313 56797 39347 56831
rect 39347 56797 39356 56831
rect 39304 56788 39356 56797
rect 43536 56788 43588 56840
rect 46204 56856 46256 56908
rect 44088 56831 44140 56840
rect 44088 56797 44097 56831
rect 44097 56797 44131 56831
rect 44131 56797 44140 56831
rect 57060 56831 57112 56840
rect 44088 56788 44140 56797
rect 57060 56797 57069 56831
rect 57069 56797 57103 56831
rect 57103 56797 57112 56831
rect 57060 56788 57112 56797
rect 57520 56831 57572 56840
rect 57520 56797 57529 56831
rect 57529 56797 57563 56831
rect 57563 56797 57572 56831
rect 57520 56788 57572 56797
rect 58348 56831 58400 56840
rect 58348 56797 58357 56831
rect 58357 56797 58391 56831
rect 58391 56797 58400 56831
rect 58348 56788 58400 56797
rect 39580 56720 39632 56772
rect 17040 56652 17092 56704
rect 25964 56652 26016 56704
rect 30104 56652 30156 56704
rect 35900 56652 35952 56704
rect 43444 56695 43496 56704
rect 43444 56661 43453 56695
rect 43453 56661 43487 56695
rect 43487 56661 43496 56695
rect 43444 56652 43496 56661
rect 43812 56763 43864 56772
rect 43812 56729 43821 56763
rect 43821 56729 43855 56763
rect 43855 56729 43864 56763
rect 43812 56720 43864 56729
rect 53380 56652 53432 56704
rect 56784 56652 56836 56704
rect 57888 56652 57940 56704
rect 58072 56652 58124 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 22008 56448 22060 56500
rect 17868 56380 17920 56432
rect 28724 56448 28776 56500
rect 28908 56448 28960 56500
rect 24768 56380 24820 56432
rect 21364 56312 21416 56364
rect 21824 56312 21876 56364
rect 22100 56312 22152 56364
rect 23480 56355 23532 56364
rect 23480 56321 23484 56355
rect 23484 56321 23518 56355
rect 23518 56321 23532 56355
rect 23848 56355 23900 56364
rect 23480 56312 23532 56321
rect 23848 56321 23856 56355
rect 23856 56321 23890 56355
rect 23890 56321 23900 56355
rect 23848 56312 23900 56321
rect 25044 56355 25096 56364
rect 25044 56321 25053 56355
rect 25053 56321 25087 56355
rect 25087 56321 25096 56355
rect 25044 56312 25096 56321
rect 25596 56380 25648 56432
rect 26240 56423 26292 56432
rect 26240 56389 26249 56423
rect 26249 56389 26283 56423
rect 26283 56389 26292 56423
rect 26240 56380 26292 56389
rect 29828 56380 29880 56432
rect 30196 56423 30248 56432
rect 30196 56389 30205 56423
rect 30205 56389 30239 56423
rect 30239 56389 30248 56423
rect 30196 56380 30248 56389
rect 30932 56448 30984 56500
rect 35164 56491 35216 56500
rect 35164 56457 35173 56491
rect 35173 56457 35207 56491
rect 35207 56457 35216 56491
rect 35164 56448 35216 56457
rect 32496 56380 32548 56432
rect 38384 56448 38436 56500
rect 43444 56448 43496 56500
rect 57060 56448 57112 56500
rect 35440 56423 35492 56432
rect 26148 56355 26200 56364
rect 26148 56321 26157 56355
rect 26157 56321 26191 56355
rect 26191 56321 26200 56355
rect 26148 56312 26200 56321
rect 27344 56312 27396 56364
rect 25596 56176 25648 56228
rect 28356 56355 28408 56364
rect 28356 56321 28366 56355
rect 28366 56321 28400 56355
rect 28400 56321 28408 56355
rect 28632 56355 28684 56364
rect 28356 56312 28408 56321
rect 28632 56321 28641 56355
rect 28641 56321 28675 56355
rect 28675 56321 28684 56355
rect 28632 56312 28684 56321
rect 29000 56312 29052 56364
rect 29092 56244 29144 56296
rect 30104 56312 30156 56364
rect 28724 56176 28776 56228
rect 23112 56108 23164 56160
rect 23296 56151 23348 56160
rect 23296 56117 23305 56151
rect 23305 56117 23339 56151
rect 23339 56117 23348 56151
rect 23296 56108 23348 56117
rect 25228 56108 25280 56160
rect 25872 56108 25924 56160
rect 27252 56108 27304 56160
rect 29920 56108 29972 56160
rect 30104 56176 30156 56228
rect 30564 56312 30616 56364
rect 31116 56312 31168 56364
rect 31300 56355 31352 56364
rect 31300 56321 31309 56355
rect 31309 56321 31343 56355
rect 31343 56321 31352 56355
rect 31484 56355 31536 56364
rect 31300 56312 31352 56321
rect 31484 56321 31487 56355
rect 31487 56321 31536 56355
rect 31484 56312 31536 56321
rect 32956 56355 33008 56364
rect 32956 56321 32960 56355
rect 32960 56321 32994 56355
rect 32994 56321 33008 56355
rect 32956 56312 33008 56321
rect 35440 56389 35449 56423
rect 35449 56389 35483 56423
rect 35483 56389 35492 56423
rect 35440 56380 35492 56389
rect 36544 56423 36596 56432
rect 36544 56389 36553 56423
rect 36553 56389 36587 56423
rect 36587 56389 36596 56423
rect 36544 56380 36596 56389
rect 33508 56312 33560 56364
rect 35348 56355 35400 56364
rect 35348 56321 35352 56355
rect 35352 56321 35386 56355
rect 35386 56321 35400 56355
rect 35348 56312 35400 56321
rect 35532 56355 35584 56364
rect 35532 56321 35541 56355
rect 35541 56321 35575 56355
rect 35575 56321 35584 56355
rect 35532 56312 35584 56321
rect 35716 56355 35768 56364
rect 35716 56321 35724 56355
rect 35724 56321 35758 56355
rect 35758 56321 35768 56355
rect 35716 56312 35768 56321
rect 35808 56355 35860 56364
rect 35808 56321 35817 56355
rect 35817 56321 35851 56355
rect 35851 56321 35860 56355
rect 35808 56312 35860 56321
rect 36452 56355 36504 56364
rect 36452 56321 36456 56355
rect 36456 56321 36490 56355
rect 36490 56321 36504 56355
rect 36452 56312 36504 56321
rect 36636 56355 36688 56364
rect 36636 56321 36645 56355
rect 36645 56321 36679 56355
rect 36679 56321 36688 56355
rect 38200 56380 38252 56432
rect 36636 56312 36688 56321
rect 36912 56355 36964 56364
rect 36912 56321 36921 56355
rect 36921 56321 36955 56355
rect 36955 56321 36964 56355
rect 39028 56380 39080 56432
rect 39212 56380 39264 56432
rect 36912 56312 36964 56321
rect 38660 56312 38712 56364
rect 36728 56244 36780 56296
rect 38844 56355 38896 56364
rect 38844 56321 38853 56355
rect 38853 56321 38887 56355
rect 38887 56321 38896 56355
rect 39304 56355 39356 56364
rect 38844 56312 38896 56321
rect 39304 56321 39313 56355
rect 39313 56321 39347 56355
rect 39347 56321 39356 56355
rect 39304 56312 39356 56321
rect 52184 56380 52236 56432
rect 57520 56380 57572 56432
rect 39580 56355 39632 56364
rect 38936 56244 38988 56296
rect 39580 56321 39589 56355
rect 39589 56321 39623 56355
rect 39623 56321 39632 56355
rect 39580 56312 39632 56321
rect 40500 56312 40552 56364
rect 41696 56312 41748 56364
rect 41512 56244 41564 56296
rect 42156 56312 42208 56364
rect 43444 56355 43496 56364
rect 43444 56321 43448 56355
rect 43448 56321 43482 56355
rect 43482 56321 43496 56355
rect 43444 56312 43496 56321
rect 42800 56244 42852 56296
rect 33416 56176 33468 56228
rect 36268 56219 36320 56228
rect 36268 56185 36277 56219
rect 36277 56185 36311 56219
rect 36311 56185 36320 56219
rect 36268 56176 36320 56185
rect 36636 56176 36688 56228
rect 33324 56108 33376 56160
rect 35716 56108 35768 56160
rect 41236 56151 41288 56160
rect 41236 56117 41245 56151
rect 41245 56117 41279 56151
rect 41279 56117 41288 56151
rect 41236 56108 41288 56117
rect 43628 56355 43680 56364
rect 43628 56321 43637 56355
rect 43637 56321 43671 56355
rect 43671 56321 43680 56355
rect 43628 56312 43680 56321
rect 43904 56355 43956 56364
rect 43904 56321 43913 56355
rect 43913 56321 43947 56355
rect 43947 56321 43956 56355
rect 43904 56312 43956 56321
rect 44088 56312 44140 56364
rect 57980 56312 58032 56364
rect 58440 56312 58492 56364
rect 44272 56176 44324 56228
rect 58164 56244 58216 56296
rect 58164 56151 58216 56160
rect 58164 56117 58173 56151
rect 58173 56117 58207 56151
rect 58207 56117 58216 56151
rect 58164 56108 58216 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 6920 55904 6972 55956
rect 23848 55904 23900 55956
rect 26148 55904 26200 55956
rect 28356 55904 28408 55956
rect 28448 55947 28500 55956
rect 28448 55913 28457 55947
rect 28457 55913 28491 55947
rect 28491 55913 28500 55947
rect 28448 55904 28500 55913
rect 29000 55904 29052 55956
rect 30104 55904 30156 55956
rect 32956 55904 33008 55956
rect 35072 55904 35124 55956
rect 36452 55904 36504 55956
rect 38200 55904 38252 55956
rect 42156 55904 42208 55956
rect 43904 55904 43956 55956
rect 58440 55904 58492 55956
rect 23756 55836 23808 55888
rect 24860 55768 24912 55820
rect 25780 55836 25832 55888
rect 30288 55879 30340 55888
rect 27068 55768 27120 55820
rect 27344 55768 27396 55820
rect 28540 55811 28592 55820
rect 1768 55700 1820 55752
rect 3424 55700 3476 55752
rect 23112 55743 23164 55752
rect 21364 55632 21416 55684
rect 23112 55709 23121 55743
rect 23121 55709 23155 55743
rect 23155 55709 23164 55743
rect 23112 55700 23164 55709
rect 23296 55743 23348 55752
rect 23296 55709 23305 55743
rect 23305 55709 23339 55743
rect 23339 55709 23348 55743
rect 23296 55700 23348 55709
rect 23940 55700 23992 55752
rect 24768 55743 24820 55752
rect 24768 55709 24777 55743
rect 24777 55709 24811 55743
rect 24811 55709 24820 55743
rect 24768 55700 24820 55709
rect 25228 55700 25280 55752
rect 25596 55743 25648 55752
rect 25596 55709 25605 55743
rect 25605 55709 25639 55743
rect 25639 55709 25648 55743
rect 25596 55700 25648 55709
rect 25780 55743 25832 55752
rect 25780 55709 25787 55743
rect 25787 55709 25832 55743
rect 25780 55700 25832 55709
rect 25872 55743 25924 55752
rect 25872 55709 25881 55743
rect 25881 55709 25915 55743
rect 25915 55709 25924 55743
rect 25872 55700 25924 55709
rect 26056 55743 26108 55752
rect 26056 55709 26070 55743
rect 26070 55709 26104 55743
rect 26104 55709 26108 55743
rect 28264 55743 28316 55752
rect 26056 55700 26108 55709
rect 28264 55709 28273 55743
rect 28273 55709 28307 55743
rect 28307 55709 28316 55743
rect 28264 55700 28316 55709
rect 28540 55777 28549 55811
rect 28549 55777 28583 55811
rect 28583 55777 28592 55811
rect 28540 55768 28592 55777
rect 30288 55845 30297 55879
rect 30297 55845 30331 55879
rect 30331 55845 30340 55879
rect 30288 55836 30340 55845
rect 29920 55743 29972 55752
rect 1676 55607 1728 55616
rect 1676 55573 1685 55607
rect 1685 55573 1719 55607
rect 1719 55573 1728 55607
rect 1676 55564 1728 55573
rect 18972 55564 19024 55616
rect 25964 55675 26016 55684
rect 25964 55641 25973 55675
rect 25973 55641 26007 55675
rect 26007 55641 26016 55675
rect 25964 55632 26016 55641
rect 29920 55709 29929 55743
rect 29929 55709 29963 55743
rect 29963 55709 29972 55743
rect 29920 55700 29972 55709
rect 30196 55743 30248 55752
rect 30196 55709 30199 55743
rect 30199 55709 30248 55743
rect 30196 55700 30248 55709
rect 31484 55700 31536 55752
rect 27068 55564 27120 55616
rect 30840 55607 30892 55616
rect 30840 55573 30849 55607
rect 30849 55573 30883 55607
rect 30883 55573 30892 55607
rect 30840 55564 30892 55573
rect 31300 55564 31352 55616
rect 32956 55700 33008 55752
rect 33140 55743 33192 55752
rect 33140 55709 33149 55743
rect 33149 55709 33183 55743
rect 33183 55709 33192 55743
rect 33140 55700 33192 55709
rect 41236 55836 41288 55888
rect 41880 55836 41932 55888
rect 43628 55836 43680 55888
rect 33508 55743 33560 55752
rect 33508 55709 33517 55743
rect 33517 55709 33551 55743
rect 33551 55709 33560 55743
rect 33508 55700 33560 55709
rect 34612 55700 34664 55752
rect 35072 55743 35124 55752
rect 35072 55709 35076 55743
rect 35076 55709 35110 55743
rect 35110 55709 35124 55743
rect 35072 55700 35124 55709
rect 35348 55700 35400 55752
rect 34796 55632 34848 55684
rect 35256 55675 35308 55684
rect 35256 55641 35265 55675
rect 35265 55641 35299 55675
rect 35299 55641 35308 55675
rect 35808 55700 35860 55752
rect 37188 55768 37240 55820
rect 36544 55743 36596 55752
rect 36544 55709 36553 55743
rect 36553 55709 36587 55743
rect 36587 55709 36596 55743
rect 36728 55743 36780 55752
rect 36544 55700 36596 55709
rect 36728 55709 36737 55743
rect 36737 55709 36771 55743
rect 36771 55709 36780 55743
rect 36728 55700 36780 55709
rect 36820 55743 36872 55752
rect 36820 55709 36829 55743
rect 36829 55709 36863 55743
rect 36863 55709 36872 55743
rect 40040 55768 40092 55820
rect 36820 55700 36872 55709
rect 38752 55743 38804 55752
rect 38752 55709 38761 55743
rect 38761 55709 38795 55743
rect 38795 55709 38804 55743
rect 38752 55700 38804 55709
rect 38936 55709 38964 55730
rect 38964 55709 38988 55730
rect 35256 55632 35308 55641
rect 35900 55632 35952 55684
rect 38936 55678 38988 55709
rect 39028 55737 39080 55752
rect 39028 55703 39037 55737
rect 39037 55703 39071 55737
rect 39071 55703 39080 55737
rect 39028 55700 39080 55703
rect 41512 55700 41564 55752
rect 34520 55564 34572 55616
rect 35532 55564 35584 55616
rect 37924 55607 37976 55616
rect 37924 55573 37933 55607
rect 37933 55573 37967 55607
rect 37967 55573 37976 55607
rect 37924 55564 37976 55573
rect 38752 55564 38804 55616
rect 41880 55675 41932 55684
rect 41880 55641 41889 55675
rect 41889 55641 41923 55675
rect 41923 55641 41932 55675
rect 42156 55743 42208 55752
rect 42156 55709 42165 55743
rect 42165 55709 42199 55743
rect 42199 55709 42208 55743
rect 42156 55700 42208 55709
rect 43444 55700 43496 55752
rect 45468 55768 45520 55820
rect 43904 55743 43956 55752
rect 43904 55709 43913 55743
rect 43913 55709 43947 55743
rect 43947 55709 43956 55743
rect 43904 55700 43956 55709
rect 58348 55743 58400 55752
rect 58348 55709 58357 55743
rect 58357 55709 58391 55743
rect 58391 55709 58400 55743
rect 58348 55700 58400 55709
rect 41880 55632 41932 55641
rect 42892 55632 42944 55684
rect 42708 55564 42760 55616
rect 43260 55607 43312 55616
rect 43260 55573 43269 55607
rect 43269 55573 43303 55607
rect 43303 55573 43312 55607
rect 43260 55564 43312 55573
rect 54576 55564 54628 55616
rect 58532 55564 58584 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 8300 55292 8352 55344
rect 30840 55360 30892 55412
rect 41052 55360 41104 55412
rect 3516 55224 3568 55276
rect 21364 55224 21416 55276
rect 21824 55224 21876 55276
rect 35256 55292 35308 55344
rect 58348 55360 58400 55412
rect 54668 55292 54720 55344
rect 27344 55224 27396 55276
rect 29000 55224 29052 55276
rect 32680 55267 32732 55276
rect 32680 55233 32689 55267
rect 32689 55233 32723 55267
rect 32723 55233 32732 55267
rect 32680 55224 32732 55233
rect 31852 55156 31904 55208
rect 36544 55224 36596 55276
rect 37740 55224 37792 55276
rect 38660 55224 38712 55276
rect 40040 55224 40092 55276
rect 43444 55224 43496 55276
rect 43720 55267 43772 55276
rect 43720 55233 43729 55267
rect 43729 55233 43763 55267
rect 43763 55233 43772 55267
rect 43720 55224 43772 55233
rect 43996 55267 44048 55276
rect 43996 55233 44005 55267
rect 44005 55233 44039 55267
rect 44039 55233 44048 55267
rect 43996 55224 44048 55233
rect 44180 55224 44232 55276
rect 57980 55224 58032 55276
rect 1676 55063 1728 55072
rect 1676 55029 1685 55063
rect 1685 55029 1719 55063
rect 1719 55029 1728 55063
rect 1676 55020 1728 55029
rect 32404 55020 32456 55072
rect 36820 55020 36872 55072
rect 40316 55063 40368 55072
rect 40316 55029 40325 55063
rect 40325 55029 40359 55063
rect 40359 55029 40368 55063
rect 40316 55020 40368 55029
rect 40868 55063 40920 55072
rect 40868 55029 40877 55063
rect 40877 55029 40911 55063
rect 40911 55029 40920 55063
rect 40868 55020 40920 55029
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 25228 54816 25280 54868
rect 40316 54816 40368 54868
rect 41052 54816 41104 54868
rect 41328 54859 41380 54868
rect 41328 54825 41337 54859
rect 41337 54825 41371 54859
rect 41371 54825 41380 54859
rect 41328 54816 41380 54825
rect 41512 54859 41564 54868
rect 41512 54825 41521 54859
rect 41521 54825 41555 54859
rect 41555 54825 41564 54859
rect 41512 54816 41564 54825
rect 33232 54748 33284 54800
rect 25136 54680 25188 54732
rect 27896 54680 27948 54732
rect 34520 54680 34572 54732
rect 21364 54655 21416 54664
rect 21364 54621 21373 54655
rect 21373 54621 21407 54655
rect 21407 54621 21416 54655
rect 21364 54612 21416 54621
rect 24768 54655 24820 54664
rect 24768 54621 24777 54655
rect 24777 54621 24811 54655
rect 24811 54621 24820 54655
rect 24768 54612 24820 54621
rect 32404 54655 32456 54664
rect 32404 54621 32413 54655
rect 32413 54621 32447 54655
rect 32447 54621 32456 54655
rect 32404 54612 32456 54621
rect 35348 54655 35400 54664
rect 35348 54621 35352 54655
rect 35352 54621 35386 54655
rect 35386 54621 35400 54655
rect 35348 54612 35400 54621
rect 42156 54748 42208 54800
rect 35716 54655 35768 54664
rect 35716 54621 35724 54655
rect 35724 54621 35758 54655
rect 35758 54621 35768 54655
rect 35716 54612 35768 54621
rect 35808 54655 35860 54664
rect 35808 54621 35817 54655
rect 35817 54621 35851 54655
rect 35851 54621 35860 54655
rect 35808 54612 35860 54621
rect 40040 54612 40092 54664
rect 20444 54544 20496 54596
rect 25044 54544 25096 54596
rect 23572 54476 23624 54528
rect 25136 54476 25188 54528
rect 32312 54519 32364 54528
rect 32312 54485 32321 54519
rect 32321 54485 32355 54519
rect 32355 54485 32364 54519
rect 32312 54476 32364 54485
rect 32772 54476 32824 54528
rect 43260 54612 43312 54664
rect 36452 54476 36504 54528
rect 37924 54476 37976 54528
rect 38568 54476 38620 54528
rect 39396 54519 39448 54528
rect 39396 54485 39405 54519
rect 39405 54485 39439 54519
rect 39439 54485 39448 54519
rect 40868 54544 40920 54596
rect 39396 54476 39448 54485
rect 41052 54476 41104 54528
rect 58348 54519 58400 54528
rect 58348 54485 58357 54519
rect 58357 54485 58391 54519
rect 58391 54485 58400 54519
rect 58348 54476 58400 54485
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 21916 54272 21968 54324
rect 20720 54204 20772 54256
rect 24768 54272 24820 54324
rect 1676 54043 1728 54052
rect 1676 54009 1685 54043
rect 1685 54009 1719 54043
rect 1719 54009 1728 54043
rect 1676 54000 1728 54009
rect 21364 54136 21416 54188
rect 23572 54179 23624 54188
rect 23572 54145 23581 54179
rect 23581 54145 23615 54179
rect 23615 54145 23624 54179
rect 23572 54136 23624 54145
rect 25044 54247 25096 54256
rect 25044 54213 25053 54247
rect 25053 54213 25087 54247
rect 25087 54213 25096 54247
rect 25044 54204 25096 54213
rect 23940 54136 23992 54188
rect 24676 54136 24728 54188
rect 24860 54179 24912 54188
rect 24860 54145 24864 54179
rect 24864 54145 24898 54179
rect 24898 54145 24912 54179
rect 24860 54136 24912 54145
rect 18880 54068 18932 54120
rect 25136 54179 25188 54188
rect 25136 54145 25181 54179
rect 25181 54145 25188 54179
rect 25136 54136 25188 54145
rect 25596 54136 25648 54188
rect 28264 54272 28316 54324
rect 32312 54272 32364 54324
rect 26424 54204 26476 54256
rect 27896 54204 27948 54256
rect 35716 54272 35768 54324
rect 37740 54272 37792 54324
rect 41880 54272 41932 54324
rect 27160 54136 27212 54188
rect 27344 54179 27396 54188
rect 27344 54145 27348 54179
rect 27348 54145 27382 54179
rect 27382 54145 27396 54179
rect 27344 54136 27396 54145
rect 29092 54136 29144 54188
rect 31852 54136 31904 54188
rect 28632 54068 28684 54120
rect 32772 54136 32824 54188
rect 32956 54179 33008 54188
rect 32956 54145 32965 54179
rect 32965 54145 32999 54179
rect 32999 54145 33008 54179
rect 32956 54136 33008 54145
rect 36728 54204 36780 54256
rect 36820 54204 36872 54256
rect 36452 54136 36504 54188
rect 37648 54179 37700 54188
rect 37648 54145 37657 54179
rect 37657 54145 37691 54179
rect 37691 54145 37700 54179
rect 37648 54136 37700 54145
rect 37740 54179 37792 54188
rect 37740 54145 37749 54179
rect 37749 54145 37783 54179
rect 37783 54145 37792 54179
rect 38660 54204 38712 54256
rect 39396 54204 39448 54256
rect 37740 54136 37792 54145
rect 38568 54179 38620 54188
rect 36728 54068 36780 54120
rect 38568 54145 38577 54179
rect 38577 54145 38611 54179
rect 38611 54145 38620 54179
rect 38568 54136 38620 54145
rect 40316 54136 40368 54188
rect 58348 54179 58400 54188
rect 58348 54145 58357 54179
rect 58357 54145 58391 54179
rect 58391 54145 58400 54179
rect 58348 54136 58400 54145
rect 25228 54000 25280 54052
rect 27344 54000 27396 54052
rect 30472 54000 30524 54052
rect 4804 53932 4856 53984
rect 23388 53932 23440 53984
rect 24124 53975 24176 53984
rect 24124 53941 24133 53975
rect 24133 53941 24167 53975
rect 24167 53941 24176 53975
rect 24124 53932 24176 53941
rect 27068 53932 27120 53984
rect 29000 53932 29052 53984
rect 32312 54000 32364 54052
rect 32404 54000 32456 54052
rect 32680 53975 32732 53984
rect 32680 53941 32689 53975
rect 32689 53941 32723 53975
rect 32723 53941 32732 53975
rect 32680 53932 32732 53941
rect 34612 54000 34664 54052
rect 35808 54000 35860 54052
rect 40040 53932 40092 53984
rect 41328 53932 41380 53984
rect 59176 53932 59228 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 27344 53728 27396 53780
rect 28448 53728 28500 53780
rect 24676 53592 24728 53644
rect 11704 53524 11756 53576
rect 23388 53524 23440 53576
rect 27068 53567 27120 53576
rect 27068 53533 27077 53567
rect 27077 53533 27111 53567
rect 27111 53533 27120 53567
rect 27068 53524 27120 53533
rect 28632 53635 28684 53644
rect 28632 53601 28641 53635
rect 28641 53601 28675 53635
rect 28675 53601 28684 53635
rect 28632 53592 28684 53601
rect 36728 53728 36780 53780
rect 38660 53771 38712 53780
rect 38660 53737 38669 53771
rect 38669 53737 38703 53771
rect 38703 53737 38712 53771
rect 38660 53728 38712 53737
rect 40316 53728 40368 53780
rect 30104 53703 30156 53712
rect 30104 53669 30113 53703
rect 30113 53669 30147 53703
rect 30147 53669 30156 53703
rect 30104 53660 30156 53669
rect 28908 53524 28960 53576
rect 29736 53524 29788 53576
rect 30012 53567 30064 53576
rect 30012 53533 30021 53567
rect 30021 53533 30055 53567
rect 30055 53533 30064 53567
rect 30012 53524 30064 53533
rect 30472 53524 30524 53576
rect 30564 53567 30616 53576
rect 30564 53533 30573 53567
rect 30573 53533 30607 53567
rect 30607 53533 30616 53567
rect 30564 53524 30616 53533
rect 32680 53592 32732 53644
rect 31852 53524 31904 53576
rect 32404 53567 32456 53576
rect 32404 53533 32413 53567
rect 32413 53533 32447 53567
rect 32447 53533 32456 53567
rect 32404 53524 32456 53533
rect 39396 53524 39448 53576
rect 58348 53567 58400 53576
rect 58348 53533 58357 53567
rect 58357 53533 58391 53567
rect 58391 53533 58400 53567
rect 58348 53524 58400 53533
rect 1676 53431 1728 53440
rect 1676 53397 1685 53431
rect 1685 53397 1719 53431
rect 1719 53397 1728 53431
rect 1676 53388 1728 53397
rect 5724 53388 5776 53440
rect 30932 53456 30984 53508
rect 38384 53499 38436 53508
rect 38384 53465 38393 53499
rect 38393 53465 38427 53499
rect 38427 53465 38436 53499
rect 40040 53499 40092 53508
rect 38384 53456 38436 53465
rect 40040 53465 40049 53499
rect 40049 53465 40083 53499
rect 40083 53465 40092 53499
rect 40040 53456 40092 53465
rect 28448 53388 28500 53440
rect 31944 53431 31996 53440
rect 31944 53397 31953 53431
rect 31953 53397 31987 53431
rect 31987 53397 31996 53431
rect 31944 53388 31996 53397
rect 59636 53388 59688 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 28264 53184 28316 53236
rect 29736 53184 29788 53236
rect 30196 53184 30248 53236
rect 31944 53184 31996 53236
rect 28908 53048 28960 53100
rect 30564 53116 30616 53168
rect 30012 53091 30064 53100
rect 30012 53057 30021 53091
rect 30021 53057 30055 53091
rect 30055 53057 30064 53091
rect 30012 53048 30064 53057
rect 31852 53048 31904 53100
rect 27896 52844 27948 52896
rect 28908 52844 28960 52896
rect 30472 52844 30524 52896
rect 38384 52844 38436 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 1676 52615 1728 52624
rect 1676 52581 1685 52615
rect 1685 52581 1719 52615
rect 1719 52581 1728 52615
rect 1676 52572 1728 52581
rect 59268 52572 59320 52624
rect 5540 52436 5592 52488
rect 58348 52479 58400 52488
rect 58348 52445 58357 52479
rect 58357 52445 58391 52479
rect 58391 52445 58400 52479
rect 58348 52436 58400 52445
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 1676 51799 1728 51808
rect 1676 51765 1685 51799
rect 1685 51765 1719 51799
rect 1719 51765 1728 51799
rect 1676 51756 1728 51765
rect 58348 52003 58400 52012
rect 58348 51969 58357 52003
rect 58357 51969 58391 52003
rect 58391 51969 58400 52003
rect 58348 51960 58400 51969
rect 4896 51756 4948 51808
rect 58992 51756 59044 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 58348 51255 58400 51264
rect 58348 51221 58357 51255
rect 58357 51221 58391 51255
rect 58391 51221 58400 51255
rect 58348 51212 58400 51221
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 16580 50872 16632 50924
rect 58348 50915 58400 50924
rect 58348 50881 58357 50915
rect 58357 50881 58391 50915
rect 58391 50881 58400 50915
rect 58348 50872 58400 50881
rect 1676 50779 1728 50788
rect 1676 50745 1685 50779
rect 1685 50745 1719 50779
rect 1719 50745 1728 50779
rect 1676 50736 1728 50745
rect 58900 50668 58952 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 58164 50328 58216 50380
rect 58624 50328 58676 50380
rect 58348 50303 58400 50312
rect 58348 50269 58357 50303
rect 58357 50269 58391 50303
rect 58391 50269 58400 50303
rect 58348 50260 58400 50269
rect 1676 50167 1728 50176
rect 1676 50133 1685 50167
rect 1685 50133 1719 50167
rect 1719 50133 1728 50167
rect 1676 50124 1728 50133
rect 2412 50167 2464 50176
rect 2412 50133 2421 50167
rect 2421 50133 2455 50167
rect 2455 50133 2464 50167
rect 2412 50124 2464 50133
rect 59084 50124 59136 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 2412 49920 2464 49972
rect 13452 49920 13504 49972
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 58348 49215 58400 49224
rect 58348 49181 58357 49215
rect 58357 49181 58391 49215
rect 58391 49181 58400 49215
rect 58348 49172 58400 49181
rect 1676 49079 1728 49088
rect 1676 49045 1685 49079
rect 1685 49045 1719 49079
rect 1719 49045 1728 49079
rect 1676 49036 1728 49045
rect 2412 49079 2464 49088
rect 2412 49045 2421 49079
rect 2421 49045 2455 49079
rect 2455 49045 2464 49079
rect 2412 49036 2464 49045
rect 58808 49036 58860 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 2412 48832 2464 48884
rect 13360 48832 13412 48884
rect 2412 48696 2464 48748
rect 58348 48739 58400 48748
rect 58348 48705 58357 48739
rect 58357 48705 58391 48739
rect 58391 48705 58400 48739
rect 58348 48696 58400 48705
rect 1676 48535 1728 48544
rect 1676 48501 1685 48535
rect 1685 48501 1719 48535
rect 1719 48501 1728 48535
rect 1676 48492 1728 48501
rect 2412 48535 2464 48544
rect 2412 48501 2421 48535
rect 2421 48501 2455 48535
rect 2455 48501 2464 48535
rect 2412 48492 2464 48501
rect 59820 48492 59872 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 58348 47991 58400 48000
rect 58348 47957 58357 47991
rect 58357 47957 58391 47991
rect 58391 47957 58400 47991
rect 58348 47948 58400 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 58348 47651 58400 47660
rect 1676 47515 1728 47524
rect 1676 47481 1685 47515
rect 1685 47481 1719 47515
rect 1719 47481 1728 47515
rect 1676 47472 1728 47481
rect 58348 47617 58357 47651
rect 58357 47617 58391 47651
rect 58391 47617 58400 47651
rect 58348 47608 58400 47617
rect 5540 47540 5592 47592
rect 17132 47540 17184 47592
rect 9220 47404 9272 47456
rect 55956 47404 56008 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 59544 47132 59596 47184
rect 58348 47039 58400 47048
rect 58348 47005 58357 47039
rect 58357 47005 58391 47039
rect 58391 47005 58400 47039
rect 58348 46996 58400 47005
rect 6644 46928 6696 46980
rect 1676 46903 1728 46912
rect 1676 46869 1685 46903
rect 1685 46869 1719 46903
rect 1719 46869 1728 46903
rect 1676 46860 1728 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 1860 45951 1912 45960
rect 1860 45917 1869 45951
rect 1869 45917 1903 45951
rect 1903 45917 1912 45951
rect 1860 45908 1912 45917
rect 58348 45951 58400 45960
rect 58348 45917 58357 45951
rect 58357 45917 58391 45951
rect 58391 45917 58400 45951
rect 58348 45908 58400 45917
rect 1676 45815 1728 45824
rect 1676 45781 1685 45815
rect 1685 45781 1719 45815
rect 1719 45781 1728 45815
rect 1676 45772 1728 45781
rect 58716 45772 58768 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 3516 45568 3568 45620
rect 7472 45568 7524 45620
rect 1676 45271 1728 45280
rect 1676 45237 1685 45271
rect 1685 45237 1719 45271
rect 1719 45237 1728 45271
rect 1676 45228 1728 45237
rect 58348 45475 58400 45484
rect 58348 45441 58357 45475
rect 58357 45441 58391 45475
rect 58391 45441 58400 45475
rect 58348 45432 58400 45441
rect 9312 45228 9364 45280
rect 57244 45228 57296 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 4896 44820 4948 44872
rect 18788 44820 18840 44872
rect 58348 44727 58400 44736
rect 58348 44693 58357 44727
rect 58357 44693 58391 44727
rect 58391 44693 58400 44727
rect 58348 44684 58400 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 1952 44344 2004 44396
rect 58348 44387 58400 44396
rect 58348 44353 58357 44387
rect 58357 44353 58391 44387
rect 58391 44353 58400 44387
rect 58348 44344 58400 44353
rect 57980 44276 58032 44328
rect 58624 44276 58676 44328
rect 1676 44251 1728 44260
rect 1676 44217 1685 44251
rect 1685 44217 1719 44251
rect 1719 44217 1728 44251
rect 1676 44208 1728 44217
rect 58624 44140 58676 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 1676 43639 1728 43648
rect 1676 43605 1685 43639
rect 1685 43605 1719 43639
rect 1719 43605 1728 43639
rect 1676 43596 1728 43605
rect 58348 43775 58400 43784
rect 58348 43741 58357 43775
rect 58357 43741 58391 43775
rect 58391 43741 58400 43775
rect 58348 43732 58400 43741
rect 5264 43596 5316 43648
rect 59728 43596 59780 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 1676 42551 1728 42560
rect 1676 42517 1685 42551
rect 1685 42517 1719 42551
rect 1719 42517 1728 42551
rect 1676 42508 1728 42517
rect 58348 42687 58400 42696
rect 58348 42653 58357 42687
rect 58357 42653 58391 42687
rect 58391 42653 58400 42687
rect 58348 42644 58400 42653
rect 6276 42508 6328 42560
rect 56968 42508 57020 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 1676 42007 1728 42016
rect 1676 41973 1685 42007
rect 1685 41973 1719 42007
rect 1719 41973 1728 42007
rect 1676 41964 1728 41973
rect 58348 42211 58400 42220
rect 58348 42177 58357 42211
rect 58357 42177 58391 42211
rect 58391 42177 58400 42211
rect 58348 42168 58400 42177
rect 2504 41964 2556 42016
rect 59452 41964 59504 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 2504 41760 2556 41812
rect 13912 41760 13964 41812
rect 58348 41463 58400 41472
rect 58348 41429 58357 41463
rect 58357 41429 58391 41463
rect 58391 41429 58400 41463
rect 58348 41420 58400 41429
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 58348 41123 58400 41132
rect 1676 40987 1728 40996
rect 1676 40953 1685 40987
rect 1685 40953 1719 40987
rect 1719 40953 1728 40987
rect 1676 40944 1728 40953
rect 58348 41089 58357 41123
rect 58357 41089 58391 41123
rect 58391 41089 58400 41123
rect 58348 41080 58400 41089
rect 3516 40876 3568 40928
rect 58164 40919 58216 40928
rect 58164 40885 58173 40919
rect 58173 40885 58207 40919
rect 58207 40885 58216 40919
rect 58164 40876 58216 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 1676 40375 1728 40384
rect 1676 40341 1685 40375
rect 1685 40341 1719 40375
rect 1719 40341 1728 40375
rect 1676 40332 1728 40341
rect 58348 40511 58400 40520
rect 58348 40477 58357 40511
rect 58357 40477 58391 40511
rect 58391 40477 58400 40511
rect 58348 40468 58400 40477
rect 3700 40332 3752 40384
rect 57336 40332 57388 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 3700 40128 3752 40180
rect 11796 40128 11848 40180
rect 58348 39856 58400 39908
rect 57888 39788 57940 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 56692 39448 56744 39500
rect 1676 39287 1728 39296
rect 1676 39253 1685 39287
rect 1685 39253 1719 39287
rect 1719 39253 1728 39287
rect 1676 39244 1728 39253
rect 56232 39380 56284 39432
rect 57980 39584 58032 39636
rect 58348 39423 58400 39432
rect 58348 39389 58357 39423
rect 58357 39389 58391 39423
rect 58391 39389 58400 39423
rect 58348 39380 58400 39389
rect 56140 39355 56192 39364
rect 56140 39321 56149 39355
rect 56149 39321 56183 39355
rect 56183 39321 56192 39355
rect 56140 39312 56192 39321
rect 59820 39312 59872 39364
rect 3424 39244 3476 39296
rect 55680 39244 55732 39296
rect 57428 39244 57480 39296
rect 57612 39244 57664 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 56140 39040 56192 39092
rect 57888 38904 57940 38956
rect 58348 38947 58400 38956
rect 58348 38913 58357 38947
rect 58357 38913 58391 38947
rect 58391 38913 58400 38947
rect 58348 38904 58400 38913
rect 18236 38768 18288 38820
rect 1676 38743 1728 38752
rect 1676 38709 1685 38743
rect 1685 38709 1719 38743
rect 1719 38709 1728 38743
rect 1676 38700 1728 38709
rect 56692 38743 56744 38752
rect 56692 38709 56701 38743
rect 56701 38709 56735 38743
rect 56735 38709 56744 38743
rect 56692 38700 56744 38709
rect 57520 38743 57572 38752
rect 57520 38709 57529 38743
rect 57529 38709 57563 38743
rect 57563 38709 57572 38743
rect 57520 38700 57572 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 55496 38496 55548 38548
rect 56232 38539 56284 38548
rect 56232 38505 56241 38539
rect 56241 38505 56275 38539
rect 56275 38505 56284 38539
rect 56232 38496 56284 38505
rect 56692 38360 56744 38412
rect 57612 38292 57664 38344
rect 57888 38335 57940 38344
rect 57888 38301 57897 38335
rect 57897 38301 57931 38335
rect 57931 38301 57940 38335
rect 57888 38292 57940 38301
rect 58256 38292 58308 38344
rect 59176 38292 59228 38344
rect 57980 38224 58032 38276
rect 58808 38224 58860 38276
rect 56600 38156 56652 38208
rect 59176 38156 59228 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 55772 37952 55824 38004
rect 55956 37952 56008 38004
rect 56784 37952 56836 38004
rect 57888 37952 57940 38004
rect 58072 37952 58124 38004
rect 1676 37723 1728 37732
rect 1676 37689 1685 37723
rect 1685 37689 1719 37723
rect 1719 37689 1728 37723
rect 1676 37680 1728 37689
rect 55496 37859 55548 37868
rect 55496 37825 55505 37859
rect 55505 37825 55539 37859
rect 55539 37825 55548 37859
rect 55496 37816 55548 37825
rect 56784 37816 56836 37868
rect 57520 37816 57572 37868
rect 58348 37859 58400 37868
rect 58348 37825 58357 37859
rect 58357 37825 58391 37859
rect 58391 37825 58400 37859
rect 58348 37816 58400 37825
rect 56692 37748 56744 37800
rect 2596 37612 2648 37664
rect 54668 37612 54720 37664
rect 55864 37612 55916 37664
rect 59820 37612 59872 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2596 37408 2648 37460
rect 15200 37408 15252 37460
rect 56232 37451 56284 37460
rect 56232 37417 56241 37451
rect 56241 37417 56275 37451
rect 56275 37417 56284 37451
rect 56232 37408 56284 37417
rect 56968 37340 57020 37392
rect 56692 37272 56744 37324
rect 57888 37247 57940 37256
rect 1676 37111 1728 37120
rect 1676 37077 1685 37111
rect 1685 37077 1719 37111
rect 1719 37077 1728 37111
rect 1676 37068 1728 37077
rect 56232 37136 56284 37188
rect 57428 37179 57480 37188
rect 57428 37145 57437 37179
rect 57437 37145 57471 37179
rect 57471 37145 57480 37179
rect 57428 37136 57480 37145
rect 57888 37213 57897 37247
rect 57897 37213 57931 37247
rect 57931 37213 57940 37247
rect 57888 37204 57940 37213
rect 57980 37136 58032 37188
rect 59544 37136 59596 37188
rect 2504 37068 2556 37120
rect 58072 37068 58124 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 56692 36907 56744 36916
rect 56692 36873 56701 36907
rect 56701 36873 56735 36907
rect 56735 36873 56744 36907
rect 56692 36864 56744 36873
rect 57428 36864 57480 36916
rect 58348 36771 58400 36780
rect 58348 36737 58357 36771
rect 58357 36737 58391 36771
rect 58391 36737 58400 36771
rect 58348 36728 58400 36737
rect 58992 36524 59044 36576
rect 59360 36524 59412 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1676 36023 1728 36032
rect 1676 35989 1685 36023
rect 1685 35989 1719 36023
rect 1719 35989 1728 36023
rect 1676 35980 1728 35989
rect 58348 36159 58400 36168
rect 58348 36125 58357 36159
rect 58357 36125 58391 36159
rect 58391 36125 58400 36159
rect 58348 36116 58400 36125
rect 7564 35980 7616 36032
rect 57704 36023 57756 36032
rect 57704 35989 57713 36023
rect 57713 35989 57747 36023
rect 57747 35989 57756 36023
rect 57704 35980 57756 35989
rect 58164 36023 58216 36032
rect 58164 35989 58173 36023
rect 58173 35989 58207 36023
rect 58207 35989 58216 36023
rect 58164 35980 58216 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 56692 35776 56744 35828
rect 57428 35776 57480 35828
rect 57980 35776 58032 35828
rect 58532 35776 58584 35828
rect 7012 35640 7064 35692
rect 57704 35640 57756 35692
rect 58348 35683 58400 35692
rect 58348 35649 58357 35683
rect 58357 35649 58391 35683
rect 58391 35649 58400 35683
rect 58348 35640 58400 35649
rect 1676 35479 1728 35488
rect 1676 35445 1685 35479
rect 1685 35445 1719 35479
rect 1719 35445 1728 35479
rect 1676 35436 1728 35445
rect 57612 35436 57664 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 53932 35232 53984 35284
rect 56232 35232 56284 35284
rect 57152 35232 57204 35284
rect 58716 35232 58768 35284
rect 3516 35164 3568 35216
rect 11244 35164 11296 35216
rect 57152 35139 57204 35148
rect 57152 35105 57170 35139
rect 57170 35105 57204 35139
rect 57152 35096 57204 35105
rect 57980 35164 58032 35216
rect 57520 35139 57572 35148
rect 57520 35105 57529 35139
rect 57529 35105 57563 35139
rect 57563 35105 57572 35139
rect 58164 35139 58216 35148
rect 57520 35096 57572 35105
rect 58164 35105 58173 35139
rect 58173 35105 58207 35139
rect 58207 35105 58216 35139
rect 58164 35096 58216 35105
rect 59084 35096 59136 35148
rect 54576 35071 54628 35080
rect 54576 35037 54585 35071
rect 54585 35037 54619 35071
rect 54619 35037 54628 35071
rect 54576 35028 54628 35037
rect 54760 35028 54812 35080
rect 58808 35028 58860 35080
rect 52368 34960 52420 35012
rect 59084 34892 59136 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 53932 34731 53984 34740
rect 53932 34697 53941 34731
rect 53941 34697 53975 34731
rect 53975 34697 53984 34731
rect 53932 34688 53984 34697
rect 54760 34688 54812 34740
rect 55220 34688 55272 34740
rect 57244 34688 57296 34740
rect 52368 34595 52420 34604
rect 52368 34561 52377 34595
rect 52377 34561 52411 34595
rect 52411 34561 52420 34595
rect 52368 34552 52420 34561
rect 8208 34484 8260 34536
rect 51448 34484 51500 34536
rect 55220 34595 55272 34604
rect 55220 34561 55238 34595
rect 55238 34561 55272 34595
rect 55220 34552 55272 34561
rect 57612 34620 57664 34672
rect 56048 34527 56100 34536
rect 56048 34493 56057 34527
rect 56057 34493 56091 34527
rect 56091 34493 56100 34527
rect 56048 34484 56100 34493
rect 57888 34552 57940 34604
rect 58440 34484 58492 34536
rect 1676 34459 1728 34468
rect 1676 34425 1685 34459
rect 1685 34425 1719 34459
rect 1719 34425 1728 34459
rect 1676 34416 1728 34425
rect 55588 34459 55640 34468
rect 55588 34425 55597 34459
rect 55597 34425 55631 34459
rect 55631 34425 55640 34459
rect 55588 34416 55640 34425
rect 56692 34416 56744 34468
rect 56968 34416 57020 34468
rect 57520 34416 57572 34468
rect 58348 34391 58400 34400
rect 58348 34357 58357 34391
rect 58357 34357 58391 34391
rect 58391 34357 58400 34391
rect 58348 34348 58400 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 55588 34144 55640 34196
rect 56600 34076 56652 34128
rect 2688 33940 2740 33992
rect 58440 33940 58492 33992
rect 1676 33847 1728 33856
rect 1676 33813 1685 33847
rect 1685 33813 1719 33847
rect 1719 33813 1728 33847
rect 1676 33804 1728 33813
rect 57888 33804 57940 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 56232 33643 56284 33652
rect 56232 33609 56241 33643
rect 56241 33609 56275 33643
rect 56275 33609 56284 33643
rect 56232 33600 56284 33609
rect 56692 33643 56744 33652
rect 56692 33609 56701 33643
rect 56701 33609 56735 33643
rect 56735 33609 56744 33643
rect 56692 33600 56744 33609
rect 57428 33600 57480 33652
rect 58256 33600 58308 33652
rect 57888 33464 57940 33516
rect 57980 33260 58032 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 56140 33056 56192 33108
rect 56692 33056 56744 33108
rect 57704 33056 57756 33108
rect 56232 32920 56284 32972
rect 58624 32988 58676 33040
rect 57704 32963 57756 32972
rect 57704 32929 57713 32963
rect 57713 32929 57747 32963
rect 57747 32929 57756 32963
rect 58348 32963 58400 32972
rect 57704 32920 57756 32929
rect 58348 32929 58357 32963
rect 58357 32929 58391 32963
rect 58391 32929 58400 32963
rect 58348 32920 58400 32929
rect 2228 32852 2280 32904
rect 57428 32895 57480 32904
rect 57428 32861 57437 32895
rect 57437 32861 57471 32895
rect 57471 32861 57480 32895
rect 57428 32852 57480 32861
rect 58624 32852 58676 32904
rect 1676 32759 1728 32768
rect 1676 32725 1685 32759
rect 1685 32725 1719 32759
rect 1719 32725 1728 32759
rect 1676 32716 1728 32725
rect 55864 32716 55916 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 56968 32512 57020 32564
rect 59728 32512 59780 32564
rect 3424 32444 3476 32496
rect 16948 32444 17000 32496
rect 56600 32487 56652 32496
rect 56600 32453 56609 32487
rect 56609 32453 56643 32487
rect 56643 32453 56652 32487
rect 56600 32444 56652 32453
rect 4620 32376 4672 32428
rect 55864 32376 55916 32428
rect 56232 32376 56284 32428
rect 58164 32376 58216 32428
rect 58348 32419 58400 32428
rect 58348 32385 58357 32419
rect 58357 32385 58391 32419
rect 58391 32385 58400 32419
rect 58348 32376 58400 32385
rect 49056 32308 49108 32360
rect 56692 32308 56744 32360
rect 1676 32215 1728 32224
rect 1676 32181 1685 32215
rect 1685 32181 1719 32215
rect 1719 32181 1728 32215
rect 1676 32172 1728 32181
rect 55956 32172 56008 32224
rect 58256 32172 58308 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 56232 31968 56284 32020
rect 58348 32011 58400 32020
rect 58348 31977 58357 32011
rect 58357 31977 58391 32011
rect 58391 31977 58400 32011
rect 58348 31968 58400 31977
rect 58164 31900 58216 31952
rect 59636 31900 59688 31952
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 58440 31424 58492 31476
rect 59268 31424 59320 31476
rect 4068 31288 4120 31340
rect 58164 31331 58216 31340
rect 58164 31297 58173 31331
rect 58173 31297 58207 31331
rect 58207 31297 58216 31331
rect 58164 31288 58216 31297
rect 1676 31195 1728 31204
rect 1676 31161 1685 31195
rect 1685 31161 1719 31195
rect 1719 31161 1728 31195
rect 1676 31152 1728 31161
rect 58348 31127 58400 31136
rect 58348 31093 58357 31127
rect 58357 31093 58391 31127
rect 58391 31093 58400 31127
rect 58348 31084 58400 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 57612 30744 57664 30796
rect 2320 30676 2372 30728
rect 57980 30676 58032 30728
rect 1676 30583 1728 30592
rect 1676 30549 1685 30583
rect 1685 30549 1719 30583
rect 1719 30549 1728 30583
rect 1676 30540 1728 30549
rect 57060 30608 57112 30660
rect 57244 30608 57296 30660
rect 58440 30608 58492 30660
rect 56784 30583 56836 30592
rect 56784 30549 56793 30583
rect 56793 30549 56827 30583
rect 56827 30549 56836 30583
rect 56784 30540 56836 30549
rect 56968 30540 57020 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 58164 30243 58216 30252
rect 58164 30209 58173 30243
rect 58173 30209 58207 30243
rect 58207 30209 58216 30243
rect 58164 30200 58216 30209
rect 56876 30039 56928 30048
rect 56876 30005 56885 30039
rect 56885 30005 56919 30039
rect 56919 30005 56928 30039
rect 56876 29996 56928 30005
rect 57244 29996 57296 30048
rect 57612 29996 57664 30048
rect 58440 29996 58492 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 56876 29656 56928 29708
rect 14648 29588 14700 29640
rect 57244 29588 57296 29640
rect 57520 29656 57572 29708
rect 57612 29699 57664 29708
rect 57612 29665 57621 29699
rect 57621 29665 57655 29699
rect 57655 29665 57664 29699
rect 58256 29699 58308 29708
rect 57612 29656 57664 29665
rect 58256 29665 58265 29699
rect 58265 29665 58299 29699
rect 58299 29665 58308 29699
rect 58256 29656 58308 29665
rect 58716 29588 58768 29640
rect 1676 29495 1728 29504
rect 1676 29461 1685 29495
rect 1685 29461 1719 29495
rect 1719 29461 1728 29495
rect 1676 29452 1728 29461
rect 9956 29495 10008 29504
rect 9956 29461 9965 29495
rect 9965 29461 9999 29495
rect 9999 29461 10008 29495
rect 9956 29452 10008 29461
rect 10692 29452 10744 29504
rect 57428 29452 57480 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 3056 29248 3108 29300
rect 9956 29248 10008 29300
rect 10692 29291 10744 29300
rect 10692 29257 10701 29291
rect 10701 29257 10735 29291
rect 10735 29257 10744 29291
rect 10692 29248 10744 29257
rect 58992 29248 59044 29300
rect 6920 29155 6972 29164
rect 1676 29019 1728 29028
rect 1676 28985 1685 29019
rect 1685 28985 1719 29019
rect 1719 28985 1728 29019
rect 1676 28976 1728 28985
rect 6920 29121 6929 29155
rect 6929 29121 6963 29155
rect 6963 29121 6972 29155
rect 8300 29155 8352 29164
rect 6920 29112 6972 29121
rect 8300 29121 8309 29155
rect 8309 29121 8343 29155
rect 8343 29121 8352 29155
rect 8300 29112 8352 29121
rect 7012 29087 7064 29096
rect 7012 29053 7021 29087
rect 7021 29053 7055 29087
rect 7055 29053 7064 29087
rect 7012 29044 7064 29053
rect 7840 29044 7892 29096
rect 57520 29180 57572 29232
rect 59360 29180 59412 29232
rect 57888 29112 57940 29164
rect 9220 29087 9272 29096
rect 9220 29053 9229 29087
rect 9229 29053 9263 29087
rect 9263 29053 9272 29087
rect 9220 29044 9272 29053
rect 57244 29044 57296 29096
rect 59452 29044 59504 29096
rect 6368 28976 6420 29028
rect 7748 29019 7800 29028
rect 7748 28985 7757 29019
rect 7757 28985 7791 29019
rect 7791 28985 7800 29019
rect 7748 28976 7800 28985
rect 10232 29019 10284 29028
rect 10232 28985 10241 29019
rect 10241 28985 10275 29019
rect 10275 28985 10284 29019
rect 10232 28976 10284 28985
rect 57520 29019 57572 29028
rect 57520 28985 57529 29019
rect 57529 28985 57563 29019
rect 57563 28985 57572 29019
rect 57520 28976 57572 28985
rect 6552 28951 6604 28960
rect 6552 28917 6561 28951
rect 6561 28917 6595 28951
rect 6595 28917 6604 28951
rect 6552 28908 6604 28917
rect 10048 28908 10100 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 3608 28704 3660 28756
rect 6920 28704 6972 28756
rect 9956 28704 10008 28756
rect 10692 28568 10744 28620
rect 6552 28543 6604 28552
rect 6552 28509 6561 28543
rect 6561 28509 6595 28543
rect 6595 28509 6604 28543
rect 6552 28500 6604 28509
rect 8300 28500 8352 28552
rect 8208 28432 8260 28484
rect 57796 28704 57848 28756
rect 13728 28679 13780 28688
rect 13728 28645 13737 28679
rect 13737 28645 13771 28679
rect 13771 28645 13780 28679
rect 13728 28636 13780 28645
rect 57888 28636 57940 28688
rect 13820 28500 13872 28552
rect 58348 28543 58400 28552
rect 58348 28509 58357 28543
rect 58357 28509 58391 28543
rect 58391 28509 58400 28543
rect 58348 28500 58400 28509
rect 6460 28364 6512 28416
rect 7840 28364 7892 28416
rect 9864 28407 9916 28416
rect 9864 28373 9873 28407
rect 9873 28373 9907 28407
rect 9907 28373 9916 28407
rect 9864 28364 9916 28373
rect 10324 28407 10376 28416
rect 10324 28373 10333 28407
rect 10333 28373 10367 28407
rect 10367 28373 10376 28407
rect 10324 28364 10376 28373
rect 10876 28364 10928 28416
rect 14372 28364 14424 28416
rect 56876 28364 56928 28416
rect 57152 28364 57204 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 2412 28160 2464 28212
rect 10324 28160 10376 28212
rect 58348 28160 58400 28212
rect 9864 28067 9916 28076
rect 1676 27931 1728 27940
rect 1676 27897 1685 27931
rect 1685 27897 1719 27931
rect 1719 27897 1728 27931
rect 1676 27888 1728 27897
rect 9864 28033 9873 28067
rect 9873 28033 9907 28067
rect 9907 28033 9916 28067
rect 9864 28024 9916 28033
rect 10048 28024 10100 28076
rect 13728 28024 13780 28076
rect 58348 28067 58400 28076
rect 58348 28033 58357 28067
rect 58357 28033 58391 28067
rect 58391 28033 58400 28067
rect 58348 28024 58400 28033
rect 59820 27888 59872 27940
rect 4896 27820 4948 27872
rect 5356 27820 5408 27872
rect 8300 27820 8352 27872
rect 9772 27820 9824 27872
rect 11612 27820 11664 27872
rect 13820 27863 13872 27872
rect 13820 27829 13829 27863
rect 13829 27829 13863 27863
rect 13863 27829 13872 27863
rect 13820 27820 13872 27829
rect 15016 27820 15068 27872
rect 15568 27863 15620 27872
rect 15568 27829 15577 27863
rect 15577 27829 15611 27863
rect 15611 27829 15620 27863
rect 15568 27820 15620 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 5724 27659 5776 27668
rect 5724 27625 5733 27659
rect 5733 27625 5767 27659
rect 5767 27625 5776 27659
rect 5724 27616 5776 27625
rect 6184 27480 6236 27532
rect 5356 27455 5408 27464
rect 5356 27421 5365 27455
rect 5365 27421 5399 27455
rect 5399 27421 5408 27455
rect 5356 27412 5408 27421
rect 5448 27412 5500 27464
rect 9496 27616 9548 27668
rect 10692 27616 10744 27668
rect 8116 27548 8168 27600
rect 7656 27480 7708 27532
rect 14188 27548 14240 27600
rect 58348 27616 58400 27668
rect 58072 27548 58124 27600
rect 13360 27523 13412 27532
rect 13360 27489 13369 27523
rect 13369 27489 13403 27523
rect 13403 27489 13412 27523
rect 13360 27480 13412 27489
rect 14004 27480 14056 27532
rect 57980 27480 58032 27532
rect 59084 27480 59136 27532
rect 58348 27455 58400 27464
rect 58348 27421 58357 27455
rect 58357 27421 58391 27455
rect 58391 27421 58400 27455
rect 58348 27412 58400 27421
rect 5264 27387 5316 27396
rect 5264 27353 5273 27387
rect 5273 27353 5307 27387
rect 5307 27353 5316 27387
rect 5264 27344 5316 27353
rect 5908 27344 5960 27396
rect 7840 27344 7892 27396
rect 10600 27344 10652 27396
rect 10784 27344 10836 27396
rect 1676 27319 1728 27328
rect 1676 27285 1685 27319
rect 1685 27285 1719 27319
rect 1719 27285 1728 27319
rect 1676 27276 1728 27285
rect 1952 27276 2004 27328
rect 8760 27276 8812 27328
rect 9220 27276 9272 27328
rect 11520 27276 11572 27328
rect 12348 27276 12400 27328
rect 15016 27276 15068 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 6184 27072 6236 27124
rect 9312 27115 9364 27124
rect 3976 27004 4028 27056
rect 7840 27004 7892 27056
rect 2596 26936 2648 26988
rect 2504 26868 2556 26920
rect 5724 26936 5776 26988
rect 9312 27081 9321 27115
rect 9321 27081 9355 27115
rect 9355 27081 9364 27115
rect 9312 27072 9364 27081
rect 9220 27047 9272 27056
rect 9220 27013 9229 27047
rect 9229 27013 9263 27047
rect 9263 27013 9272 27047
rect 9220 27004 9272 27013
rect 10324 26936 10376 26988
rect 10784 26979 10836 26988
rect 10784 26945 10793 26979
rect 10793 26945 10827 26979
rect 10827 26945 10836 26979
rect 10784 26936 10836 26945
rect 12072 27072 12124 27124
rect 58348 27115 58400 27124
rect 58348 27081 58357 27115
rect 58357 27081 58391 27115
rect 58391 27081 58400 27115
rect 58348 27072 58400 27081
rect 13452 27047 13504 27056
rect 13452 27013 13461 27047
rect 13461 27013 13495 27047
rect 13495 27013 13504 27047
rect 13452 27004 13504 27013
rect 13820 27004 13872 27056
rect 15108 27004 15160 27056
rect 12348 26979 12400 26988
rect 12348 26945 12357 26979
rect 12357 26945 12391 26979
rect 12391 26945 12400 26979
rect 12348 26936 12400 26945
rect 14740 26979 14792 26988
rect 9496 26911 9548 26920
rect 9496 26877 9505 26911
rect 9505 26877 9539 26911
rect 9539 26877 9548 26911
rect 9496 26868 9548 26877
rect 10600 26911 10652 26920
rect 10600 26877 10609 26911
rect 10609 26877 10643 26911
rect 10643 26877 10652 26911
rect 10600 26868 10652 26877
rect 2872 26732 2924 26784
rect 5448 26800 5500 26852
rect 7564 26800 7616 26852
rect 11520 26868 11572 26920
rect 11980 26868 12032 26920
rect 14740 26945 14749 26979
rect 14749 26945 14783 26979
rect 14783 26945 14792 26979
rect 14740 26936 14792 26945
rect 13452 26868 13504 26920
rect 14004 26868 14056 26920
rect 15016 26868 15068 26920
rect 17500 26868 17552 26920
rect 13360 26800 13412 26852
rect 5632 26732 5684 26784
rect 5908 26775 5960 26784
rect 5908 26741 5917 26775
rect 5917 26741 5951 26775
rect 5951 26741 5960 26775
rect 5908 26732 5960 26741
rect 6828 26732 6880 26784
rect 8484 26732 8536 26784
rect 12716 26732 12768 26784
rect 12992 26775 13044 26784
rect 12992 26741 13001 26775
rect 13001 26741 13035 26775
rect 13035 26741 13044 26775
rect 12992 26732 13044 26741
rect 15752 26775 15804 26784
rect 15752 26741 15761 26775
rect 15761 26741 15795 26775
rect 15795 26741 15804 26775
rect 15752 26732 15804 26741
rect 17592 26775 17644 26784
rect 17592 26741 17601 26775
rect 17601 26741 17635 26775
rect 17635 26741 17644 26775
rect 17592 26732 17644 26741
rect 57152 26732 57204 26784
rect 57520 26775 57572 26784
rect 57520 26741 57529 26775
rect 57529 26741 57563 26775
rect 57563 26741 57572 26775
rect 57520 26732 57572 26741
rect 57796 26732 57848 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4068 26528 4120 26580
rect 1676 26503 1728 26512
rect 1676 26469 1685 26503
rect 1685 26469 1719 26503
rect 1719 26469 1728 26503
rect 1676 26460 1728 26469
rect 2136 26392 2188 26444
rect 3976 26392 4028 26444
rect 8668 26528 8720 26580
rect 9312 26528 9364 26580
rect 9956 26528 10008 26580
rect 10600 26528 10652 26580
rect 2872 26324 2924 26376
rect 4620 26324 4672 26376
rect 8208 26460 8260 26512
rect 8300 26460 8352 26512
rect 9496 26460 9548 26512
rect 12164 26460 12216 26512
rect 13268 26528 13320 26580
rect 14740 26571 14792 26580
rect 14740 26537 14749 26571
rect 14749 26537 14783 26571
rect 14783 26537 14792 26571
rect 14740 26528 14792 26537
rect 15016 26528 15068 26580
rect 13820 26460 13872 26512
rect 15108 26460 15160 26512
rect 6184 26392 6236 26444
rect 6644 26435 6696 26444
rect 6644 26401 6653 26435
rect 6653 26401 6687 26435
rect 6687 26401 6696 26435
rect 6644 26392 6696 26401
rect 6552 26324 6604 26376
rect 2044 26256 2096 26308
rect 2596 26256 2648 26308
rect 5448 26256 5500 26308
rect 5632 26256 5684 26308
rect 10416 26392 10468 26444
rect 17592 26460 17644 26512
rect 12992 26324 13044 26376
rect 13452 26324 13504 26376
rect 15476 26324 15528 26376
rect 15752 26324 15804 26376
rect 57336 26435 57388 26444
rect 16764 26324 16816 26376
rect 9128 26299 9180 26308
rect 9128 26265 9137 26299
rect 9137 26265 9171 26299
rect 9171 26265 9180 26299
rect 9128 26256 9180 26265
rect 57336 26401 57354 26435
rect 57354 26401 57388 26435
rect 57336 26392 57388 26401
rect 57980 26460 58032 26512
rect 57796 26392 57848 26444
rect 58440 26392 58492 26444
rect 57152 26367 57204 26376
rect 57152 26333 57161 26367
rect 57161 26333 57195 26367
rect 57195 26333 57204 26367
rect 57152 26324 57204 26333
rect 3700 26188 3752 26240
rect 6736 26231 6788 26240
rect 6736 26197 6745 26231
rect 6745 26197 6779 26231
rect 6779 26197 6788 26231
rect 6736 26188 6788 26197
rect 7196 26188 7248 26240
rect 19432 26256 19484 26308
rect 58440 26256 58492 26308
rect 14096 26188 14148 26240
rect 15936 26231 15988 26240
rect 15936 26197 15945 26231
rect 15945 26197 15979 26231
rect 15979 26197 15988 26231
rect 15936 26188 15988 26197
rect 16396 26231 16448 26240
rect 16396 26197 16405 26231
rect 16405 26197 16439 26231
rect 16439 26197 16448 26231
rect 16396 26188 16448 26197
rect 17040 26188 17092 26240
rect 17500 26231 17552 26240
rect 17500 26197 17509 26231
rect 17509 26197 17543 26231
rect 17543 26197 17552 26231
rect 44364 26231 44416 26240
rect 17500 26188 17552 26197
rect 44364 26197 44373 26231
rect 44373 26197 44407 26231
rect 44407 26197 44416 26231
rect 44364 26188 44416 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 2780 25984 2832 26036
rect 1860 25916 1912 25968
rect 9128 25916 9180 25968
rect 1768 25848 1820 25900
rect 3700 25891 3752 25900
rect 3700 25857 3709 25891
rect 3709 25857 3743 25891
rect 3743 25857 3752 25891
rect 3700 25848 3752 25857
rect 3976 25848 4028 25900
rect 7196 25891 7248 25900
rect 7196 25857 7205 25891
rect 7205 25857 7239 25891
rect 7239 25857 7248 25891
rect 7196 25848 7248 25857
rect 2136 25823 2188 25832
rect 2136 25789 2145 25823
rect 2145 25789 2179 25823
rect 2179 25789 2188 25823
rect 2136 25780 2188 25789
rect 2320 25823 2372 25832
rect 2320 25789 2329 25823
rect 2329 25789 2363 25823
rect 2363 25789 2372 25823
rect 2320 25780 2372 25789
rect 2688 25780 2740 25832
rect 3332 25780 3384 25832
rect 8392 25848 8444 25900
rect 6552 25712 6604 25764
rect 8300 25780 8352 25832
rect 2412 25644 2464 25696
rect 3884 25687 3936 25696
rect 3884 25653 3893 25687
rect 3893 25653 3927 25687
rect 3927 25653 3936 25687
rect 3884 25644 3936 25653
rect 9312 25712 9364 25764
rect 15384 25984 15436 26036
rect 16396 25984 16448 26036
rect 56048 25984 56100 26036
rect 58808 25984 58860 26036
rect 10324 25848 10376 25900
rect 10600 25891 10652 25900
rect 10600 25857 10609 25891
rect 10609 25857 10643 25891
rect 10643 25857 10652 25891
rect 10600 25848 10652 25857
rect 10692 25823 10744 25832
rect 10692 25789 10701 25823
rect 10701 25789 10735 25823
rect 10735 25789 10744 25823
rect 10692 25780 10744 25789
rect 15476 25848 15528 25900
rect 15936 25848 15988 25900
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 57520 25891 57572 25900
rect 57520 25857 57529 25891
rect 57529 25857 57563 25891
rect 57563 25857 57572 25891
rect 57520 25848 57572 25857
rect 58348 25891 58400 25900
rect 58348 25857 58357 25891
rect 58357 25857 58391 25891
rect 58391 25857 58400 25891
rect 58348 25848 58400 25857
rect 14280 25823 14332 25832
rect 14280 25789 14289 25823
rect 14289 25789 14323 25823
rect 14323 25789 14332 25823
rect 14280 25780 14332 25789
rect 14464 25823 14516 25832
rect 14464 25789 14473 25823
rect 14473 25789 14507 25823
rect 14507 25789 14516 25823
rect 14464 25780 14516 25789
rect 14004 25712 14056 25764
rect 9128 25644 9180 25696
rect 9404 25644 9456 25696
rect 13176 25687 13228 25696
rect 13176 25653 13185 25687
rect 13185 25653 13219 25687
rect 13219 25653 13228 25687
rect 13176 25644 13228 25653
rect 15384 25687 15436 25696
rect 15384 25653 15393 25687
rect 15393 25653 15427 25687
rect 15427 25653 15436 25687
rect 15384 25644 15436 25653
rect 15936 25644 15988 25696
rect 17500 25644 17552 25696
rect 19248 25644 19300 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1676 25483 1728 25492
rect 1676 25449 1685 25483
rect 1685 25449 1719 25483
rect 1719 25449 1728 25483
rect 1676 25440 1728 25449
rect 3148 25483 3200 25492
rect 3148 25449 3157 25483
rect 3157 25449 3191 25483
rect 3191 25449 3200 25483
rect 3148 25440 3200 25449
rect 5356 25440 5408 25492
rect 6736 25440 6788 25492
rect 8392 25440 8444 25492
rect 10692 25440 10744 25492
rect 14464 25483 14516 25492
rect 14464 25449 14473 25483
rect 14473 25449 14507 25483
rect 14507 25449 14516 25483
rect 14464 25440 14516 25449
rect 5540 25372 5592 25424
rect 3240 25304 3292 25356
rect 15292 25372 15344 25424
rect 2228 25236 2280 25288
rect 2412 25279 2464 25288
rect 2412 25245 2421 25279
rect 2421 25245 2455 25279
rect 2455 25245 2464 25279
rect 2412 25236 2464 25245
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 57336 25347 57388 25356
rect 57336 25313 57354 25347
rect 57354 25313 57388 25347
rect 57336 25304 57388 25313
rect 58900 25372 58952 25424
rect 57796 25304 57848 25356
rect 58256 25304 58308 25356
rect 57152 25279 57204 25288
rect 57152 25245 57161 25279
rect 57161 25245 57195 25279
rect 57195 25245 57204 25279
rect 58164 25279 58216 25288
rect 57152 25236 57204 25245
rect 58164 25245 58173 25279
rect 58173 25245 58207 25279
rect 58207 25245 58216 25279
rect 58164 25236 58216 25245
rect 17408 25168 17460 25220
rect 1768 25100 1820 25152
rect 3148 25100 3200 25152
rect 10324 25100 10376 25152
rect 14280 25100 14332 25152
rect 15476 25100 15528 25152
rect 16764 25143 16816 25152
rect 16764 25109 16773 25143
rect 16773 25109 16807 25143
rect 16807 25109 16816 25143
rect 16764 25100 16816 25109
rect 57980 25100 58032 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 2412 24760 2464 24812
rect 58348 24803 58400 24812
rect 58348 24769 58357 24803
rect 58357 24769 58391 24803
rect 58391 24769 58400 24803
rect 58348 24760 58400 24769
rect 2136 24692 2188 24744
rect 2596 24692 2648 24744
rect 1676 24667 1728 24676
rect 1676 24633 1685 24667
rect 1685 24633 1719 24667
rect 1719 24633 1728 24667
rect 1676 24624 1728 24633
rect 56692 24624 56744 24676
rect 57796 24624 57848 24676
rect 58624 24624 58676 24676
rect 2228 24556 2280 24608
rect 3516 24599 3568 24608
rect 3516 24565 3525 24599
rect 3525 24565 3559 24599
rect 3559 24565 3568 24599
rect 3516 24556 3568 24565
rect 14280 24556 14332 24608
rect 14648 24556 14700 24608
rect 57152 24556 57204 24608
rect 57336 24556 57388 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2596 24352 2648 24404
rect 19432 24352 19484 24404
rect 58348 24352 58400 24404
rect 57244 24284 57296 24336
rect 3516 24148 3568 24200
rect 58348 24191 58400 24200
rect 58348 24157 58357 24191
rect 58357 24157 58391 24191
rect 58391 24157 58400 24191
rect 58348 24148 58400 24157
rect 6368 24080 6420 24132
rect 18604 24080 18656 24132
rect 1676 24055 1728 24064
rect 1676 24021 1685 24055
rect 1685 24021 1719 24055
rect 1719 24021 1728 24055
rect 1676 24012 1728 24021
rect 2412 24055 2464 24064
rect 2412 24021 2421 24055
rect 2421 24021 2455 24055
rect 2455 24021 2464 24055
rect 2412 24012 2464 24021
rect 20444 24055 20496 24064
rect 20444 24021 20453 24055
rect 20453 24021 20487 24055
rect 20487 24021 20496 24055
rect 20444 24012 20496 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 2412 23808 2464 23860
rect 18420 23808 18472 23860
rect 58900 23808 58952 23860
rect 3332 23740 3384 23792
rect 5080 23740 5132 23792
rect 5540 23783 5592 23792
rect 5540 23749 5549 23783
rect 5549 23749 5583 23783
rect 5583 23749 5592 23783
rect 5540 23740 5592 23749
rect 8944 23740 8996 23792
rect 9312 23740 9364 23792
rect 6644 23672 6696 23724
rect 2136 23647 2188 23656
rect 2136 23613 2145 23647
rect 2145 23613 2179 23647
rect 2179 23613 2188 23647
rect 2136 23604 2188 23613
rect 2412 23604 2464 23656
rect 2596 23604 2648 23656
rect 2688 23604 2740 23656
rect 6644 23536 6696 23588
rect 2320 23468 2372 23520
rect 10140 23604 10192 23656
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4068 23264 4120 23316
rect 10232 23264 10284 23316
rect 2596 23196 2648 23248
rect 6644 23171 6696 23180
rect 6644 23137 6653 23171
rect 6653 23137 6687 23171
rect 6687 23137 6696 23171
rect 6644 23128 6696 23137
rect 11612 23128 11664 23180
rect 57980 23128 58032 23180
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 2688 23060 2740 23112
rect 12440 23103 12492 23112
rect 12440 23069 12449 23103
rect 12449 23069 12483 23103
rect 12483 23069 12492 23103
rect 12440 23060 12492 23069
rect 53104 23060 53156 23112
rect 5356 22992 5408 23044
rect 11888 22992 11940 23044
rect 1676 22967 1728 22976
rect 1676 22933 1685 22967
rect 1685 22933 1719 22967
rect 1719 22933 1728 22967
rect 1676 22924 1728 22933
rect 3148 22967 3200 22976
rect 3148 22933 3157 22967
rect 3157 22933 3191 22967
rect 3191 22933 3200 22967
rect 3148 22924 3200 22933
rect 4068 22967 4120 22976
rect 4068 22933 4077 22967
rect 4077 22933 4111 22967
rect 4111 22933 4120 22967
rect 4068 22924 4120 22933
rect 10600 22924 10652 22976
rect 18420 22967 18472 22976
rect 18420 22933 18429 22967
rect 18429 22933 18463 22967
rect 18463 22933 18472 22967
rect 18420 22924 18472 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2504 22720 2556 22772
rect 2688 22763 2740 22772
rect 2688 22729 2697 22763
rect 2697 22729 2731 22763
rect 2731 22729 2740 22763
rect 2688 22720 2740 22729
rect 3240 22763 3292 22772
rect 3240 22729 3249 22763
rect 3249 22729 3283 22763
rect 3283 22729 3292 22763
rect 3240 22720 3292 22729
rect 8576 22720 8628 22772
rect 11704 22720 11756 22772
rect 11888 22720 11940 22772
rect 14188 22763 14240 22772
rect 2136 22559 2188 22568
rect 2136 22525 2145 22559
rect 2145 22525 2179 22559
rect 2179 22525 2188 22559
rect 2136 22516 2188 22525
rect 5080 22652 5132 22704
rect 5356 22652 5408 22704
rect 12716 22695 12768 22704
rect 12716 22661 12725 22695
rect 12725 22661 12759 22695
rect 12759 22661 12768 22695
rect 12716 22652 12768 22661
rect 14188 22729 14197 22763
rect 14197 22729 14231 22763
rect 14231 22729 14240 22763
rect 14188 22720 14240 22729
rect 10140 22627 10192 22636
rect 10140 22593 10149 22627
rect 10149 22593 10183 22627
rect 10183 22593 10192 22627
rect 12440 22627 12492 22636
rect 10140 22584 10192 22593
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 13820 22584 13872 22636
rect 56784 22720 56836 22772
rect 19248 22652 19300 22704
rect 58348 22627 58400 22636
rect 58348 22593 58357 22627
rect 58357 22593 58391 22627
rect 58391 22593 58400 22627
rect 58348 22584 58400 22593
rect 3332 22516 3384 22568
rect 8208 22516 8260 22568
rect 18420 22516 18472 22568
rect 17408 22448 17460 22500
rect 15660 22380 15712 22432
rect 20352 22380 20404 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1676 22219 1728 22228
rect 1676 22185 1685 22219
rect 1685 22185 1719 22219
rect 1719 22185 1728 22219
rect 1676 22176 1728 22185
rect 3148 22176 3200 22228
rect 15936 22176 15988 22228
rect 2136 22040 2188 22092
rect 16764 22083 16816 22092
rect 16764 22049 16773 22083
rect 16773 22049 16807 22083
rect 16807 22049 16816 22083
rect 16764 22040 16816 22049
rect 1860 22015 1912 22024
rect 1860 21981 1869 22015
rect 1869 21981 1903 22015
rect 1903 21981 1912 22015
rect 1860 21972 1912 21981
rect 2504 21836 2556 21888
rect 5264 21904 5316 21956
rect 6000 21904 6052 21956
rect 6644 21972 6696 22024
rect 58348 22015 58400 22024
rect 58348 21981 58357 22015
rect 58357 21981 58391 22015
rect 58391 21981 58400 22015
rect 58348 21972 58400 21981
rect 15200 21904 15252 21956
rect 16028 21904 16080 21956
rect 19248 21836 19300 21888
rect 58716 21836 58768 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 2872 21632 2924 21684
rect 16212 21632 16264 21684
rect 58164 21675 58216 21684
rect 58164 21641 58173 21675
rect 58173 21641 58207 21675
rect 58207 21641 58216 21675
rect 58164 21632 58216 21641
rect 13820 21564 13872 21616
rect 15200 21564 15252 21616
rect 2596 21496 2648 21548
rect 17592 21564 17644 21616
rect 20168 21496 20220 21548
rect 58348 21539 58400 21548
rect 58348 21505 58357 21539
rect 58357 21505 58391 21539
rect 58391 21505 58400 21539
rect 58348 21496 58400 21505
rect 11796 21428 11848 21480
rect 13820 21428 13872 21480
rect 15292 21471 15344 21480
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 1676 21403 1728 21412
rect 1676 21369 1685 21403
rect 1685 21369 1719 21403
rect 1719 21369 1728 21403
rect 1676 21360 1728 21369
rect 2780 21292 2832 21344
rect 2964 21292 3016 21344
rect 14096 21292 14148 21344
rect 20168 21335 20220 21344
rect 20168 21301 20177 21335
rect 20177 21301 20211 21335
rect 20211 21301 20220 21335
rect 20168 21292 20220 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 11980 21131 12032 21140
rect 11980 21097 11989 21131
rect 11989 21097 12023 21131
rect 12023 21097 12032 21131
rect 11980 21088 12032 21097
rect 14372 21088 14424 21140
rect 18236 21131 18288 21140
rect 18236 21097 18245 21131
rect 18245 21097 18279 21131
rect 18279 21097 18288 21131
rect 18236 21088 18288 21097
rect 2964 20952 3016 21004
rect 12440 20952 12492 21004
rect 15200 20952 15252 21004
rect 15568 20995 15620 21004
rect 15568 20961 15577 20995
rect 15577 20961 15611 20995
rect 15611 20961 15620 20995
rect 15568 20952 15620 20961
rect 58256 21088 58308 21140
rect 20168 20952 20220 21004
rect 20628 20952 20680 21004
rect 3056 20884 3108 20936
rect 12348 20884 12400 20936
rect 19432 20884 19484 20936
rect 58348 20927 58400 20936
rect 58348 20893 58357 20927
rect 58357 20893 58391 20927
rect 58391 20893 58400 20927
rect 58348 20884 58400 20893
rect 1860 20816 1912 20868
rect 4160 20816 4212 20868
rect 13360 20816 13412 20868
rect 16028 20816 16080 20868
rect 2688 20791 2740 20800
rect 2688 20757 2697 20791
rect 2697 20757 2731 20791
rect 2731 20757 2740 20791
rect 2688 20748 2740 20757
rect 3056 20748 3108 20800
rect 3424 20748 3476 20800
rect 3792 20748 3844 20800
rect 4804 20748 4856 20800
rect 10784 20748 10836 20800
rect 19340 20748 19392 20800
rect 20628 20791 20680 20800
rect 20628 20757 20637 20791
rect 20637 20757 20671 20791
rect 20671 20757 20680 20791
rect 20628 20748 20680 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 1676 20587 1728 20596
rect 1676 20553 1685 20587
rect 1685 20553 1719 20587
rect 1719 20553 1728 20587
rect 1676 20544 1728 20553
rect 4712 20544 4764 20596
rect 10876 20587 10928 20596
rect 10876 20553 10885 20587
rect 10885 20553 10919 20587
rect 10919 20553 10928 20587
rect 10876 20544 10928 20553
rect 11612 20544 11664 20596
rect 14924 20544 14976 20596
rect 18788 20544 18840 20596
rect 5264 20476 5316 20528
rect 8944 20476 8996 20528
rect 2136 20408 2188 20460
rect 2688 20408 2740 20460
rect 19340 20408 19392 20460
rect 19524 20451 19576 20460
rect 19524 20417 19533 20451
rect 19533 20417 19567 20451
rect 19567 20417 19576 20451
rect 19524 20408 19576 20417
rect 3884 20340 3936 20392
rect 6000 20383 6052 20392
rect 6000 20349 6009 20383
rect 6009 20349 6043 20383
rect 6043 20349 6052 20383
rect 6000 20340 6052 20349
rect 8300 20340 8352 20392
rect 9772 20340 9824 20392
rect 4712 20272 4764 20324
rect 16028 20204 16080 20256
rect 19984 20204 20036 20256
rect 20444 20247 20496 20256
rect 20444 20213 20453 20247
rect 20453 20213 20487 20247
rect 20487 20213 20496 20247
rect 20444 20204 20496 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 18420 20000 18472 20052
rect 18788 20043 18840 20052
rect 18788 20009 18797 20043
rect 18797 20009 18831 20043
rect 18831 20009 18840 20043
rect 18788 20000 18840 20009
rect 15200 19864 15252 19916
rect 15660 19907 15712 19916
rect 15660 19873 15669 19907
rect 15669 19873 15703 19907
rect 15703 19873 15712 19907
rect 15660 19864 15712 19873
rect 2044 19796 2096 19848
rect 58348 19839 58400 19848
rect 58348 19805 58357 19839
rect 58357 19805 58391 19839
rect 58391 19805 58400 19839
rect 58348 19796 58400 19805
rect 5724 19771 5776 19780
rect 5724 19737 5733 19771
rect 5733 19737 5767 19771
rect 5767 19737 5776 19771
rect 5724 19728 5776 19737
rect 16120 19728 16172 19780
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 5264 19660 5316 19712
rect 19524 19703 19576 19712
rect 19524 19669 19533 19703
rect 19533 19669 19567 19703
rect 19567 19669 19576 19703
rect 19524 19660 19576 19669
rect 20536 19660 20588 19712
rect 58072 19660 58124 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4160 19456 4212 19508
rect 8760 19456 8812 19508
rect 14648 19499 14700 19508
rect 14648 19465 14657 19499
rect 14657 19465 14691 19499
rect 14691 19465 14700 19499
rect 14648 19456 14700 19465
rect 56600 19456 56652 19508
rect 5264 19388 5316 19440
rect 2228 19320 2280 19372
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 8300 19388 8352 19440
rect 9036 19388 9088 19440
rect 6000 19320 6052 19329
rect 12440 19320 12492 19372
rect 12624 19320 12676 19372
rect 4712 19252 4764 19304
rect 8116 19252 8168 19304
rect 13176 19295 13228 19304
rect 13176 19261 13185 19295
rect 13185 19261 13219 19295
rect 13219 19261 13228 19295
rect 13176 19252 13228 19261
rect 1676 19159 1728 19168
rect 1676 19125 1685 19159
rect 1685 19125 1719 19159
rect 1719 19125 1728 19159
rect 1676 19116 1728 19125
rect 12348 19116 12400 19168
rect 16120 19388 16172 19440
rect 58348 19363 58400 19372
rect 58348 19329 58357 19363
rect 58357 19329 58391 19363
rect 58391 19329 58400 19363
rect 58348 19320 58400 19329
rect 57244 19295 57296 19304
rect 57244 19261 57253 19295
rect 57253 19261 57287 19295
rect 57287 19261 57296 19295
rect 57244 19252 57296 19261
rect 57520 19295 57572 19304
rect 57520 19261 57529 19295
rect 57529 19261 57563 19295
rect 57563 19261 57572 19295
rect 57520 19252 57572 19261
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 7656 18912 7708 18964
rect 58348 18955 58400 18964
rect 1860 18751 1912 18760
rect 1860 18717 1869 18751
rect 1869 18717 1903 18751
rect 1903 18717 1912 18751
rect 1860 18708 1912 18717
rect 2688 18708 2740 18760
rect 1676 18615 1728 18624
rect 1676 18581 1685 18615
rect 1685 18581 1719 18615
rect 1719 18581 1728 18615
rect 1676 18572 1728 18581
rect 2504 18615 2556 18624
rect 2504 18581 2513 18615
rect 2513 18581 2547 18615
rect 2547 18581 2556 18615
rect 2504 18572 2556 18581
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 58348 18921 58357 18955
rect 58357 18921 58391 18955
rect 58391 18921 58400 18955
rect 58348 18912 58400 18921
rect 12624 18819 12676 18828
rect 12624 18785 12633 18819
rect 12633 18785 12667 18819
rect 12667 18785 12676 18819
rect 12624 18776 12676 18785
rect 15108 18819 15160 18828
rect 15108 18785 15117 18819
rect 15117 18785 15151 18819
rect 15151 18785 15160 18819
rect 15108 18776 15160 18785
rect 17132 18819 17184 18828
rect 17132 18785 17141 18819
rect 17141 18785 17175 18819
rect 17175 18785 17184 18819
rect 17132 18776 17184 18785
rect 19984 18708 20036 18760
rect 20260 18708 20312 18760
rect 12256 18640 12308 18692
rect 15292 18640 15344 18692
rect 16120 18640 16172 18692
rect 21180 18640 21232 18692
rect 19984 18572 20036 18624
rect 45836 18572 45888 18624
rect 57244 18572 57296 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 1952 18368 2004 18420
rect 2688 18411 2740 18420
rect 2688 18377 2697 18411
rect 2697 18377 2731 18411
rect 2731 18377 2740 18411
rect 2688 18368 2740 18377
rect 5908 18368 5960 18420
rect 12256 18368 12308 18420
rect 17132 18368 17184 18420
rect 20260 18411 20312 18420
rect 20260 18377 20269 18411
rect 20269 18377 20303 18411
rect 20303 18377 20312 18411
rect 20260 18368 20312 18377
rect 9036 18300 9088 18352
rect 15108 18300 15160 18352
rect 15292 18300 15344 18352
rect 21456 18300 21508 18352
rect 2964 18232 3016 18284
rect 11060 18232 11112 18284
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 20168 18232 20220 18284
rect 58348 18275 58400 18284
rect 58348 18241 58357 18275
rect 58357 18241 58391 18275
rect 58391 18241 58400 18275
rect 58348 18232 58400 18241
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 2504 18164 2556 18216
rect 6184 18164 6236 18216
rect 6828 18164 6880 18216
rect 9220 18207 9272 18216
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 11060 18071 11112 18080
rect 11060 18037 11069 18071
rect 11069 18037 11103 18071
rect 11103 18037 11112 18071
rect 11060 18028 11112 18037
rect 20444 18028 20496 18080
rect 57428 18028 57480 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 15384 17824 15436 17876
rect 18236 17824 18288 17876
rect 21456 17867 21508 17876
rect 21456 17833 21465 17867
rect 21465 17833 21499 17867
rect 21499 17833 21508 17867
rect 21456 17824 21508 17833
rect 2964 17756 3016 17808
rect 2136 17688 2188 17740
rect 2412 17688 2464 17740
rect 14004 17688 14056 17740
rect 16028 17688 16080 17740
rect 1768 17552 1820 17604
rect 2136 17552 2188 17604
rect 2688 17527 2740 17536
rect 2688 17493 2697 17527
rect 2697 17493 2731 17527
rect 2731 17493 2740 17527
rect 2688 17484 2740 17493
rect 3332 17620 3384 17672
rect 15200 17620 15252 17672
rect 11704 17552 11756 17604
rect 16672 17552 16724 17604
rect 20168 17552 20220 17604
rect 3976 17484 4028 17536
rect 19432 17484 19484 17536
rect 20076 17527 20128 17536
rect 20076 17493 20085 17527
rect 20085 17493 20119 17527
rect 20119 17493 20128 17527
rect 20076 17484 20128 17493
rect 21640 17663 21692 17672
rect 21640 17629 21649 17663
rect 21649 17629 21683 17663
rect 21683 17629 21692 17663
rect 21640 17620 21692 17629
rect 58348 17663 58400 17672
rect 58348 17629 58357 17663
rect 58357 17629 58391 17663
rect 58391 17629 58400 17663
rect 58348 17620 58400 17629
rect 20628 17484 20680 17536
rect 23480 17484 23532 17536
rect 58716 17484 58768 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 19340 17280 19392 17332
rect 20076 17280 20128 17332
rect 4896 17212 4948 17264
rect 16304 17212 16356 17264
rect 2228 17144 2280 17196
rect 2688 17144 2740 17196
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 2964 16983 3016 16992
rect 2964 16949 2973 16983
rect 2973 16949 3007 16983
rect 3007 16949 3016 16983
rect 2964 16940 3016 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 21180 16779 21232 16788
rect 21180 16745 21189 16779
rect 21189 16745 21223 16779
rect 21223 16745 21232 16779
rect 21180 16736 21232 16745
rect 21640 16736 21692 16788
rect 2504 16600 2556 16652
rect 9128 16643 9180 16652
rect 9128 16609 9137 16643
rect 9137 16609 9171 16643
rect 9171 16609 9180 16643
rect 9128 16600 9180 16609
rect 9404 16643 9456 16652
rect 9404 16609 9413 16643
rect 9413 16609 9447 16643
rect 9447 16609 9456 16643
rect 9404 16600 9456 16609
rect 1584 16532 1636 16584
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 16948 16532 17000 16584
rect 19340 16532 19392 16584
rect 19432 16532 19484 16584
rect 20352 16532 20404 16584
rect 20444 16532 20496 16584
rect 21180 16600 21232 16652
rect 58348 16575 58400 16584
rect 58348 16541 58357 16575
rect 58357 16541 58391 16575
rect 58391 16541 58400 16575
rect 58348 16532 58400 16541
rect 5356 16464 5408 16516
rect 9036 16464 9088 16516
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 2412 16396 2464 16448
rect 10692 16396 10744 16448
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 22284 16396 22336 16448
rect 56784 16396 56836 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 9128 16192 9180 16244
rect 3332 16056 3384 16108
rect 9588 16099 9640 16108
rect 9588 16065 9597 16099
rect 9597 16065 9631 16099
rect 9631 16065 9640 16099
rect 12992 16099 13044 16108
rect 9588 16056 9640 16065
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 58348 16099 58400 16108
rect 58348 16065 58357 16099
rect 58357 16065 58391 16099
rect 58391 16065 58400 16099
rect 58348 16056 58400 16065
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2964 15852 3016 15904
rect 3332 15895 3384 15904
rect 3332 15861 3341 15895
rect 3341 15861 3375 15895
rect 3375 15861 3384 15895
rect 3332 15852 3384 15861
rect 12532 15852 12584 15904
rect 15200 15852 15252 15904
rect 15384 15852 15436 15904
rect 57796 15852 57848 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2044 15648 2096 15700
rect 3240 15691 3292 15700
rect 3240 15657 3249 15691
rect 3249 15657 3283 15691
rect 3283 15657 3292 15691
rect 3240 15648 3292 15657
rect 10416 15648 10468 15700
rect 16948 15648 17000 15700
rect 58348 15691 58400 15700
rect 58348 15657 58357 15691
rect 58357 15657 58391 15691
rect 58391 15657 58400 15691
rect 58348 15648 58400 15657
rect 4252 15512 4304 15564
rect 6184 15512 6236 15564
rect 6828 15512 6880 15564
rect 15384 15555 15436 15564
rect 15384 15521 15393 15555
rect 15393 15521 15427 15555
rect 15427 15521 15436 15555
rect 15384 15512 15436 15521
rect 19432 15512 19484 15564
rect 2964 15444 3016 15496
rect 12532 15444 12584 15496
rect 3240 15376 3292 15428
rect 5356 15376 5408 15428
rect 9036 15376 9088 15428
rect 11704 15376 11756 15428
rect 12072 15376 12124 15428
rect 16672 15376 16724 15428
rect 2688 15351 2740 15360
rect 2688 15317 2697 15351
rect 2697 15317 2731 15351
rect 2731 15317 2740 15351
rect 2688 15308 2740 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4252 15104 4304 15156
rect 5356 15104 5408 15156
rect 6552 15147 6604 15156
rect 5724 15036 5776 15088
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 7748 15104 7800 15156
rect 6460 15036 6512 15088
rect 9036 15036 9088 15088
rect 2688 14968 2740 15020
rect 6920 14968 6972 15020
rect 20168 15011 20220 15020
rect 20168 14977 20177 15011
rect 20177 14977 20211 15011
rect 20211 14977 20220 15011
rect 20168 14968 20220 14977
rect 58348 15011 58400 15020
rect 58348 14977 58357 15011
rect 58357 14977 58391 15011
rect 58391 14977 58400 15011
rect 58348 14968 58400 14977
rect 8944 14900 8996 14952
rect 1676 14875 1728 14884
rect 1676 14841 1685 14875
rect 1685 14841 1719 14875
rect 1719 14841 1728 14875
rect 1676 14832 1728 14841
rect 20444 14943 20496 14952
rect 20444 14909 20453 14943
rect 20453 14909 20487 14943
rect 20487 14909 20496 14943
rect 20444 14900 20496 14909
rect 6552 14764 6604 14816
rect 11060 14764 11112 14816
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 20076 14764 20128 14816
rect 57336 14764 57388 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2964 14424 3016 14476
rect 13268 14560 13320 14612
rect 13820 14560 13872 14612
rect 22100 14560 22152 14612
rect 19432 14492 19484 14544
rect 12164 14424 12216 14476
rect 12532 14467 12584 14476
rect 12532 14433 12541 14467
rect 12541 14433 12575 14467
rect 12575 14433 12584 14467
rect 12532 14424 12584 14433
rect 15384 14424 15436 14476
rect 18788 14424 18840 14476
rect 20352 14424 20404 14476
rect 20536 14467 20588 14476
rect 20536 14433 20545 14467
rect 20545 14433 20579 14467
rect 20579 14433 20588 14467
rect 20536 14424 20588 14433
rect 19984 14356 20036 14408
rect 22192 14356 22244 14408
rect 58348 14399 58400 14408
rect 58348 14365 58357 14399
rect 58357 14365 58391 14399
rect 58391 14365 58400 14399
rect 58348 14356 58400 14365
rect 1768 14288 1820 14340
rect 2136 14288 2188 14340
rect 11704 14288 11756 14340
rect 16672 14288 16724 14340
rect 2228 14263 2280 14272
rect 2228 14229 2237 14263
rect 2237 14229 2271 14263
rect 2271 14229 2280 14263
rect 2228 14220 2280 14229
rect 2688 14263 2740 14272
rect 2688 14229 2697 14263
rect 2697 14229 2731 14263
rect 2731 14229 2740 14263
rect 2688 14220 2740 14229
rect 18788 14263 18840 14272
rect 18788 14229 18797 14263
rect 18797 14229 18831 14263
rect 18831 14229 18840 14263
rect 18788 14220 18840 14229
rect 19984 14220 20036 14272
rect 20536 14220 20588 14272
rect 57980 14220 58032 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 1676 14059 1728 14068
rect 1676 14025 1685 14059
rect 1685 14025 1719 14059
rect 1719 14025 1728 14059
rect 1676 14016 1728 14025
rect 3884 14016 3936 14068
rect 11060 14059 11112 14068
rect 11060 14025 11069 14059
rect 11069 14025 11103 14059
rect 11103 14025 11112 14059
rect 11060 14016 11112 14025
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 2688 13880 2740 13932
rect 11704 13991 11756 14000
rect 11704 13957 11713 13991
rect 11713 13957 11747 13991
rect 11747 13957 11756 13991
rect 11704 13948 11756 13957
rect 15384 13948 15436 14000
rect 18052 14016 18104 14068
rect 22192 14059 22244 14068
rect 22192 14025 22201 14059
rect 22201 14025 22235 14059
rect 22235 14025 22244 14059
rect 22192 14016 22244 14025
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 23480 14016 23532 14025
rect 12072 13923 12124 13932
rect 12072 13889 12081 13923
rect 12081 13889 12115 13923
rect 12115 13889 12124 13923
rect 12072 13880 12124 13889
rect 16672 13948 16724 14000
rect 56692 13948 56744 14000
rect 56876 13948 56928 14000
rect 57704 13948 57756 14000
rect 20076 13880 20128 13932
rect 20536 13880 20588 13932
rect 22284 13880 22336 13932
rect 2412 13812 2464 13864
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 6276 13812 6328 13864
rect 11704 13812 11756 13864
rect 22100 13812 22152 13864
rect 56048 13855 56100 13864
rect 19432 13744 19484 13796
rect 56048 13821 56057 13855
rect 56057 13821 56091 13855
rect 56091 13821 56100 13855
rect 56048 13812 56100 13821
rect 23480 13744 23532 13796
rect 11704 13676 11756 13728
rect 22560 13676 22612 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 3608 13472 3660 13524
rect 16212 13515 16264 13524
rect 2228 13404 2280 13456
rect 16212 13481 16221 13515
rect 16221 13481 16255 13515
rect 16255 13481 16264 13515
rect 16212 13472 16264 13481
rect 19340 13472 19392 13524
rect 22100 13515 22152 13524
rect 22100 13481 22109 13515
rect 22109 13481 22143 13515
rect 22143 13481 22152 13515
rect 22100 13472 22152 13481
rect 22560 13515 22612 13524
rect 22560 13481 22569 13515
rect 22569 13481 22603 13515
rect 22603 13481 22612 13515
rect 22560 13472 22612 13481
rect 16672 13404 16724 13456
rect 3884 13336 3936 13388
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 18052 13336 18104 13388
rect 57152 13379 57204 13388
rect 57152 13345 57161 13379
rect 57161 13345 57195 13379
rect 57195 13345 57204 13379
rect 57152 13336 57204 13345
rect 57336 13379 57388 13388
rect 57336 13345 57354 13379
rect 57354 13345 57388 13379
rect 57336 13336 57388 13345
rect 58072 13404 58124 13456
rect 57704 13379 57756 13388
rect 57704 13345 57713 13379
rect 57713 13345 57747 13379
rect 57747 13345 57756 13379
rect 57704 13336 57756 13345
rect 58532 13336 58584 13388
rect 2044 13268 2096 13320
rect 6920 13268 6972 13320
rect 13820 13268 13872 13320
rect 2320 13200 2372 13252
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 5172 13200 5224 13252
rect 12164 13200 12216 13252
rect 13452 13243 13504 13252
rect 13452 13209 13461 13243
rect 13461 13209 13495 13243
rect 13495 13209 13504 13243
rect 13452 13200 13504 13209
rect 16672 13200 16724 13252
rect 17776 13200 17828 13252
rect 19984 13268 20036 13320
rect 58256 13268 58308 13320
rect 11060 13132 11112 13184
rect 17960 13132 18012 13184
rect 56140 13132 56192 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 9956 12928 10008 12980
rect 13452 12928 13504 12980
rect 22468 12928 22520 12980
rect 22560 12928 22612 12980
rect 23480 12928 23532 12980
rect 57152 12928 57204 12980
rect 3056 12903 3108 12912
rect 3056 12869 3065 12903
rect 3065 12869 3099 12903
rect 3099 12869 3108 12903
rect 3056 12860 3108 12869
rect 5448 12860 5500 12912
rect 8484 12860 8536 12912
rect 9036 12860 9088 12912
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 19432 12792 19484 12844
rect 20628 12792 20680 12844
rect 22744 12792 22796 12844
rect 57704 12792 57756 12844
rect 58348 12835 58400 12844
rect 58348 12801 58357 12835
rect 58357 12801 58391 12835
rect 58391 12801 58400 12835
rect 58348 12792 58400 12801
rect 2044 12724 2096 12776
rect 4804 12724 4856 12776
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 2412 12656 2464 12708
rect 16580 12724 16632 12776
rect 11060 12656 11112 12708
rect 11980 12656 12032 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 2320 12588 2372 12640
rect 3056 12588 3108 12640
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 20444 12767 20496 12776
rect 20444 12733 20453 12767
rect 20453 12733 20487 12767
rect 20487 12733 20496 12767
rect 20444 12724 20496 12733
rect 23480 12724 23532 12776
rect 19432 12588 19484 12640
rect 19800 12631 19852 12640
rect 19800 12597 19809 12631
rect 19809 12597 19843 12631
rect 19843 12597 19852 12631
rect 19800 12588 19852 12597
rect 22652 12588 22704 12640
rect 58164 12631 58216 12640
rect 58164 12597 58173 12631
rect 58173 12597 58207 12631
rect 58207 12597 58216 12631
rect 58164 12588 58216 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 14924 12384 14976 12436
rect 18788 12384 18840 12436
rect 22468 12427 22520 12436
rect 22468 12393 22477 12427
rect 22477 12393 22511 12427
rect 22511 12393 22520 12427
rect 22468 12384 22520 12393
rect 57704 12427 57756 12436
rect 57704 12393 57713 12427
rect 57713 12393 57747 12427
rect 57747 12393 57756 12427
rect 57704 12384 57756 12393
rect 1860 12180 1912 12232
rect 2964 12248 3016 12300
rect 6920 12248 6972 12300
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 17960 12248 18012 12300
rect 2320 12180 2372 12189
rect 8116 12180 8168 12232
rect 8300 12180 8352 12232
rect 5356 12112 5408 12164
rect 16212 12112 16264 12164
rect 16764 12112 16816 12164
rect 17776 12180 17828 12232
rect 19800 12223 19852 12232
rect 19800 12189 19809 12223
rect 19809 12189 19843 12223
rect 19843 12189 19852 12223
rect 19800 12180 19852 12189
rect 22652 12223 22704 12232
rect 22652 12189 22661 12223
rect 22661 12189 22695 12223
rect 22695 12189 22704 12223
rect 22652 12180 22704 12189
rect 58348 12223 58400 12232
rect 58348 12189 58357 12223
rect 58357 12189 58391 12223
rect 58391 12189 58400 12223
rect 58348 12180 58400 12189
rect 10784 12044 10836 12096
rect 13360 12044 13412 12096
rect 13452 12044 13504 12096
rect 57612 12044 57664 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 2596 11840 2648 11892
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 12164 11840 12216 11892
rect 3148 11772 3200 11824
rect 5356 11772 5408 11824
rect 9680 11772 9732 11824
rect 10784 11815 10836 11824
rect 10784 11781 10793 11815
rect 10793 11781 10827 11815
rect 10827 11781 10836 11815
rect 10784 11772 10836 11781
rect 13360 11840 13412 11892
rect 56324 11840 56376 11892
rect 57152 11840 57204 11892
rect 16672 11772 16724 11824
rect 2964 11636 3016 11688
rect 6920 11704 6972 11756
rect 16212 11704 16264 11756
rect 18144 11704 18196 11756
rect 20076 11704 20128 11756
rect 22744 11704 22796 11756
rect 56324 11747 56376 11756
rect 56324 11713 56333 11747
rect 56333 11713 56367 11747
rect 56367 11713 56376 11747
rect 56600 11747 56652 11756
rect 56324 11704 56376 11713
rect 56600 11713 56609 11747
rect 56609 11713 56643 11747
rect 56643 11713 56652 11747
rect 56600 11704 56652 11713
rect 8300 11636 8352 11688
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 13452 11679 13504 11688
rect 13452 11645 13461 11679
rect 13461 11645 13495 11679
rect 13495 11645 13504 11679
rect 13452 11636 13504 11645
rect 13820 11636 13872 11688
rect 20352 11679 20404 11688
rect 20352 11645 20361 11679
rect 20361 11645 20395 11679
rect 20395 11645 20404 11679
rect 20352 11636 20404 11645
rect 2596 11500 2648 11552
rect 19892 11500 19944 11552
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 23112 11679 23164 11688
rect 23112 11645 23121 11679
rect 23121 11645 23155 11679
rect 23155 11645 23164 11679
rect 23112 11636 23164 11645
rect 57980 11704 58032 11756
rect 58348 11747 58400 11756
rect 58348 11713 58357 11747
rect 58357 11713 58391 11747
rect 58391 11713 58400 11747
rect 58348 11704 58400 11713
rect 56876 11611 56928 11620
rect 56876 11577 56885 11611
rect 56885 11577 56919 11611
rect 56919 11577 56928 11611
rect 56876 11568 56928 11577
rect 58072 11636 58124 11688
rect 57980 11568 58032 11620
rect 21364 11500 21416 11509
rect 22560 11500 22612 11552
rect 55312 11500 55364 11552
rect 55772 11500 55824 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2964 11296 3016 11348
rect 9036 11296 9088 11348
rect 20352 11296 20404 11348
rect 57152 11339 57204 11348
rect 2596 11092 2648 11144
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 57152 11305 57161 11339
rect 57161 11305 57195 11339
rect 57195 11305 57204 11339
rect 57152 11296 57204 11305
rect 20720 11228 20772 11280
rect 56692 11228 56744 11280
rect 22192 11160 22244 11212
rect 23112 11160 23164 11212
rect 56876 11160 56928 11212
rect 22560 11135 22612 11144
rect 22560 11101 22569 11135
rect 22569 11101 22603 11135
rect 22603 11101 22612 11135
rect 22560 11092 22612 11101
rect 58440 11092 58492 11144
rect 1492 10956 1544 11008
rect 18880 10956 18932 11008
rect 21364 10956 21416 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 9588 10727 9640 10736
rect 9588 10693 9597 10727
rect 9597 10693 9631 10727
rect 9631 10693 9640 10727
rect 12992 10727 13044 10736
rect 9588 10684 9640 10693
rect 12992 10693 13001 10727
rect 13001 10693 13035 10727
rect 13035 10693 13044 10727
rect 12992 10684 13044 10693
rect 20720 10752 20772 10804
rect 57520 10795 57572 10804
rect 57520 10761 57529 10795
rect 57529 10761 57563 10795
rect 57563 10761 57572 10795
rect 57520 10752 57572 10761
rect 58348 10795 58400 10804
rect 58348 10761 58357 10795
rect 58357 10761 58391 10795
rect 58391 10761 58400 10795
rect 58348 10752 58400 10761
rect 18144 10684 18196 10736
rect 18880 10727 18932 10736
rect 18880 10693 18889 10727
rect 18889 10693 18923 10727
rect 18923 10693 18932 10727
rect 18880 10684 18932 10693
rect 20076 10616 20128 10668
rect 55312 10659 55364 10668
rect 55312 10625 55321 10659
rect 55321 10625 55355 10659
rect 55355 10625 55364 10659
rect 55312 10616 55364 10625
rect 2412 10548 2464 10600
rect 10140 10548 10192 10600
rect 13820 10548 13872 10600
rect 16764 10548 16816 10600
rect 2596 10412 2648 10464
rect 16304 10412 16356 10464
rect 20444 10591 20496 10600
rect 20444 10557 20453 10591
rect 20453 10557 20487 10591
rect 20487 10557 20496 10591
rect 20444 10548 20496 10557
rect 23388 10548 23440 10600
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 51724 10412 51776 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 16304 10251 16356 10260
rect 16304 10217 16313 10251
rect 16313 10217 16347 10251
rect 16347 10217 16356 10251
rect 16304 10208 16356 10217
rect 57980 10140 58032 10192
rect 58348 10140 58400 10192
rect 16764 10072 16816 10124
rect 23388 10072 23440 10124
rect 56876 10072 56928 10124
rect 9496 10004 9548 10056
rect 16672 10004 16724 10056
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 57980 10004 58032 10056
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 2780 9868 2832 9920
rect 22100 9979 22152 9988
rect 22100 9945 22109 9979
rect 22109 9945 22143 9979
rect 22143 9945 22152 9979
rect 22100 9936 22152 9945
rect 57060 9936 57112 9988
rect 22652 9868 22704 9920
rect 22744 9868 22796 9920
rect 50160 9868 50212 9920
rect 57336 9868 57388 9920
rect 57428 9868 57480 9920
rect 58164 9936 58216 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 2780 9596 2832 9648
rect 40868 9664 40920 9716
rect 50160 9664 50212 9716
rect 3792 9596 3844 9648
rect 55404 9596 55456 9648
rect 56232 9639 56284 9648
rect 56232 9605 56241 9639
rect 56241 9605 56275 9639
rect 56275 9605 56284 9639
rect 56232 9596 56284 9605
rect 57060 9596 57112 9648
rect 2412 9503 2464 9512
rect 2412 9469 2421 9503
rect 2421 9469 2455 9503
rect 2455 9469 2464 9503
rect 2412 9460 2464 9469
rect 11060 9528 11112 9580
rect 12072 9528 12124 9580
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 56876 9528 56928 9580
rect 57796 9528 57848 9580
rect 3424 9460 3476 9512
rect 9772 9460 9824 9512
rect 19432 9460 19484 9512
rect 5356 9392 5408 9444
rect 8760 9392 8812 9444
rect 12164 9392 12216 9444
rect 14832 9392 14884 9444
rect 14924 9392 14976 9444
rect 22100 9392 22152 9444
rect 58256 9392 58308 9444
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 3792 9324 3844 9376
rect 13728 9324 13780 9376
rect 19524 9367 19576 9376
rect 19524 9333 19533 9367
rect 19533 9333 19567 9367
rect 19567 9333 19576 9367
rect 19524 9324 19576 9333
rect 19616 9324 19668 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2412 9120 2464 9172
rect 14924 9120 14976 9172
rect 19616 9120 19668 9172
rect 2780 8984 2832 9036
rect 3424 8984 3476 9036
rect 3516 8984 3568 9036
rect 9496 8984 9548 9036
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 11244 8984 11296 9036
rect 13728 8984 13780 9036
rect 19524 8984 19576 9036
rect 23480 9120 23532 9172
rect 57796 9120 57848 9172
rect 58072 9120 58124 9172
rect 57060 9052 57112 9104
rect 23388 8984 23440 9036
rect 57796 8984 57848 9036
rect 3148 8916 3200 8968
rect 7380 8916 7432 8968
rect 5356 8848 5408 8900
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 3700 8780 3752 8832
rect 8300 8780 8352 8832
rect 13820 8916 13872 8968
rect 14832 8916 14884 8968
rect 22468 8916 22520 8968
rect 58348 8959 58400 8968
rect 58348 8925 58357 8959
rect 58357 8925 58391 8959
rect 58391 8925 58400 8959
rect 58348 8916 58400 8925
rect 10324 8848 10376 8900
rect 12164 8848 12216 8900
rect 14648 8848 14700 8900
rect 10508 8780 10560 8832
rect 19984 8780 20036 8832
rect 20076 8823 20128 8832
rect 20076 8789 20085 8823
rect 20085 8789 20119 8823
rect 20119 8789 20128 8823
rect 21916 8823 21968 8832
rect 20076 8780 20128 8789
rect 21916 8789 21925 8823
rect 21925 8789 21959 8823
rect 21959 8789 21968 8823
rect 21916 8780 21968 8789
rect 22560 8780 22612 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 2596 8576 2648 8628
rect 3424 8508 3476 8560
rect 8300 8551 8352 8560
rect 8300 8517 8309 8551
rect 8309 8517 8343 8551
rect 8343 8517 8352 8551
rect 8300 8508 8352 8517
rect 8760 8508 8812 8560
rect 2412 8440 2464 8492
rect 2964 8440 3016 8492
rect 7380 8372 7432 8424
rect 9496 8372 9548 8424
rect 12900 8508 12952 8560
rect 18788 8576 18840 8628
rect 19248 8576 19300 8628
rect 58348 8576 58400 8628
rect 6644 8304 6696 8356
rect 13820 8372 13872 8424
rect 14372 8372 14424 8424
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22560 8440 22612 8449
rect 58348 8483 58400 8492
rect 58348 8449 58357 8483
rect 58357 8449 58391 8483
rect 58391 8449 58400 8483
rect 58348 8440 58400 8449
rect 19432 8372 19484 8424
rect 20628 8372 20680 8424
rect 21732 8304 21784 8356
rect 57980 8304 58032 8356
rect 57428 8236 57480 8288
rect 57704 8236 57756 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 3148 8075 3200 8084
rect 3148 8041 3157 8075
rect 3157 8041 3191 8075
rect 3191 8041 3200 8075
rect 3148 8032 3200 8041
rect 3424 8032 3476 8084
rect 14648 8032 14700 8084
rect 18604 7964 18656 8016
rect 21916 7964 21968 8016
rect 2504 7896 2556 7948
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 23480 8032 23532 8084
rect 56876 7964 56928 8016
rect 57152 8007 57204 8016
rect 57152 7973 57161 8007
rect 57161 7973 57195 8007
rect 57195 7973 57204 8007
rect 57152 7964 57204 7973
rect 58716 8032 58768 8084
rect 57612 7896 57664 7948
rect 57704 7939 57756 7948
rect 57704 7905 57713 7939
rect 57713 7905 57747 7939
rect 57747 7905 57756 7939
rect 57704 7896 57756 7905
rect 2780 7828 2832 7880
rect 7380 7828 7432 7880
rect 19984 7828 20036 7880
rect 56600 7828 56652 7880
rect 56876 7828 56928 7880
rect 6644 7760 6696 7812
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 18788 7692 18840 7701
rect 21548 7735 21600 7744
rect 21548 7701 21557 7735
rect 21557 7701 21591 7735
rect 21591 7701 21600 7735
rect 21548 7692 21600 7701
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22468 7735 22520 7744
rect 22100 7692 22152 7701
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 58440 7692 58492 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 3976 7531 4028 7540
rect 3976 7497 3985 7531
rect 3985 7497 4019 7531
rect 4019 7497 4028 7531
rect 3976 7488 4028 7497
rect 18604 7531 18656 7540
rect 18604 7497 18613 7531
rect 18613 7497 18647 7531
rect 18647 7497 18656 7531
rect 18604 7488 18656 7497
rect 56600 7488 56652 7540
rect 9588 7463 9640 7472
rect 9588 7429 9597 7463
rect 9597 7429 9631 7463
rect 9631 7429 9640 7463
rect 9588 7420 9640 7429
rect 18144 7420 18196 7472
rect 56968 7463 57020 7472
rect 56968 7429 56977 7463
rect 56977 7429 57011 7463
rect 57011 7429 57020 7463
rect 56968 7420 57020 7429
rect 57704 7420 57756 7472
rect 22836 7352 22888 7404
rect 2780 7284 2832 7336
rect 4068 7284 4120 7336
rect 7380 7284 7432 7336
rect 14372 7284 14424 7336
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 21732 7284 21784 7336
rect 23388 7327 23440 7336
rect 23388 7293 23397 7327
rect 23397 7293 23431 7327
rect 23431 7293 23440 7327
rect 23388 7284 23440 7293
rect 2872 7216 2924 7268
rect 3148 7216 3200 7268
rect 3976 7216 4028 7268
rect 58348 7395 58400 7404
rect 58348 7361 58357 7395
rect 58357 7361 58391 7395
rect 58391 7361 58400 7395
rect 58348 7352 58400 7361
rect 57152 7284 57204 7336
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 19156 7191 19208 7200
rect 19156 7157 19165 7191
rect 19165 7157 19199 7191
rect 19199 7157 19208 7191
rect 19156 7148 19208 7157
rect 23112 7148 23164 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3516 6944 3568 6996
rect 23480 6987 23532 6996
rect 23480 6953 23489 6987
rect 23489 6953 23523 6987
rect 23523 6953 23532 6987
rect 23480 6944 23532 6953
rect 56324 6944 56376 6996
rect 56968 6944 57020 6996
rect 4068 6919 4120 6928
rect 4068 6885 4077 6919
rect 4077 6885 4111 6919
rect 4111 6885 4120 6919
rect 4068 6876 4120 6885
rect 57152 6876 57204 6928
rect 57336 6876 57388 6928
rect 2872 6808 2924 6860
rect 3240 6851 3292 6860
rect 3240 6817 3249 6851
rect 3249 6817 3283 6851
rect 3283 6817 3292 6851
rect 3240 6808 3292 6817
rect 10140 6808 10192 6860
rect 19156 6808 19208 6860
rect 20628 6851 20680 6860
rect 20628 6817 20637 6851
rect 20637 6817 20671 6851
rect 20671 6817 20680 6851
rect 20628 6808 20680 6817
rect 22192 6808 22244 6860
rect 56324 6851 56376 6860
rect 56324 6817 56333 6851
rect 56333 6817 56367 6851
rect 56367 6817 56376 6851
rect 56324 6808 56376 6817
rect 56784 6808 56836 6860
rect 3700 6740 3752 6792
rect 4068 6740 4120 6792
rect 7380 6740 7432 6792
rect 15476 6740 15528 6792
rect 15936 6740 15988 6792
rect 22100 6740 22152 6792
rect 22836 6740 22888 6792
rect 23112 6740 23164 6792
rect 56416 6740 56468 6792
rect 57152 6740 57204 6792
rect 58348 6783 58400 6792
rect 3516 6672 3568 6724
rect 6644 6672 6696 6724
rect 13912 6672 13964 6724
rect 21548 6672 21600 6724
rect 22468 6672 22520 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2504 6604 2556 6656
rect 15108 6604 15160 6656
rect 18144 6604 18196 6656
rect 19432 6647 19484 6656
rect 19432 6613 19441 6647
rect 19441 6613 19475 6647
rect 19475 6613 19484 6647
rect 19432 6604 19484 6613
rect 21180 6647 21232 6656
rect 21180 6613 21189 6647
rect 21189 6613 21223 6647
rect 21223 6613 21232 6647
rect 21180 6604 21232 6613
rect 22100 6647 22152 6656
rect 22100 6613 22109 6647
rect 22109 6613 22143 6647
rect 22143 6613 22152 6647
rect 22560 6647 22612 6656
rect 22100 6604 22152 6613
rect 22560 6613 22569 6647
rect 22569 6613 22603 6647
rect 22603 6613 22612 6647
rect 22560 6604 22612 6613
rect 55588 6604 55640 6656
rect 55772 6604 55824 6656
rect 56416 6604 56468 6656
rect 58348 6749 58357 6783
rect 58357 6749 58391 6783
rect 58391 6749 58400 6783
rect 58348 6740 58400 6749
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 2872 6400 2924 6452
rect 7472 6332 7524 6384
rect 22100 6400 22152 6452
rect 56968 6443 57020 6452
rect 56968 6409 56977 6443
rect 56977 6409 57011 6443
rect 57011 6409 57020 6443
rect 56968 6400 57020 6409
rect 57336 6400 57388 6452
rect 58348 6400 58400 6452
rect 9680 6332 9732 6384
rect 13912 6332 13964 6384
rect 15108 6332 15160 6384
rect 21180 6332 21232 6384
rect 2320 6264 2372 6316
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 19432 6307 19484 6316
rect 19432 6273 19441 6307
rect 19441 6273 19475 6307
rect 19475 6273 19484 6307
rect 19432 6264 19484 6273
rect 19800 6264 19852 6316
rect 22560 6307 22612 6316
rect 22560 6273 22569 6307
rect 22569 6273 22603 6307
rect 22603 6273 22612 6307
rect 22560 6264 22612 6273
rect 22836 6264 22888 6316
rect 23112 6264 23164 6316
rect 58348 6307 58400 6316
rect 58348 6273 58357 6307
rect 58357 6273 58391 6307
rect 58391 6273 58400 6307
rect 58348 6264 58400 6273
rect 9496 6196 9548 6248
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 9588 6060 9640 6112
rect 16856 6196 16908 6248
rect 18604 6196 18656 6248
rect 16948 6128 17000 6180
rect 44824 6128 44876 6180
rect 53104 6128 53156 6180
rect 56784 6128 56836 6180
rect 57336 6128 57388 6180
rect 11612 6060 11664 6112
rect 19340 6060 19392 6112
rect 22192 6060 22244 6112
rect 22652 6060 22704 6112
rect 57060 6060 57112 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1676 5899 1728 5908
rect 1676 5865 1685 5899
rect 1685 5865 1719 5899
rect 1719 5865 1728 5899
rect 1676 5856 1728 5865
rect 2688 5856 2740 5908
rect 2320 5788 2372 5840
rect 9496 5856 9548 5908
rect 16948 5856 17000 5908
rect 19800 5899 19852 5908
rect 19800 5865 19809 5899
rect 19809 5865 19843 5899
rect 19843 5865 19852 5899
rect 19800 5856 19852 5865
rect 22652 5899 22704 5908
rect 22652 5865 22661 5899
rect 22661 5865 22695 5899
rect 22695 5865 22704 5899
rect 22652 5856 22704 5865
rect 56692 5856 56744 5908
rect 57612 5856 57664 5908
rect 10140 5831 10192 5840
rect 10140 5797 10149 5831
rect 10149 5797 10183 5831
rect 10183 5797 10192 5831
rect 10140 5788 10192 5797
rect 16580 5788 16632 5840
rect 56784 5788 56836 5840
rect 57244 5788 57296 5840
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 9588 5720 9640 5772
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 20444 5763 20496 5772
rect 20444 5729 20453 5763
rect 20453 5729 20487 5763
rect 20487 5729 20496 5763
rect 20444 5720 20496 5729
rect 57060 5720 57112 5772
rect 57428 5763 57480 5772
rect 57428 5729 57437 5763
rect 57437 5729 57471 5763
rect 57471 5729 57480 5763
rect 57428 5720 57480 5729
rect 57612 5720 57664 5772
rect 2596 5652 2648 5704
rect 14372 5652 14424 5704
rect 18604 5652 18656 5704
rect 19432 5652 19484 5704
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 56692 5695 56744 5704
rect 56692 5661 56701 5695
rect 56701 5661 56735 5695
rect 56735 5661 56744 5695
rect 56692 5652 56744 5661
rect 57704 5695 57756 5704
rect 57704 5661 57713 5695
rect 57713 5661 57747 5695
rect 57747 5661 57756 5695
rect 57704 5652 57756 5661
rect 6644 5584 6696 5636
rect 9680 5584 9732 5636
rect 10324 5584 10376 5636
rect 18236 5627 18288 5636
rect 17592 5516 17644 5568
rect 18236 5593 18245 5627
rect 18245 5593 18279 5627
rect 18279 5593 18288 5627
rect 18236 5584 18288 5593
rect 18144 5516 18196 5568
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 22836 5516 22888 5568
rect 56968 5516 57020 5568
rect 57704 5516 57756 5568
rect 58256 5516 58308 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 4804 5312 4856 5364
rect 2688 5176 2740 5228
rect 1676 5083 1728 5092
rect 1676 5049 1685 5083
rect 1685 5049 1719 5083
rect 1719 5049 1728 5083
rect 1676 5040 1728 5049
rect 12900 5244 12952 5296
rect 13636 5312 13688 5364
rect 18236 5312 18288 5364
rect 20352 5312 20404 5364
rect 20536 5312 20588 5364
rect 56968 5355 57020 5364
rect 56968 5321 56977 5355
rect 56977 5321 57011 5355
rect 57011 5321 57020 5355
rect 56968 5312 57020 5321
rect 57244 5312 57296 5364
rect 58532 5312 58584 5364
rect 19340 5244 19392 5296
rect 14372 5176 14424 5228
rect 58348 5219 58400 5228
rect 58348 5185 58357 5219
rect 58357 5185 58391 5219
rect 58391 5185 58400 5219
rect 58348 5176 58400 5185
rect 20168 5108 20220 5160
rect 20444 5151 20496 5160
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 20260 4972 20312 5024
rect 22836 4972 22888 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2872 4768 2924 4820
rect 3976 4768 4028 4820
rect 16580 4768 16632 4820
rect 20168 4768 20220 4820
rect 56508 4811 56560 4820
rect 56508 4777 56517 4811
rect 56517 4777 56551 4811
rect 56551 4777 56560 4811
rect 56508 4768 56560 4777
rect 57520 4811 57572 4820
rect 57520 4777 57529 4811
rect 57529 4777 57563 4811
rect 57563 4777 57572 4811
rect 57520 4768 57572 4777
rect 58164 4811 58216 4820
rect 58164 4777 58173 4811
rect 58173 4777 58207 4811
rect 58207 4777 58216 4811
rect 58164 4768 58216 4777
rect 2504 4564 2556 4616
rect 57704 4607 57756 4616
rect 57704 4573 57713 4607
rect 57713 4573 57747 4607
rect 57747 4573 57756 4607
rect 57704 4564 57756 4573
rect 58348 4607 58400 4616
rect 58348 4573 58357 4607
rect 58357 4573 58391 4607
rect 58391 4573 58400 4607
rect 58348 4564 58400 4573
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 1676 4428 1728 4437
rect 20168 4428 20220 4480
rect 21364 4428 21416 4480
rect 23020 4428 23072 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 2412 4224 2464 4276
rect 19248 4267 19300 4276
rect 19248 4233 19257 4267
rect 19257 4233 19291 4267
rect 19291 4233 19300 4267
rect 19248 4224 19300 4233
rect 3332 4156 3384 4208
rect 2688 4020 2740 4072
rect 4712 4088 4764 4140
rect 7932 4020 7984 4072
rect 9864 4088 9916 4140
rect 19432 4088 19484 4140
rect 19524 4088 19576 4140
rect 23204 4224 23256 4276
rect 22468 4156 22520 4208
rect 24124 4088 24176 4140
rect 30012 4088 30064 4140
rect 55680 4088 55732 4140
rect 57796 4088 57848 4140
rect 16396 4020 16448 4072
rect 2872 3952 2924 4004
rect 3424 3952 3476 4004
rect 11152 3952 11204 4004
rect 16764 3952 16816 4004
rect 2412 3884 2464 3936
rect 3608 3927 3660 3936
rect 3608 3893 3617 3927
rect 3617 3893 3651 3927
rect 3651 3893 3660 3927
rect 3608 3884 3660 3893
rect 3976 3884 4028 3936
rect 7288 3884 7340 3936
rect 11060 3884 11112 3936
rect 11980 3884 12032 3936
rect 17776 3884 17828 3936
rect 20076 3952 20128 4004
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 20628 4020 20680 4072
rect 23204 4063 23256 4072
rect 23204 4029 23213 4063
rect 23213 4029 23247 4063
rect 23247 4029 23256 4063
rect 23204 4020 23256 4029
rect 23756 4020 23808 4072
rect 28908 4020 28960 4072
rect 56140 4020 56192 4072
rect 53380 3952 53432 4004
rect 19524 3884 19576 3936
rect 19708 3927 19760 3936
rect 19708 3893 19717 3927
rect 19717 3893 19751 3927
rect 19751 3893 19760 3927
rect 19708 3884 19760 3893
rect 22100 3884 22152 3936
rect 56508 3884 56560 3936
rect 58164 3884 58216 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2504 3612 2556 3664
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 8944 3680 8996 3732
rect 2872 3544 2924 3596
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 11980 3680 12032 3732
rect 14280 3680 14332 3732
rect 16396 3723 16448 3732
rect 16396 3689 16405 3723
rect 16405 3689 16439 3723
rect 16439 3689 16448 3723
rect 16396 3680 16448 3689
rect 40868 3723 40920 3732
rect 13728 3612 13780 3664
rect 2596 3476 2648 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 6920 3476 6972 3528
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 14280 3476 14332 3528
rect 1584 3408 1636 3460
rect 5080 3408 5132 3460
rect 6552 3408 6604 3460
rect 6828 3408 6880 3460
rect 9036 3408 9088 3460
rect 10324 3408 10376 3460
rect 13636 3408 13688 3460
rect 1952 3340 2004 3392
rect 2228 3340 2280 3392
rect 2964 3383 3016 3392
rect 2964 3349 2973 3383
rect 2973 3349 3007 3383
rect 3007 3349 3016 3383
rect 2964 3340 3016 3349
rect 4436 3340 4488 3392
rect 7012 3340 7064 3392
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 14740 3340 14792 3392
rect 18604 3476 18656 3528
rect 19708 3476 19760 3528
rect 20352 3544 20404 3596
rect 40868 3689 40877 3723
rect 40877 3689 40911 3723
rect 40911 3689 40920 3723
rect 40868 3680 40920 3689
rect 23204 3587 23256 3596
rect 23204 3553 23213 3587
rect 23213 3553 23247 3587
rect 23247 3553 23256 3587
rect 23204 3544 23256 3553
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 22100 3519 22152 3528
rect 22100 3485 22109 3519
rect 22109 3485 22143 3519
rect 22143 3485 22152 3519
rect 22100 3476 22152 3485
rect 40868 3476 40920 3528
rect 55956 3680 56008 3732
rect 53748 3612 53800 3664
rect 57336 3612 57388 3664
rect 55312 3544 55364 3596
rect 55588 3544 55640 3596
rect 54668 3519 54720 3528
rect 54668 3485 54677 3519
rect 54677 3485 54711 3519
rect 54711 3485 54720 3519
rect 54668 3476 54720 3485
rect 55680 3519 55732 3528
rect 55680 3485 55689 3519
rect 55689 3485 55723 3519
rect 55723 3485 55732 3519
rect 55680 3476 55732 3485
rect 56600 3476 56652 3528
rect 57428 3519 57480 3528
rect 57428 3485 57437 3519
rect 57437 3485 57471 3519
rect 57471 3485 57480 3519
rect 57428 3476 57480 3485
rect 58256 3519 58308 3528
rect 58256 3485 58265 3519
rect 58265 3485 58299 3519
rect 58299 3485 58308 3519
rect 58256 3476 58308 3485
rect 17592 3408 17644 3460
rect 18328 3340 18380 3392
rect 19984 3340 20036 3392
rect 20444 3340 20496 3392
rect 20536 3340 20588 3392
rect 23204 3408 23256 3460
rect 22376 3340 22428 3392
rect 22744 3340 22796 3392
rect 40316 3340 40368 3392
rect 48044 3340 48096 3392
rect 54484 3383 54536 3392
rect 54484 3349 54493 3383
rect 54493 3349 54527 3383
rect 54527 3349 54536 3383
rect 54484 3340 54536 3349
rect 55496 3383 55548 3392
rect 55496 3349 55505 3383
rect 55505 3349 55539 3383
rect 55539 3349 55548 3383
rect 55496 3340 55548 3349
rect 56140 3383 56192 3392
rect 56140 3349 56149 3383
rect 56149 3349 56183 3383
rect 56183 3349 56192 3383
rect 56140 3340 56192 3349
rect 56784 3383 56836 3392
rect 56784 3349 56793 3383
rect 56793 3349 56827 3383
rect 56827 3349 56836 3383
rect 56784 3340 56836 3349
rect 57980 3340 58032 3392
rect 58072 3383 58124 3392
rect 58072 3349 58081 3383
rect 58081 3349 58115 3383
rect 58115 3349 58124 3383
rect 58072 3340 58124 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 1768 3179 1820 3188
rect 1768 3145 1777 3179
rect 1777 3145 1811 3179
rect 1811 3145 1820 3179
rect 1768 3136 1820 3145
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 2596 3136 2648 3188
rect 3976 3136 4028 3188
rect 5080 3136 5132 3188
rect 13728 3136 13780 3188
rect 4436 3068 4488 3120
rect 6644 3068 6696 3120
rect 9036 3068 9088 3120
rect 9588 3068 9640 3120
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 2964 3000 3016 3052
rect 3608 3000 3660 3052
rect 2688 2932 2740 2984
rect 6920 3000 6972 3052
rect 7288 3000 7340 3052
rect 13636 3068 13688 3120
rect 23204 3179 23256 3188
rect 23204 3145 23213 3179
rect 23213 3145 23247 3179
rect 23247 3145 23256 3179
rect 23204 3136 23256 3145
rect 27252 3179 27304 3188
rect 27252 3145 27261 3179
rect 27261 3145 27295 3179
rect 27295 3145 27304 3179
rect 27252 3136 27304 3145
rect 28908 3136 28960 3188
rect 30012 3136 30064 3188
rect 30932 3179 30984 3188
rect 30932 3145 30941 3179
rect 30941 3145 30975 3179
rect 30975 3145 30984 3179
rect 30932 3136 30984 3145
rect 33324 3136 33376 3188
rect 43628 3136 43680 3188
rect 44364 3136 44416 3188
rect 44824 3179 44876 3188
rect 44824 3145 44833 3179
rect 44833 3145 44867 3179
rect 44867 3145 44876 3179
rect 44824 3136 44876 3145
rect 45836 3179 45888 3188
rect 45836 3145 45845 3179
rect 45845 3145 45879 3179
rect 45879 3145 45888 3179
rect 45836 3136 45888 3145
rect 51448 3179 51500 3188
rect 51448 3145 51457 3179
rect 51457 3145 51491 3179
rect 51491 3145 51500 3179
rect 51448 3136 51500 3145
rect 53748 3179 53800 3188
rect 53748 3145 53757 3179
rect 53757 3145 53791 3179
rect 53791 3145 53800 3179
rect 53748 3136 53800 3145
rect 54668 3136 54720 3188
rect 56692 3179 56744 3188
rect 56692 3145 56701 3179
rect 56701 3145 56735 3179
rect 56735 3145 56744 3179
rect 56692 3136 56744 3145
rect 17592 3068 17644 3120
rect 18328 3111 18380 3120
rect 18328 3077 18337 3111
rect 18337 3077 18371 3111
rect 18371 3077 18380 3111
rect 18328 3068 18380 3077
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 19340 3043 19392 3052
rect 18604 3000 18656 3009
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 21088 3000 21140 3052
rect 21364 3043 21416 3052
rect 21364 3009 21373 3043
rect 21373 3009 21407 3043
rect 21407 3009 21416 3043
rect 21364 3000 21416 3009
rect 22376 3043 22428 3052
rect 22376 3009 22385 3043
rect 22385 3009 22419 3043
rect 22419 3009 22428 3043
rect 22376 3000 22428 3009
rect 22836 3043 22888 3052
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 23020 3043 23072 3052
rect 23020 3009 23029 3043
rect 23029 3009 23063 3043
rect 23063 3009 23072 3043
rect 23020 3000 23072 3009
rect 30288 3068 30340 3120
rect 32312 3111 32364 3120
rect 32312 3077 32321 3111
rect 32321 3077 32355 3111
rect 32355 3077 32364 3111
rect 32312 3068 32364 3077
rect 37740 3068 37792 3120
rect 58072 3068 58124 3120
rect 55956 3000 56008 3052
rect 56048 3043 56100 3052
rect 56048 3009 56057 3043
rect 56057 3009 56091 3043
rect 56091 3009 56100 3043
rect 56048 3000 56100 3009
rect 56508 3000 56560 3052
rect 57336 3000 57388 3052
rect 58440 3000 58492 3052
rect 2872 2864 2924 2916
rect 18880 2932 18932 2984
rect 38660 2975 38712 2984
rect 38660 2941 38669 2975
rect 38669 2941 38703 2975
rect 38703 2941 38712 2975
rect 38660 2932 38712 2941
rect 56140 2932 56192 2984
rect 7012 2864 7064 2916
rect 16672 2864 16724 2916
rect 16764 2864 16816 2916
rect 19432 2864 19484 2916
rect 20444 2864 20496 2916
rect 39212 2864 39264 2916
rect 7840 2796 7892 2848
rect 10048 2796 10100 2848
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 12256 2796 12308 2848
rect 15568 2796 15620 2848
rect 23480 2796 23532 2848
rect 24400 2839 24452 2848
rect 24400 2805 24409 2839
rect 24409 2805 24443 2839
rect 24443 2805 24452 2839
rect 24400 2796 24452 2805
rect 25504 2839 25556 2848
rect 25504 2805 25513 2839
rect 25513 2805 25547 2839
rect 25547 2805 25556 2839
rect 25504 2796 25556 2805
rect 27712 2796 27764 2848
rect 35992 2839 36044 2848
rect 35992 2805 36001 2839
rect 36001 2805 36035 2839
rect 36035 2805 36044 2839
rect 35992 2796 36044 2805
rect 50620 2796 50672 2848
rect 54576 2796 54628 2848
rect 56048 2796 56100 2848
rect 57152 2796 57204 2848
rect 57336 2839 57388 2848
rect 57336 2805 57345 2839
rect 57345 2805 57379 2839
rect 57379 2805 57388 2839
rect 57336 2796 57388 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4712 2592 4764 2644
rect 4804 2592 4856 2644
rect 22468 2635 22520 2644
rect 22468 2601 22477 2635
rect 22477 2601 22511 2635
rect 22511 2601 22520 2635
rect 22468 2592 22520 2601
rect 22744 2592 22796 2644
rect 28632 2592 28684 2644
rect 2780 2524 2832 2576
rect 4068 2524 4120 2576
rect 15936 2567 15988 2576
rect 15936 2533 15945 2567
rect 15945 2533 15979 2567
rect 15979 2533 15988 2567
rect 15936 2524 15988 2533
rect 18788 2524 18840 2576
rect 2596 2456 2648 2508
rect 7932 2499 7984 2508
rect 7932 2465 7941 2499
rect 7941 2465 7975 2499
rect 7975 2465 7984 2499
rect 7932 2456 7984 2465
rect 10508 2456 10560 2508
rect 19156 2456 19208 2508
rect 20076 2499 20128 2508
rect 20076 2465 20085 2499
rect 20085 2465 20119 2499
rect 20119 2465 20128 2499
rect 20076 2456 20128 2465
rect 20260 2456 20312 2508
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 4528 2388 4580 2440
rect 5632 2388 5684 2440
rect 6920 2388 6972 2440
rect 8576 2388 8628 2440
rect 8944 2388 8996 2440
rect 12256 2388 12308 2440
rect 17776 2388 17828 2440
rect 7840 2320 7892 2372
rect 10048 2320 10100 2372
rect 11152 2320 11204 2372
rect 13360 2320 13412 2372
rect 14464 2320 14516 2372
rect 14740 2363 14792 2372
rect 14740 2329 14749 2363
rect 14749 2329 14783 2363
rect 14783 2329 14792 2363
rect 14740 2320 14792 2329
rect 15568 2320 15620 2372
rect 16672 2320 16724 2372
rect 22192 2320 22244 2372
rect 23480 2388 23532 2440
rect 38384 2524 38436 2576
rect 27896 2499 27948 2508
rect 27896 2465 27905 2499
rect 27905 2465 27939 2499
rect 27939 2465 27948 2499
rect 27896 2456 27948 2465
rect 28908 2431 28960 2440
rect 28908 2397 28917 2431
rect 28917 2397 28951 2431
rect 28951 2397 28960 2431
rect 28908 2388 28960 2397
rect 30012 2431 30064 2440
rect 30012 2397 30021 2431
rect 30021 2397 30055 2431
rect 30055 2397 30064 2431
rect 30012 2388 30064 2397
rect 30932 2388 30984 2440
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 33324 2431 33376 2440
rect 33324 2397 33333 2431
rect 33333 2397 33367 2431
rect 33367 2397 33376 2431
rect 33324 2388 33376 2397
rect 24400 2320 24452 2372
rect 25504 2320 25556 2372
rect 3884 2252 3936 2304
rect 4620 2252 4672 2304
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 5908 2295 5960 2304
rect 5908 2261 5917 2295
rect 5917 2261 5951 2295
rect 5951 2261 5960 2295
rect 5908 2252 5960 2261
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 13544 2295 13596 2304
rect 13544 2261 13553 2295
rect 13553 2261 13587 2295
rect 13587 2261 13596 2295
rect 13544 2252 13596 2261
rect 21364 2295 21416 2304
rect 21364 2261 21373 2295
rect 21373 2261 21407 2295
rect 21407 2261 21416 2295
rect 21364 2252 21416 2261
rect 22836 2252 22888 2304
rect 26608 2295 26660 2304
rect 26608 2261 26617 2295
rect 26617 2261 26651 2295
rect 26651 2261 26660 2295
rect 35992 2388 36044 2440
rect 37740 2431 37792 2440
rect 37740 2397 37749 2431
rect 37749 2397 37783 2431
rect 37783 2397 37792 2431
rect 37740 2388 37792 2397
rect 38660 2388 38712 2440
rect 39212 2431 39264 2440
rect 39212 2397 39221 2431
rect 39221 2397 39255 2431
rect 39255 2397 39264 2431
rect 39212 2388 39264 2397
rect 40316 2431 40368 2440
rect 40316 2397 40325 2431
rect 40325 2397 40359 2431
rect 40359 2397 40368 2431
rect 40316 2388 40368 2397
rect 36360 2363 36412 2372
rect 36360 2329 36369 2363
rect 36369 2329 36403 2363
rect 36403 2329 36412 2363
rect 36360 2320 36412 2329
rect 55680 2592 55732 2644
rect 57428 2592 57480 2644
rect 43628 2431 43680 2440
rect 43628 2397 43637 2431
rect 43637 2397 43671 2431
rect 43671 2397 43680 2431
rect 43628 2388 43680 2397
rect 44824 2388 44876 2440
rect 45836 2388 45888 2440
rect 48044 2431 48096 2440
rect 48044 2397 48053 2431
rect 48053 2397 48087 2431
rect 48087 2397 48096 2431
rect 48044 2388 48096 2397
rect 49056 2431 49108 2440
rect 49056 2397 49065 2431
rect 49065 2397 49099 2431
rect 49099 2397 49108 2431
rect 49056 2388 49108 2397
rect 50620 2431 50672 2440
rect 50620 2397 50629 2431
rect 50629 2397 50663 2431
rect 50663 2397 50672 2431
rect 50620 2388 50672 2397
rect 57336 2524 57388 2576
rect 51448 2388 51500 2440
rect 53380 2388 53432 2440
rect 54484 2388 54536 2440
rect 55496 2388 55548 2440
rect 55588 2388 55640 2440
rect 56784 2456 56836 2508
rect 55956 2388 56008 2440
rect 56416 2388 56468 2440
rect 57520 2431 57572 2440
rect 57520 2397 57529 2431
rect 57529 2397 57563 2431
rect 57563 2397 57572 2431
rect 57520 2388 57572 2397
rect 57980 2388 58032 2440
rect 55680 2320 55732 2372
rect 58164 2320 58216 2372
rect 26608 2252 26660 2261
rect 28816 2252 28868 2304
rect 29920 2252 29972 2304
rect 31024 2252 31076 2304
rect 32128 2252 32180 2304
rect 33232 2252 33284 2304
rect 34336 2295 34388 2304
rect 34336 2261 34345 2295
rect 34345 2261 34379 2295
rect 34379 2261 34388 2295
rect 34336 2252 34388 2261
rect 36544 2252 36596 2304
rect 37648 2252 37700 2304
rect 38752 2252 38804 2304
rect 39856 2252 39908 2304
rect 40960 2252 41012 2304
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 42064 2252 42116 2304
rect 43168 2252 43220 2304
rect 44272 2252 44324 2304
rect 45376 2252 45428 2304
rect 46480 2252 46532 2304
rect 47584 2252 47636 2304
rect 48688 2252 48740 2304
rect 49792 2252 49844 2304
rect 50896 2252 50948 2304
rect 52000 2252 52052 2304
rect 53104 2252 53156 2304
rect 54208 2252 54260 2304
rect 55312 2252 55364 2304
rect 56876 2252 56928 2304
rect 57520 2252 57572 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 4804 2048 4856 2100
rect 23020 2048 23072 2100
rect 36360 2048 36412 2100
rect 55404 2048 55456 2100
rect 3792 1980 3844 2032
rect 13544 1980 13596 2032
rect 41880 1980 41932 2032
rect 51724 1980 51776 2032
rect 3516 1912 3568 1964
rect 10232 1912 10284 1964
rect 5908 1844 5960 1896
rect 21364 1844 21416 1896
rect 2228 1776 2280 1828
rect 9312 1776 9364 1828
<< metal2 >>
rect 1858 59200 1914 60000
rect 3054 59200 3110 60000
rect 4250 59200 4306 60000
rect 5446 59200 5502 60000
rect 6642 59200 6698 60000
rect 7838 59200 7894 60000
rect 9034 59200 9090 60000
rect 10230 59200 10286 60000
rect 11426 59200 11482 60000
rect 12622 59200 12678 60000
rect 13818 59200 13874 60000
rect 15014 59200 15070 60000
rect 16210 59200 16266 60000
rect 17406 59200 17462 60000
rect 18602 59200 18658 60000
rect 19798 59200 19854 60000
rect 20994 59200 21050 60000
rect 22190 59200 22246 60000
rect 23386 59200 23442 60000
rect 24582 59200 24638 60000
rect 25778 59200 25834 60000
rect 26974 59200 27030 60000
rect 28170 59200 28226 60000
rect 29366 59200 29422 60000
rect 30562 59200 30618 60000
rect 31758 59200 31814 60000
rect 32954 59200 33010 60000
rect 34150 59200 34206 60000
rect 35346 59200 35402 60000
rect 36542 59200 36598 60000
rect 37738 59200 37794 60000
rect 38934 59200 38990 60000
rect 40130 59200 40186 60000
rect 41326 59200 41382 60000
rect 42522 59200 42578 60000
rect 43718 59200 43774 60000
rect 44914 59200 44970 60000
rect 46110 59200 46166 60000
rect 47306 59200 47362 60000
rect 48502 59200 48558 60000
rect 49698 59200 49754 60000
rect 50894 59200 50950 60000
rect 52090 59200 52146 60000
rect 53286 59200 53342 60000
rect 54482 59200 54538 60000
rect 55678 59200 55734 60000
rect 56874 59200 56930 60000
rect 58070 59200 58126 60000
rect 1872 57458 1900 59200
rect 2228 57860 2280 57866
rect 2228 57802 2280 57808
rect 2240 57458 2268 57802
rect 3068 57458 3096 59200
rect 4264 57458 4292 59200
rect 1860 57452 1912 57458
rect 1860 57394 1912 57400
rect 2228 57452 2280 57458
rect 2228 57394 2280 57400
rect 3056 57452 3108 57458
rect 3056 57394 3108 57400
rect 4252 57452 4304 57458
rect 4252 57394 4304 57400
rect 4620 57452 4672 57458
rect 5460 57440 5488 59200
rect 6656 57458 6684 59200
rect 7852 57458 7880 59200
rect 9048 57458 9076 59200
rect 10244 57458 10272 59200
rect 11440 57526 11468 59200
rect 11428 57520 11480 57526
rect 11428 57462 11480 57468
rect 12636 57458 12664 59200
rect 13832 57526 13860 59200
rect 13820 57520 13872 57526
rect 13820 57462 13872 57468
rect 15028 57458 15056 59200
rect 16224 57526 16252 59200
rect 16212 57520 16264 57526
rect 16212 57462 16264 57468
rect 17420 57458 17448 59200
rect 18616 57458 18644 59200
rect 19812 57848 19840 59200
rect 19812 57820 20024 57848
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 19996 57458 20024 57820
rect 21008 57458 21036 59200
rect 21640 57792 21692 57798
rect 21640 57734 21692 57740
rect 5540 57452 5592 57458
rect 5460 57412 5540 57440
rect 4620 57394 4672 57400
rect 5540 57394 5592 57400
rect 6000 57452 6052 57458
rect 6000 57394 6052 57400
rect 6644 57452 6696 57458
rect 6644 57394 6696 57400
rect 7840 57452 7892 57458
rect 7840 57394 7892 57400
rect 8484 57452 8536 57458
rect 8484 57394 8536 57400
rect 9036 57452 9088 57458
rect 9036 57394 9088 57400
rect 10232 57452 10284 57458
rect 10232 57394 10284 57400
rect 12624 57452 12676 57458
rect 12624 57394 12676 57400
rect 15016 57452 15068 57458
rect 15016 57394 15068 57400
rect 17408 57452 17460 57458
rect 17408 57394 17460 57400
rect 18604 57452 18656 57458
rect 18604 57394 18656 57400
rect 19984 57452 20036 57458
rect 19984 57394 20036 57400
rect 20996 57452 21048 57458
rect 20996 57394 21048 57400
rect 1872 57050 1900 57394
rect 3068 57050 3096 57394
rect 3424 57248 3476 57254
rect 3424 57190 3476 57196
rect 1860 57044 1912 57050
rect 1860 56986 1912 56992
rect 3056 57044 3108 57050
rect 3056 56986 3108 56992
rect 3436 55758 3464 57190
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4632 57050 4660 57394
rect 5724 57384 5776 57390
rect 5724 57326 5776 57332
rect 4620 57044 4672 57050
rect 4620 56986 4672 56992
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 1768 55752 1820 55758
rect 1674 55720 1730 55729
rect 1768 55694 1820 55700
rect 3424 55752 3476 55758
rect 3424 55694 3476 55700
rect 1674 55655 1730 55664
rect 1688 55622 1716 55655
rect 1676 55616 1728 55622
rect 1676 55558 1728 55564
rect 1676 55072 1728 55078
rect 1676 55014 1728 55020
rect 1688 54913 1716 55014
rect 1674 54904 1730 54913
rect 1674 54839 1730 54848
rect 1674 54088 1730 54097
rect 1674 54023 1676 54032
rect 1728 54023 1730 54032
rect 1676 53994 1728 54000
rect 1676 53440 1728 53446
rect 1676 53382 1728 53388
rect 1688 53281 1716 53382
rect 1674 53272 1730 53281
rect 1674 53207 1730 53216
rect 1676 52624 1728 52630
rect 1676 52566 1728 52572
rect 1688 52465 1716 52566
rect 1674 52456 1730 52465
rect 1674 52391 1730 52400
rect 1676 51808 1728 51814
rect 1676 51750 1728 51756
rect 1688 51649 1716 51750
rect 1674 51640 1730 51649
rect 1674 51575 1730 51584
rect 1674 50824 1730 50833
rect 1674 50759 1676 50768
rect 1728 50759 1730 50768
rect 1676 50730 1728 50736
rect 1676 50176 1728 50182
rect 1676 50118 1728 50124
rect 1688 50017 1716 50118
rect 1674 50008 1730 50017
rect 1674 49943 1730 49952
rect 1674 49192 1730 49201
rect 1674 49127 1730 49136
rect 1688 49094 1716 49127
rect 1676 49088 1728 49094
rect 1676 49030 1728 49036
rect 1676 48544 1728 48550
rect 1676 48486 1728 48492
rect 1688 48385 1716 48486
rect 1674 48376 1730 48385
rect 1674 48311 1730 48320
rect 1674 47560 1730 47569
rect 1674 47495 1676 47504
rect 1728 47495 1730 47504
rect 1676 47466 1728 47472
rect 1676 46912 1728 46918
rect 1676 46854 1728 46860
rect 1688 46753 1716 46854
rect 1674 46744 1730 46753
rect 1674 46679 1730 46688
rect 1674 45928 1730 45937
rect 1674 45863 1730 45872
rect 1688 45830 1716 45863
rect 1676 45824 1728 45830
rect 1676 45766 1728 45772
rect 1676 45280 1728 45286
rect 1676 45222 1728 45228
rect 1688 45121 1716 45222
rect 1674 45112 1730 45121
rect 1674 45047 1730 45056
rect 1674 44296 1730 44305
rect 1674 44231 1676 44240
rect 1728 44231 1730 44240
rect 1676 44202 1728 44208
rect 1676 43648 1728 43654
rect 1676 43590 1728 43596
rect 1688 43489 1716 43590
rect 1674 43480 1730 43489
rect 1674 43415 1730 43424
rect 1674 42664 1730 42673
rect 1674 42599 1730 42608
rect 1688 42566 1716 42599
rect 1676 42560 1728 42566
rect 1676 42502 1728 42508
rect 1676 42016 1728 42022
rect 1676 41958 1728 41964
rect 1688 41857 1716 41958
rect 1674 41848 1730 41857
rect 1674 41783 1730 41792
rect 1674 41032 1730 41041
rect 1674 40967 1676 40976
rect 1728 40967 1730 40976
rect 1676 40938 1728 40944
rect 1676 40384 1728 40390
rect 1676 40326 1728 40332
rect 1688 40225 1716 40326
rect 1674 40216 1730 40225
rect 1674 40151 1730 40160
rect 1674 39400 1730 39409
rect 1674 39335 1730 39344
rect 1688 39302 1716 39335
rect 1676 39296 1728 39302
rect 1676 39238 1728 39244
rect 1676 38752 1728 38758
rect 1676 38694 1728 38700
rect 1688 38593 1716 38694
rect 1674 38584 1730 38593
rect 1674 38519 1730 38528
rect 1674 37768 1730 37777
rect 1674 37703 1676 37712
rect 1728 37703 1730 37712
rect 1676 37674 1728 37680
rect 1676 37120 1728 37126
rect 1676 37062 1728 37068
rect 1688 36961 1716 37062
rect 1674 36952 1730 36961
rect 1674 36887 1730 36896
rect 1674 36136 1730 36145
rect 1674 36071 1730 36080
rect 1688 36038 1716 36071
rect 1676 36032 1728 36038
rect 1676 35974 1728 35980
rect 1676 35488 1728 35494
rect 1676 35430 1728 35436
rect 1688 35329 1716 35430
rect 1674 35320 1730 35329
rect 1674 35255 1730 35264
rect 1674 34504 1730 34513
rect 1674 34439 1676 34448
rect 1728 34439 1730 34448
rect 1676 34410 1728 34416
rect 1676 33856 1728 33862
rect 1676 33798 1728 33804
rect 1688 33697 1716 33798
rect 1674 33688 1730 33697
rect 1674 33623 1730 33632
rect 1674 32872 1730 32881
rect 1674 32807 1730 32816
rect 1688 32774 1716 32807
rect 1676 32768 1728 32774
rect 1676 32710 1728 32716
rect 1676 32224 1728 32230
rect 1676 32166 1728 32172
rect 1688 32065 1716 32166
rect 1674 32056 1730 32065
rect 1674 31991 1730 32000
rect 1674 31240 1730 31249
rect 1674 31175 1676 31184
rect 1728 31175 1730 31184
rect 1676 31146 1728 31152
rect 1676 30592 1728 30598
rect 1676 30534 1728 30540
rect 1688 30433 1716 30534
rect 1674 30424 1730 30433
rect 1674 30359 1730 30368
rect 1674 29608 1730 29617
rect 1674 29543 1730 29552
rect 1688 29510 1716 29543
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1676 29028 1728 29034
rect 1676 28970 1728 28976
rect 1688 28801 1716 28970
rect 1674 28792 1730 28801
rect 1674 28727 1730 28736
rect 1674 27976 1730 27985
rect 1674 27911 1676 27920
rect 1728 27911 1730 27920
rect 1676 27882 1728 27888
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1688 27169 1716 27270
rect 1674 27160 1730 27169
rect 1674 27095 1730 27104
rect 1676 26512 1728 26518
rect 1676 26454 1728 26460
rect 1688 26353 1716 26454
rect 1674 26344 1730 26353
rect 1674 26279 1730 26288
rect 1780 26234 1808 55694
rect 3516 55276 3568 55282
rect 3516 55218 3568 55224
rect 2412 50176 2464 50182
rect 2412 50118 2464 50124
rect 2424 49978 2452 50118
rect 2412 49972 2464 49978
rect 2412 49914 2464 49920
rect 2412 49088 2464 49094
rect 2412 49030 2464 49036
rect 2424 48890 2452 49030
rect 2412 48884 2464 48890
rect 2412 48826 2464 48832
rect 2412 48748 2464 48754
rect 2412 48690 2464 48696
rect 2424 48550 2452 48690
rect 2412 48544 2464 48550
rect 2412 48486 2464 48492
rect 1860 45960 1912 45966
rect 1860 45902 1912 45908
rect 1504 26206 1808 26234
rect 1504 11014 1532 26206
rect 1872 25974 1900 45902
rect 1952 44396 2004 44402
rect 1952 44338 2004 44344
rect 1964 27334 1992 44338
rect 2228 32904 2280 32910
rect 2228 32846 2280 32852
rect 1952 27328 2004 27334
rect 1952 27270 2004 27276
rect 2136 26444 2188 26450
rect 2136 26386 2188 26392
rect 2044 26308 2096 26314
rect 2044 26250 2096 26256
rect 1860 25968 1912 25974
rect 1860 25910 1912 25916
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 1674 25528 1730 25537
rect 1674 25463 1676 25472
rect 1728 25463 1730 25472
rect 1676 25434 1728 25440
rect 1780 25158 1808 25842
rect 1768 25152 1820 25158
rect 1768 25094 1820 25100
rect 1674 24712 1730 24721
rect 1674 24647 1676 24656
rect 1728 24647 1730 24656
rect 1676 24618 1728 24624
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1688 23905 1716 24006
rect 1674 23896 1730 23905
rect 1674 23831 1730 23840
rect 1674 23080 1730 23089
rect 1674 23015 1730 23024
rect 1688 22982 1716 23015
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1674 22264 1730 22273
rect 1674 22199 1676 22208
rect 1728 22199 1730 22208
rect 1676 22170 1728 22176
rect 1674 21448 1730 21457
rect 1674 21383 1676 21392
rect 1728 21383 1730 21392
rect 1676 21354 1728 21360
rect 1674 20632 1730 20641
rect 1674 20567 1676 20576
rect 1728 20567 1730 20576
rect 1676 20538 1728 20544
rect 1674 19816 1730 19825
rect 1674 19751 1730 19760
rect 1688 19718 1716 19751
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1688 19009 1716 19110
rect 1674 19000 1730 19009
rect 1674 18935 1730 18944
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 18193 1716 18566
rect 1674 18184 1730 18193
rect 1674 18119 1730 18128
rect 1780 17610 1808 25094
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1872 20874 1900 21966
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 2056 19938 2084 26250
rect 2148 25838 2176 26386
rect 2136 25832 2188 25838
rect 2136 25774 2188 25780
rect 2148 24750 2176 25774
rect 2240 25378 2268 32846
rect 2320 30728 2372 30734
rect 2320 30670 2372 30676
rect 2332 25838 2360 30670
rect 2424 28218 2452 48486
rect 3528 45626 3556 55218
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4804 53984 4856 53990
rect 4804 53926 4856 53932
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 3516 45620 3568 45626
rect 3516 45562 3568 45568
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 2504 42016 2556 42022
rect 2504 41958 2556 41964
rect 2516 41818 2544 41958
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 2504 41812 2556 41818
rect 2504 41754 2556 41760
rect 3516 40928 3568 40934
rect 3516 40870 3568 40876
rect 3424 39296 3476 39302
rect 3424 39238 3476 39244
rect 2596 37664 2648 37670
rect 2596 37606 2648 37612
rect 2608 37466 2636 37606
rect 2596 37460 2648 37466
rect 2596 37402 2648 37408
rect 2504 37120 2556 37126
rect 2504 37062 2556 37068
rect 2412 28212 2464 28218
rect 2412 28154 2464 28160
rect 2516 26926 2544 37062
rect 2688 33992 2740 33998
rect 2688 33934 2740 33940
rect 2596 26988 2648 26994
rect 2596 26930 2648 26936
rect 2504 26920 2556 26926
rect 2504 26862 2556 26868
rect 2608 26314 2636 26930
rect 2596 26308 2648 26314
rect 2596 26250 2648 26256
rect 2700 25922 2728 33934
rect 3436 32502 3464 39238
rect 3528 35222 3556 40870
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 3700 40384 3752 40390
rect 3700 40326 3752 40332
rect 3712 40186 3740 40326
rect 3700 40180 3752 40186
rect 3700 40122 3752 40128
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3516 35216 3568 35222
rect 3516 35158 3568 35164
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3424 32496 3476 32502
rect 3424 32438 3476 32444
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4068 31340 4120 31346
rect 4068 31282 4120 31288
rect 3056 29300 3108 29306
rect 3056 29242 3108 29248
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 2884 26382 2912 26726
rect 2872 26376 2924 26382
rect 2872 26318 2924 26324
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2516 25894 2728 25922
rect 2320 25832 2372 25838
rect 2320 25774 2372 25780
rect 2412 25696 2464 25702
rect 2412 25638 2464 25644
rect 2240 25350 2360 25378
rect 2228 25288 2280 25294
rect 2228 25230 2280 25236
rect 2136 24744 2188 24750
rect 2136 24686 2188 24692
rect 2148 23662 2176 24686
rect 2240 24614 2268 25230
rect 2228 24608 2280 24614
rect 2228 24550 2280 24556
rect 2136 23656 2188 23662
rect 2136 23598 2188 23604
rect 2148 22574 2176 23598
rect 2240 22930 2268 24550
rect 2332 23746 2360 25350
rect 2424 25294 2452 25638
rect 2412 25288 2464 25294
rect 2412 25230 2464 25236
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2424 24070 2452 24754
rect 2412 24064 2464 24070
rect 2412 24006 2464 24012
rect 2424 23866 2452 24006
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 2332 23718 2452 23746
rect 2424 23662 2452 23718
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2320 23520 2372 23526
rect 2320 23462 2372 23468
rect 2332 23118 2360 23462
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2240 22902 2360 22930
rect 2136 22568 2188 22574
rect 2136 22510 2188 22516
rect 2148 22098 2176 22510
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 1964 19910 2084 19938
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 1768 17604 1820 17610
rect 1768 17546 1820 17552
rect 1674 17368 1730 17377
rect 1674 17303 1676 17312
rect 1728 17303 1730 17312
rect 1676 17274 1728 17280
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1674 16552 1730 16561
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1596 3466 1624 16526
rect 1674 16487 1730 16496
rect 1688 16454 1716 16487
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1674 14920 1730 14929
rect 1674 14855 1676 14864
rect 1728 14855 1730 14864
rect 1676 14826 1728 14832
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1674 14104 1730 14113
rect 1674 14039 1676 14048
rect 1728 14039 1730 14048
rect 1676 14010 1728 14016
rect 1674 13288 1730 13297
rect 1674 13223 1730 13232
rect 1688 13190 1716 13223
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12481 1716 12582
rect 1674 12472 1730 12481
rect 1674 12407 1730 12416
rect 1674 11656 1730 11665
rect 1674 11591 1730 11600
rect 1688 11354 1716 11591
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1674 10840 1730 10849
rect 1674 10775 1676 10784
rect 1728 10775 1730 10784
rect 1676 10746 1728 10752
rect 1674 10024 1730 10033
rect 1674 9959 1730 9968
rect 1688 9926 1716 9959
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1674 9208 1730 9217
rect 1674 9143 1730 9152
rect 1688 8634 1716 9143
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1674 8392 1730 8401
rect 1674 8327 1730 8336
rect 1688 8090 1716 8327
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1674 6760 1730 6769
rect 1674 6695 1730 6704
rect 1688 6458 1716 6695
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1674 5944 1730 5953
rect 1674 5879 1676 5888
rect 1728 5879 1730 5888
rect 1676 5850 1728 5856
rect 1674 5128 1730 5137
rect 1674 5063 1676 5072
rect 1728 5063 1730 5072
rect 1676 5034 1728 5040
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1688 4321 1716 4422
rect 1674 4312 1730 4321
rect 1674 4247 1730 4256
rect 1584 3460 1636 3466
rect 1584 3402 1636 3408
rect 1780 3194 1808 14282
rect 1872 12238 1900 18702
rect 1964 18426 1992 19910
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1964 3398 1992 18362
rect 2056 15706 2084 19790
rect 2148 17746 2176 20402
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 2240 18222 2268 19314
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2136 17604 2188 17610
rect 2136 17546 2188 17552
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2148 14346 2176 17546
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2240 14278 2268 17138
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 13462 2268 14214
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 12782 2084 13262
rect 2332 13258 2360 22902
rect 2516 22778 2544 25894
rect 2688 25832 2740 25838
rect 2688 25774 2740 25780
rect 2596 24744 2648 24750
rect 2596 24686 2648 24692
rect 2608 24410 2636 24686
rect 2596 24404 2648 24410
rect 2596 24346 2648 24352
rect 2700 23662 2728 25774
rect 2596 23656 2648 23662
rect 2596 23598 2648 23604
rect 2688 23656 2740 23662
rect 2688 23598 2740 23604
rect 2608 23254 2636 23598
rect 2596 23248 2648 23254
rect 2596 23190 2648 23196
rect 2688 23112 2740 23118
rect 2688 23054 2740 23060
rect 2700 22778 2728 23054
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2516 21894 2544 22714
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2596 21548 2648 21554
rect 2596 21490 2648 21496
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2516 18222 2544 18566
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2424 16454 2452 17682
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2516 16658 2544 16934
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2424 13190 2452 13806
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2424 12714 2452 13126
rect 2412 12708 2464 12714
rect 2412 12650 2464 12656
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2332 12238 2360 12582
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2332 6914 2360 12174
rect 2608 11898 2636 21490
rect 2792 21350 2820 25978
rect 2884 21690 2912 26318
rect 3068 22094 3096 29242
rect 3608 28756 3660 28762
rect 3608 28698 3660 28704
rect 3332 25832 3384 25838
rect 3332 25774 3384 25780
rect 3148 25492 3200 25498
rect 3148 25434 3200 25440
rect 3160 25158 3188 25434
rect 3240 25356 3292 25362
rect 3240 25298 3292 25304
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 3148 22976 3200 22982
rect 3148 22918 3200 22924
rect 3160 22234 3188 22918
rect 3252 22778 3280 25298
rect 3344 23798 3372 25774
rect 3516 24608 3568 24614
rect 3516 24550 3568 24556
rect 3528 24206 3556 24550
rect 3516 24200 3568 24206
rect 3516 24142 3568 24148
rect 3332 23792 3384 23798
rect 3332 23734 3384 23740
rect 3344 22930 3372 23734
rect 3344 22902 3464 22930
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3436 22658 3464 22902
rect 3252 22630 3464 22658
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 3068 22066 3188 22094
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2976 21010 3004 21286
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2700 20466 2728 20742
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2700 18426 2728 18702
rect 2976 18630 3004 20946
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 3068 20806 3096 20878
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2976 18290 3004 18566
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2976 17814 3004 18226
rect 2964 17808 3016 17814
rect 2964 17750 3016 17756
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 17202 2728 17478
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2976 16998 3004 17750
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2976 15910 3004 16934
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 15502 3004 15846
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 15026 2728 15302
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2976 14482 3004 15438
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 13938 2728 14214
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2976 13870 3004 14418
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 12306 3004 13806
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 3068 12646 3096 12854
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2608 11558 2636 11834
rect 2976 11694 3004 12242
rect 3160 11830 3188 22066
rect 3252 15706 3280 22630
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3344 17678 3372 22510
rect 3620 22094 3648 28698
rect 3976 27056 4028 27062
rect 3976 26998 4028 27004
rect 3988 26450 4016 26998
rect 4080 26586 4108 31282
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 3976 26444 4028 26450
rect 3976 26386 4028 26392
rect 3700 26240 3752 26246
rect 3700 26182 3752 26188
rect 3712 25906 3740 26182
rect 3988 25906 4016 26386
rect 4632 26382 4660 32370
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3976 25900 4028 25906
rect 3976 25842 4028 25848
rect 3884 25696 3936 25702
rect 3884 25638 3936 25644
rect 3436 22066 3648 22094
rect 3436 20806 3464 22066
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3344 15910 3372 16050
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3252 15434 3280 15642
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2976 11354 3004 11630
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 3160 11150 3188 11766
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 10266 2452 10542
rect 2608 10470 2636 11086
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2424 9178 2452 9454
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2424 8498 2452 9114
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2516 7954 2544 8774
rect 2608 8634 2636 10406
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9654 2820 9862
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2792 9042 2820 9590
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 3160 8974 3188 11086
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2976 8498 3004 8774
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7585 2452 7686
rect 2410 7576 2466 7585
rect 2410 7511 2466 7520
rect 2792 7342 2820 7822
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 3160 7274 3188 8026
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 2332 6886 2636 6914
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2332 6322 2360 6598
rect 2516 6322 2544 6598
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2332 5846 2360 6258
rect 2320 5840 2372 5846
rect 2608 5794 2636 6886
rect 2884 6866 2912 7210
rect 3252 6866 3280 15370
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 2884 6458 2912 6802
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2700 5914 2728 6054
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2320 5782 2372 5788
rect 2424 5766 2636 5794
rect 2424 4282 2452 5766
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 2240 1834 2268 3334
rect 2424 2446 2452 3878
rect 2516 3670 2544 4558
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 2516 3194 2544 3606
rect 2608 3534 2636 5646
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2700 4078 2728 5170
rect 2884 4826 2912 6394
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2608 3194 2636 3470
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 2514 2636 2994
rect 2700 2990 2728 4014
rect 2884 4010 2912 4762
rect 3344 4214 3372 15846
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3620 12986 3648 13466
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3804 9654 3832 20742
rect 3896 20398 3924 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 4080 22982 4108 23258
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22094 4660 26318
rect 4632 22066 4752 22094
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 3884 20392 3936 20398
rect 4172 20346 4200 20810
rect 4724 20602 4752 22066
rect 4816 20806 4844 53926
rect 5736 53446 5764 57326
rect 6012 57050 6040 57394
rect 6656 57050 6684 57394
rect 8300 57384 8352 57390
rect 8300 57326 8352 57332
rect 6920 57248 6972 57254
rect 6920 57190 6972 57196
rect 6000 57044 6052 57050
rect 6000 56986 6052 56992
rect 6644 57044 6696 57050
rect 6644 56986 6696 56992
rect 6932 55962 6960 57190
rect 6920 55956 6972 55962
rect 6920 55898 6972 55904
rect 8312 55350 8340 57326
rect 8496 57050 8524 57394
rect 9048 57050 9076 57394
rect 9312 57248 9364 57254
rect 9312 57190 9364 57196
rect 11888 57248 11940 57254
rect 11888 57190 11940 57196
rect 8484 57044 8536 57050
rect 8484 56986 8536 56992
rect 9036 57044 9088 57050
rect 9036 56986 9088 56992
rect 9324 56982 9352 57190
rect 9312 56976 9364 56982
rect 9312 56918 9364 56924
rect 11900 56914 11928 57190
rect 12636 57050 12664 57394
rect 12900 57248 12952 57254
rect 12900 57190 12952 57196
rect 12624 57044 12676 57050
rect 12624 56986 12676 56992
rect 11888 56908 11940 56914
rect 11888 56850 11940 56856
rect 12912 56846 12940 57190
rect 15028 57050 15056 57394
rect 16304 57248 16356 57254
rect 16304 57190 16356 57196
rect 17040 57248 17092 57254
rect 17040 57190 17092 57196
rect 16316 57050 16344 57190
rect 15016 57044 15068 57050
rect 15016 56986 15068 56992
rect 16304 57044 16356 57050
rect 16304 56986 16356 56992
rect 12900 56840 12952 56846
rect 12900 56782 12952 56788
rect 17052 56710 17080 57190
rect 17420 56778 17448 57394
rect 18972 57384 19024 57390
rect 18972 57326 19024 57332
rect 18880 57248 18932 57254
rect 18880 57190 18932 57196
rect 17868 56976 17920 56982
rect 17868 56918 17920 56924
rect 17408 56772 17460 56778
rect 17408 56714 17460 56720
rect 17040 56704 17092 56710
rect 17040 56646 17092 56652
rect 17880 56438 17908 56918
rect 17868 56432 17920 56438
rect 17868 56374 17920 56380
rect 8300 55344 8352 55350
rect 8300 55286 8352 55292
rect 18892 54126 18920 57190
rect 18984 55622 19012 57326
rect 19996 57050 20024 57394
rect 20812 57316 20864 57322
rect 20812 57258 20864 57264
rect 19984 57044 20036 57050
rect 19984 56986 20036 56992
rect 20444 56908 20496 56914
rect 20444 56850 20496 56856
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 18972 55616 19024 55622
rect 18972 55558 19024 55564
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 20456 54602 20484 56850
rect 20824 56846 20852 57258
rect 21652 57050 21680 57734
rect 22008 57588 22060 57594
rect 22008 57530 22060 57536
rect 21916 57520 21968 57526
rect 21916 57462 21968 57468
rect 21640 57044 21692 57050
rect 21640 56986 21692 56992
rect 20720 56840 20772 56846
rect 20720 56782 20772 56788
rect 20812 56840 20864 56846
rect 20812 56782 20864 56788
rect 20444 54596 20496 54602
rect 20444 54538 20496 54544
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 20732 54262 20760 56782
rect 21364 56772 21416 56778
rect 21364 56714 21416 56720
rect 21376 56370 21404 56714
rect 21364 56364 21416 56370
rect 21364 56306 21416 56312
rect 21824 56364 21876 56370
rect 21824 56306 21876 56312
rect 21364 55684 21416 55690
rect 21364 55626 21416 55632
rect 21376 55282 21404 55626
rect 21836 55282 21864 56306
rect 21364 55276 21416 55282
rect 21364 55218 21416 55224
rect 21824 55276 21876 55282
rect 21824 55218 21876 55224
rect 21376 54670 21404 55218
rect 21364 54664 21416 54670
rect 21364 54606 21416 54612
rect 20720 54256 20772 54262
rect 20720 54198 20772 54204
rect 21376 54194 21404 54606
rect 21928 54330 21956 57462
rect 22020 56506 22048 57530
rect 22204 57458 22232 59200
rect 23400 57458 23428 59200
rect 24596 57458 24624 59200
rect 25792 57594 25820 59200
rect 26240 57860 26292 57866
rect 26240 57802 26292 57808
rect 25780 57588 25832 57594
rect 25780 57530 25832 57536
rect 22192 57452 22244 57458
rect 22192 57394 22244 57400
rect 23388 57452 23440 57458
rect 23388 57394 23440 57400
rect 24584 57452 24636 57458
rect 24584 57394 24636 57400
rect 22204 57050 22232 57394
rect 22284 57248 22336 57254
rect 22284 57190 22336 57196
rect 22468 57248 22520 57254
rect 22468 57190 22520 57196
rect 22192 57044 22244 57050
rect 22192 56986 22244 56992
rect 22100 56976 22152 56982
rect 22100 56918 22152 56924
rect 22008 56500 22060 56506
rect 22008 56442 22060 56448
rect 22112 56370 22140 56918
rect 22296 56914 22324 57190
rect 22480 56982 22508 57190
rect 24596 57050 24624 57394
rect 25044 57316 25096 57322
rect 25044 57258 25096 57264
rect 24860 57248 24912 57254
rect 24860 57190 24912 57196
rect 24584 57044 24636 57050
rect 24584 56986 24636 56992
rect 22468 56976 22520 56982
rect 22468 56918 22520 56924
rect 22284 56908 22336 56914
rect 22284 56850 22336 56856
rect 24768 56432 24820 56438
rect 24768 56374 24820 56380
rect 22100 56364 22152 56370
rect 22100 56306 22152 56312
rect 23480 56364 23532 56370
rect 23480 56306 23532 56312
rect 23848 56364 23900 56370
rect 23848 56306 23900 56312
rect 23112 56160 23164 56166
rect 23112 56102 23164 56108
rect 23296 56160 23348 56166
rect 23296 56102 23348 56108
rect 23124 55758 23152 56102
rect 23308 55758 23336 56102
rect 23492 55865 23520 56306
rect 23860 55962 23888 56306
rect 23848 55956 23900 55962
rect 23848 55898 23900 55904
rect 23756 55888 23808 55894
rect 23478 55856 23534 55865
rect 23756 55830 23808 55836
rect 23478 55791 23534 55800
rect 23112 55752 23164 55758
rect 23112 55694 23164 55700
rect 23296 55752 23348 55758
rect 23296 55694 23348 55700
rect 23572 54528 23624 54534
rect 23572 54470 23624 54476
rect 21916 54324 21968 54330
rect 21916 54266 21968 54272
rect 23584 54194 23612 54470
rect 21364 54188 21416 54194
rect 21364 54130 21416 54136
rect 23572 54188 23624 54194
rect 23572 54130 23624 54136
rect 18880 54120 18932 54126
rect 18880 54062 18932 54068
rect 23388 53984 23440 53990
rect 23388 53926 23440 53932
rect 23400 53582 23428 53926
rect 11704 53576 11756 53582
rect 11704 53518 11756 53524
rect 23388 53576 23440 53582
rect 23388 53518 23440 53524
rect 5724 53440 5776 53446
rect 5724 53382 5776 53388
rect 5540 52488 5592 52494
rect 5540 52430 5592 52436
rect 4896 51808 4948 51814
rect 4896 51750 4948 51756
rect 4908 44878 4936 51750
rect 5552 47598 5580 52430
rect 5540 47592 5592 47598
rect 5540 47534 5592 47540
rect 9220 47456 9272 47462
rect 9220 47398 9272 47404
rect 6644 46980 6696 46986
rect 6644 46922 6696 46928
rect 4896 44872 4948 44878
rect 4896 44814 4948 44820
rect 5264 43648 5316 43654
rect 5264 43590 5316 43596
rect 4896 27872 4948 27878
rect 4896 27814 4948 27820
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 3884 20334 3936 20340
rect 4080 20318 4200 20346
rect 4712 20324 4764 20330
rect 4080 19938 4108 20318
rect 4712 20266 4764 20272
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4080 19910 4200 19938
rect 4172 19514 4200 19910
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4724 19310 4752 20266
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3896 13394 3924 14010
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3436 9042 3464 9454
rect 3804 9382 3832 9590
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3528 9042 3556 9318
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3436 8566 3464 8978
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3436 8090 3464 8502
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 7002 3556 7142
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3712 6798 3740 8774
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3332 4208 3384 4214
rect 3332 4150 3384 4156
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 2884 3602 2912 3946
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2884 2922 2912 3538
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3058 3004 3334
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2884 2774 2912 2858
rect 2792 2746 2912 2774
rect 2792 2582 2820 2746
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2424 2122 2452 2382
rect 2332 2094 2452 2122
rect 2228 1828 2280 1834
rect 2228 1770 2280 1776
rect 2332 800 2360 2094
rect 3436 800 3464 3946
rect 3528 1970 3556 6666
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3620 3058 3648 3878
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3804 2038 3832 9318
rect 3988 7546 4016 17478
rect 4908 17270 4936 27814
rect 5276 27402 5304 43590
rect 6276 42560 6328 42566
rect 6276 42502 6328 42508
rect 5356 27872 5408 27878
rect 5356 27814 5408 27820
rect 5368 27470 5396 27814
rect 5724 27668 5776 27674
rect 5724 27610 5776 27616
rect 5356 27464 5408 27470
rect 5356 27406 5408 27412
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5264 27396 5316 27402
rect 5264 27338 5316 27344
rect 5368 25498 5396 27406
rect 5460 26858 5488 27406
rect 5736 26994 5764 27610
rect 6184 27532 6236 27538
rect 6184 27474 6236 27480
rect 5908 27396 5960 27402
rect 5908 27338 5960 27344
rect 5724 26988 5776 26994
rect 5724 26930 5776 26936
rect 5448 26852 5500 26858
rect 5448 26794 5500 26800
rect 5460 26314 5488 26794
rect 5920 26790 5948 27338
rect 6196 27130 6224 27474
rect 6184 27124 6236 27130
rect 6184 27066 6236 27072
rect 5632 26784 5684 26790
rect 5632 26726 5684 26732
rect 5908 26784 5960 26790
rect 5908 26726 5960 26732
rect 5644 26314 5672 26726
rect 5448 26308 5500 26314
rect 5448 26250 5500 26256
rect 5632 26308 5684 26314
rect 5632 26250 5684 26256
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 5080 23792 5132 23798
rect 5080 23734 5132 23740
rect 5092 22710 5120 23734
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 5368 22710 5396 22986
rect 5080 22704 5132 22710
rect 5080 22646 5132 22652
rect 5356 22704 5408 22710
rect 5356 22646 5408 22652
rect 5092 21978 5120 22646
rect 5092 21962 5304 21978
rect 5092 21956 5316 21962
rect 5092 21950 5264 21956
rect 5264 21898 5316 21904
rect 5276 20534 5304 21898
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5276 19718 5304 20470
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5276 19446 5304 19654
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4264 15162 4292 15506
rect 5368 15434 5396 16458
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5368 15162 5396 15370
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3988 7274 4016 7482
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 3988 7154 4016 7210
rect 3896 7126 4016 7154
rect 3896 2310 3924 7126
rect 4080 6934 4108 7278
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3988 3942 4016 4762
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 3194 4016 3470
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4080 2582 4108 6734
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4816 5370 4844 12718
rect 5184 12434 5212 13194
rect 5460 12918 5488 26250
rect 5540 25424 5592 25430
rect 5540 25366 5592 25372
rect 5552 23798 5580 25366
rect 5540 23792 5592 23798
rect 5540 23734 5592 23740
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5736 15094 5764 19722
rect 5920 18426 5948 26726
rect 6196 26450 6224 27066
rect 6184 26444 6236 26450
rect 6184 26386 6236 26392
rect 6000 21956 6052 21962
rect 6000 21898 6052 21904
rect 6012 20398 6040 21898
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 6012 19378 6040 20334
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6196 16590 6224 18158
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 15570 6224 16526
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 6288 13870 6316 42502
rect 6368 29028 6420 29034
rect 6368 28970 6420 28976
rect 6380 24138 6408 28970
rect 6552 28960 6604 28966
rect 6552 28902 6604 28908
rect 6564 28558 6592 28902
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6460 28416 6512 28422
rect 6460 28358 6512 28364
rect 6368 24132 6420 24138
rect 6368 24074 6420 24080
rect 6472 15094 6500 28358
rect 6656 26450 6684 46922
rect 7472 45620 7524 45626
rect 7472 45562 7524 45568
rect 7012 35692 7064 35698
rect 7012 35634 7064 35640
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 6932 28762 6960 29106
rect 7024 29102 7052 35634
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6644 26444 6696 26450
rect 6644 26386 6696 26392
rect 6552 26376 6604 26382
rect 6552 26318 6604 26324
rect 6564 25770 6592 26318
rect 6552 25764 6604 25770
rect 6552 25706 6604 25712
rect 6656 23730 6684 26386
rect 6736 26240 6788 26246
rect 6736 26182 6788 26188
rect 6748 25498 6776 26182
rect 6736 25492 6788 25498
rect 6736 25434 6788 25440
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6644 23588 6696 23594
rect 6644 23530 6696 23536
rect 6656 23186 6684 23530
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6656 22030 6684 23122
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6840 18222 6868 26726
rect 7196 26240 7248 26246
rect 7196 26182 7248 26188
rect 7208 25906 7236 26182
rect 7196 25900 7248 25906
rect 7196 25842 7248 25848
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6460 15088 6512 15094
rect 6460 15030 6512 15036
rect 6564 14822 6592 15098
rect 6840 15008 6868 15506
rect 6920 15020 6972 15026
rect 6840 14980 6920 15008
rect 6920 14962 6972 14968
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5184 12406 5396 12434
rect 5368 12170 5396 12406
rect 6932 12306 6960 13262
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5368 11830 5396 12106
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5368 9450 5396 11766
rect 6932 11762 6960 12242
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5368 8906 5396 9386
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 7392 8430 7420 8910
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6656 7954 6684 8298
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 7392 7886 7420 8366
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6656 6730 6684 7754
rect 7392 7342 7420 7822
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7392 6798 7420 7278
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6656 5642 6684 6666
rect 7392 5778 7420 6734
rect 7484 6390 7512 45562
rect 7564 36032 7616 36038
rect 7564 35974 7616 35980
rect 7576 26858 7604 35974
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 7840 29096 7892 29102
rect 7840 29038 7892 29044
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7656 27532 7708 27538
rect 7656 27474 7708 27480
rect 7564 26852 7616 26858
rect 7564 26794 7616 26800
rect 7668 18970 7696 27474
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7760 15162 7788 28970
rect 7852 28422 7880 29038
rect 8220 28490 8248 34478
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 8312 28558 8340 29106
rect 9232 29102 9260 47398
rect 9312 45280 9364 45286
rect 9312 45222 9364 45228
rect 9220 29096 9272 29102
rect 9220 29038 9272 29044
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8208 28484 8260 28490
rect 8208 28426 8260 28432
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 7852 27402 7880 28358
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8116 27600 8168 27606
rect 8116 27542 8168 27548
rect 7840 27396 7892 27402
rect 7840 27338 7892 27344
rect 7852 27062 7880 27338
rect 7840 27056 7892 27062
rect 7840 26998 7892 27004
rect 8128 19310 8156 27542
rect 8312 26518 8340 27814
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 8484 26784 8536 26790
rect 8484 26726 8536 26732
rect 8208 26512 8260 26518
rect 8208 26454 8260 26460
rect 8300 26512 8352 26518
rect 8300 26454 8352 26460
rect 8220 22574 8248 26454
rect 8312 25838 8340 26454
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8404 25498 8432 25842
rect 8392 25492 8444 25498
rect 8392 25434 8444 25440
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8312 19446 8340 20334
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 8312 17338 8340 19382
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 8496 12918 8524 26726
rect 8668 26580 8720 26586
rect 8668 26522 8720 26528
rect 8576 22772 8628 22778
rect 8680 22760 8708 26522
rect 8628 22732 8708 22760
rect 8576 22714 8628 22720
rect 8772 19514 8800 27270
rect 9232 27062 9260 27270
rect 9324 27130 9352 45222
rect 11244 35216 11296 35222
rect 11244 35158 11296 35164
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 9968 29306 9996 29446
rect 10704 29306 10732 29446
rect 9956 29300 10008 29306
rect 9956 29242 10008 29248
rect 10692 29300 10744 29306
rect 10692 29242 10744 29248
rect 9968 28762 9996 29242
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 10048 28960 10100 28966
rect 10048 28902 10100 28908
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 9864 28416 9916 28422
rect 9864 28358 9916 28364
rect 9876 28082 9904 28358
rect 10060 28082 10088 28902
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 10048 28076 10100 28082
rect 10048 28018 10100 28024
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9496 27668 9548 27674
rect 9496 27610 9548 27616
rect 9312 27124 9364 27130
rect 9312 27066 9364 27072
rect 9220 27056 9272 27062
rect 9220 26998 9272 27004
rect 9324 26586 9352 27066
rect 9508 26926 9536 27610
rect 9496 26920 9548 26926
rect 9496 26862 9548 26868
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 9508 26518 9536 26862
rect 9496 26512 9548 26518
rect 9496 26454 9548 26460
rect 9128 26308 9180 26314
rect 9128 26250 9180 26256
rect 9140 25974 9168 26250
rect 9128 25968 9180 25974
rect 9128 25910 9180 25916
rect 9312 25764 9364 25770
rect 9312 25706 9364 25712
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 9140 25294 9168 25638
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 9324 23798 9352 25706
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 8944 23792 8996 23798
rect 8944 23734 8996 23740
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 8956 20534 8984 23734
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8956 19530 8984 20470
rect 8760 19508 8812 19514
rect 8956 19502 9076 19530
rect 8760 19450 8812 19456
rect 9048 19446 9076 19502
rect 9036 19440 9088 19446
rect 9036 19382 9088 19388
rect 9048 18358 9076 19382
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9048 16522 9076 18294
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9128 16652 9180 16658
rect 9232 16640 9260 18158
rect 9416 16658 9444 25638
rect 9784 20398 9812 27814
rect 9956 26580 10008 26586
rect 9956 26522 10008 26528
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9180 16612 9260 16640
rect 9404 16652 9456 16658
rect 9128 16594 9180 16600
rect 9404 16594 9456 16600
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9048 15434 9076 16458
rect 9140 16250 9168 16594
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9600 16114 9628 17138
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 9048 15094 9076 15370
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8128 12238 8156 12718
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8312 11694 8340 12174
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8312 10810 8340 11630
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8312 8566 8340 8774
rect 8772 8566 8800 9386
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 3126 4476 3334
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2650 4752 4082
rect 6656 3482 6684 5578
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3738 7328 3878
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 6564 3466 6684 3482
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 6552 3460 6684 3466
rect 6604 3454 6684 3460
rect 6552 3402 6604 3408
rect 5092 3194 5120 3402
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 6656 3126 6684 3454
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 4528 2440 4580 2446
rect 4816 2394 4844 2586
rect 4528 2382 4580 2388
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3792 2032 3844 2038
rect 3792 1974 3844 1980
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 4540 800 4568 2382
rect 4632 2366 4844 2394
rect 5632 2440 5684 2446
rect 6840 2394 6868 3402
rect 6932 3058 6960 3470
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7024 2922 7052 3334
rect 7300 3058 7328 3674
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 6920 2440 6972 2446
rect 5632 2382 5684 2388
rect 6748 2388 6920 2394
rect 6748 2382 6972 2388
rect 4632 2310 4660 2366
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4816 2106 4844 2246
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 5644 800 5672 2382
rect 6748 2366 6960 2382
rect 7852 2378 7880 2790
rect 7944 2514 7972 4014
rect 8956 3738 8984 14894
rect 9048 12918 9076 15030
rect 9968 12986 9996 26522
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10152 22642 10180 23598
rect 10244 23322 10272 28970
rect 10704 28626 10732 29242
rect 10692 28620 10744 28626
rect 10692 28562 10744 28568
rect 10324 28416 10376 28422
rect 10324 28358 10376 28364
rect 10336 28218 10364 28358
rect 10324 28212 10376 28218
rect 10324 28154 10376 28160
rect 10704 27674 10732 28562
rect 10876 28416 10928 28422
rect 10876 28358 10928 28364
rect 10692 27668 10744 27674
rect 10692 27610 10744 27616
rect 10600 27396 10652 27402
rect 10600 27338 10652 27344
rect 10784 27396 10836 27402
rect 10784 27338 10836 27344
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10336 25906 10364 26930
rect 10612 26926 10640 27338
rect 10796 26994 10824 27338
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10612 26586 10640 26862
rect 10600 26580 10652 26586
rect 10600 26522 10652 26528
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10336 25158 10364 25842
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9048 11354 9076 11630
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9042 9536 9998
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9508 8430 9536 8978
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9600 7478 9628 10678
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9692 6390 9720 11766
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9784 9042 9812 9454
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 10152 6866 10180 10542
rect 10336 8906 10364 25094
rect 10428 15706 10456 26386
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10612 22982 10640 25842
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 10704 25498 10732 25774
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10612 16436 10640 22918
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10692 16448 10744 16454
rect 10612 16408 10692 16436
rect 10692 16390 10744 16396
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10796 12102 10824 20742
rect 10888 20602 10916 28358
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11072 18086 11100 18226
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 14822 11100 18022
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11072 14074 11100 14758
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12714 11100 13126
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10796 11830 10824 12038
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9508 5914 9536 6190
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9600 5778 9628 6054
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9600 3534 9628 5714
rect 9692 5642 9720 6326
rect 10152 5846 10180 6802
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9876 3602 9904 4082
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8588 2446 8616 3334
rect 9048 3126 9076 3402
rect 9600 3126 9628 3470
rect 10336 3466 10364 5578
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 7840 2372 7892 2378
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5920 1902 5948 2246
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 6748 800 6776 2366
rect 7840 2314 7892 2320
rect 7852 800 7880 2314
rect 8956 800 8984 2382
rect 10060 2378 10088 2790
rect 10520 2514 10548 8774
rect 11072 3942 11100 9522
rect 11164 4010 11192 12786
rect 11256 9042 11284 35158
rect 11612 27872 11664 27878
rect 11612 27814 11664 27820
rect 11520 27328 11572 27334
rect 11520 27270 11572 27276
rect 11532 26926 11560 27270
rect 11520 26920 11572 26926
rect 11520 26862 11572 26868
rect 11624 23186 11652 27814
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11716 22930 11744 53518
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 16580 50924 16632 50930
rect 16580 50866 16632 50872
rect 13452 49972 13504 49978
rect 13452 49914 13504 49920
rect 13360 48884 13412 48890
rect 13360 48826 13412 48832
rect 11796 40180 11848 40186
rect 11796 40122 11848 40128
rect 11624 22902 11744 22930
rect 11624 20602 11652 22902
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11716 17610 11744 22714
rect 11808 21486 11836 40122
rect 13372 27538 13400 48826
rect 13360 27532 13412 27538
rect 13360 27474 13412 27480
rect 12348 27328 12400 27334
rect 12348 27270 12400 27276
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11900 22778 11928 22986
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11992 21146 12020 26862
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11716 15434 11744 17546
rect 12084 15434 12112 27066
rect 12360 26994 12388 27270
rect 13464 27062 13492 49914
rect 13912 41812 13964 41818
rect 13912 41754 13964 41760
rect 13728 28688 13780 28694
rect 13728 28630 13780 28636
rect 13740 28082 13768 28630
rect 13820 28552 13872 28558
rect 13820 28494 13872 28500
rect 13728 28076 13780 28082
rect 13728 28018 13780 28024
rect 13832 27878 13860 28494
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13832 27062 13860 27814
rect 13452 27056 13504 27062
rect 13280 27004 13452 27010
rect 13280 26998 13504 27004
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 13280 26982 13492 26998
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 12164 26512 12216 26518
rect 12164 26454 12216 26460
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11716 14346 11744 15370
rect 12176 14482 12204 26454
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12452 22642 12480 23054
rect 12728 22710 12756 26726
rect 13004 26382 13032 26726
rect 13280 26586 13308 26982
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 13360 26852 13412 26858
rect 13360 26794 13412 26800
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12716 22704 12768 22710
rect 12716 22646 12768 22652
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12452 21010 12480 22578
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12360 19174 12388 20878
rect 12452 19378 12480 20946
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12360 18714 12388 19110
rect 12636 18834 12664 19314
rect 13188 19310 13216 25638
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12268 18698 12388 18714
rect 12256 18692 12388 18698
rect 12308 18686 12388 18692
rect 12256 18634 12308 18640
rect 12268 18426 12296 18634
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13004 16114 13032 18226
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12544 15502 12572 15846
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 14482 12572 15438
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11716 14006 11744 14282
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11716 13734 11744 13806
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13394 11744 13670
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 11992 11898 12020 12650
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12084 10266 12112 13874
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12176 11898 12204 13194
rect 13004 12646 13032 16050
rect 13280 14618 13308 26522
rect 13372 20874 13400 26794
rect 13464 26382 13492 26862
rect 13832 26518 13860 26998
rect 13820 26512 13872 26518
rect 13820 26454 13872 26460
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13832 21622 13860 22578
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13360 20868 13412 20874
rect 13360 20810 13412 20816
rect 13832 14618 13860 21422
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13832 14074 13860 14554
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13464 12986 13492 13194
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12084 9586 12112 10202
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12176 9450 12204 11834
rect 13004 10742 13032 12582
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13372 11898 13400 12038
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13464 11694 13492 12038
rect 13832 11694 13860 13262
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 13832 10606 13860 11630
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 12176 8906 12204 9386
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9042 13768 9318
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5778 11652 6054
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 12912 5302 12940 8502
rect 13832 8430 13860 8910
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13924 6730 13952 41754
rect 15200 37460 15252 37466
rect 15200 37402 15252 37408
rect 15212 35894 15240 37402
rect 15212 35866 15424 35894
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 14372 28416 14424 28422
rect 14372 28358 14424 28364
rect 14188 27600 14240 27606
rect 14188 27542 14240 27548
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 14016 26926 14044 27474
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14096 26240 14148 26246
rect 14096 26182 14148 26188
rect 14004 25764 14056 25770
rect 14004 25706 14056 25712
rect 14016 17746 14044 25706
rect 14108 21350 14136 26182
rect 14200 22778 14228 27542
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 14292 25158 14320 25774
rect 14280 25152 14332 25158
rect 14280 25094 14332 25100
rect 14292 24614 14320 25094
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 14384 21146 14412 28358
rect 14660 26234 14688 29582
rect 15016 27872 15068 27878
rect 15016 27814 15068 27820
rect 15028 27334 15056 27814
rect 15016 27328 15068 27334
rect 15016 27270 15068 27276
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14752 26586 14780 26930
rect 15028 26926 15056 27270
rect 15108 27056 15160 27062
rect 15108 26998 15160 27004
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15028 26586 15056 26862
rect 14740 26580 14792 26586
rect 14740 26522 14792 26528
rect 15016 26580 15068 26586
rect 15016 26522 15068 26528
rect 15120 26518 15148 26998
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 14660 26206 14780 26234
rect 14464 25832 14516 25838
rect 14464 25774 14516 25780
rect 14476 25498 14504 25774
rect 14464 25492 14516 25498
rect 14464 25434 14516 25440
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14660 19514 14688 24550
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 14752 10248 14780 26206
rect 15396 26042 15424 35866
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15476 26376 15528 26382
rect 15476 26318 15528 26324
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15396 25702 15424 25978
rect 15488 25906 15516 26318
rect 15476 25900 15528 25906
rect 15476 25842 15528 25848
rect 15384 25696 15436 25702
rect 15384 25638 15436 25644
rect 15292 25424 15344 25430
rect 15292 25366 15344 25372
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15212 21622 15240 21898
rect 15200 21616 15252 21622
rect 15200 21558 15252 21564
rect 15212 21010 15240 21558
rect 15304 21486 15332 25366
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 14936 12442 14964 20538
rect 15212 19922 15240 20946
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15212 19394 15240 19858
rect 15120 19366 15240 19394
rect 15120 18834 15148 19366
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15120 18358 15148 18770
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15304 18358 15332 18634
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15396 17882 15424 25638
rect 15488 25158 15516 25842
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 15910 15240 17614
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 15570 15424 15846
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15396 14482 15424 15506
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 14006 15424 14418
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14752 10220 14964 10248
rect 14936 9450 14964 10220
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14844 8974 14872 9386
rect 14936 9178 14964 9386
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 7342 14412 8366
rect 14660 8090 14688 8842
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13924 6390 13952 6666
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 14384 5710 14412 7278
rect 15488 6798 15516 25094
rect 15580 21010 15608 27814
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 15764 26382 15792 26726
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15936 26240 15988 26246
rect 15936 26182 15988 26188
rect 16396 26240 16448 26246
rect 16592 26234 16620 50866
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 17132 47592 17184 47598
rect 17132 47534 17184 47540
rect 16948 32496 17000 32502
rect 16948 32438 17000 32444
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16776 26234 16804 26318
rect 16592 26206 16804 26234
rect 16396 26182 16448 26188
rect 15948 25906 15976 26182
rect 16408 26042 16436 26182
rect 16396 26036 16448 26042
rect 16396 25978 16448 25984
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15672 19922 15700 22374
rect 15948 22234 15976 25638
rect 16776 25158 16804 26206
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 16776 22098 16804 25094
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 16040 20874 16068 21898
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16028 20868 16080 20874
rect 16028 20810 16080 20816
rect 16040 20346 16068 20810
rect 16040 20318 16160 20346
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 16040 17746 16068 20198
rect 16132 19786 16160 20318
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16132 19446 16160 19722
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 16132 18698 16160 19382
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16224 13530 16252 21626
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16304 17264 16356 17270
rect 16304 17206 16356 17212
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 16224 11762 16252 12106
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16316 10470 16344 17206
rect 16684 15434 16712 17546
rect 16960 16590 16988 32438
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 17052 25906 17080 26182
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17144 18834 17172 47534
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 18788 44872 18840 44878
rect 18788 44814 18840 44820
rect 18236 38820 18288 38826
rect 18236 38762 18288 38768
rect 17500 26920 17552 26926
rect 17500 26862 17552 26868
rect 17512 26246 17540 26862
rect 17592 26784 17644 26790
rect 17592 26726 17644 26732
rect 17604 26518 17632 26726
rect 17592 26512 17644 26518
rect 17592 26454 17644 26460
rect 17500 26240 17552 26246
rect 17500 26182 17552 26188
rect 17512 25702 17540 26182
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 17408 25220 17460 25226
rect 17408 25162 17460 25168
rect 17420 22506 17448 25162
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17604 21622 17632 26454
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 18248 21146 18276 38762
rect 18604 24132 18656 24138
rect 18604 24074 18656 24080
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18432 22982 18460 23802
rect 18420 22976 18472 22982
rect 18420 22918 18472 22924
rect 18432 22574 18460 22918
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18236 21140 18288 21146
rect 18236 21082 18288 21088
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17144 18426 17172 18770
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 18248 17882 18276 21082
rect 18432 20058 18460 22510
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 15706 16988 16526
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16684 14346 16712 15370
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16684 14006 16712 14282
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16672 13456 16724 13462
rect 16724 13404 16896 13410
rect 16672 13398 16896 13404
rect 16684 13382 16896 13398
rect 18064 13394 18092 14010
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 10266 16344 10406
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15120 6390 15148 6598
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11992 3738 12020 3878
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 13648 3466 13676 5306
rect 14384 5234 14412 5646
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13648 3126 13676 3402
rect 13740 3194 13768 3606
rect 14292 3534 14320 3674
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 14384 3058 14412 5170
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 11164 2378 11192 2790
rect 12268 2446 12296 2790
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9324 1834 9352 2246
rect 9312 1828 9364 1834
rect 9312 1770 9364 1776
rect 10060 800 10088 2314
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10244 1970 10272 2246
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 11164 800 11192 2314
rect 12268 800 12296 2382
rect 14752 2378 14780 3334
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15580 2378 15608 2790
rect 15948 2582 15976 6734
rect 16592 5846 16620 12718
rect 16684 11830 16712 13194
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16684 10062 16712 11766
rect 16776 10606 16804 12106
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16776 10130 16804 10542
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16868 7426 16896 13382
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 17788 12238 17816 13194
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17972 12306 18000 13126
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18156 10742 18184 11698
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 18156 7478 18184 10678
rect 18616 8022 18644 24074
rect 18800 20602 18828 44814
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 19260 22710 19288 25638
rect 19444 24410 19472 26250
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19260 21894 19288 22646
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 18788 20596 18840 20602
rect 18788 20538 18840 20544
rect 18800 20058 18828 20538
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18800 14482 18828 19994
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18800 12442 18828 14214
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18892 10742 18920 10950
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 19260 8634 19288 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 20180 21350 20208 21490
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 20180 21010 20208 21286
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20466 19380 20742
rect 19444 20482 19472 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19444 20466 19564 20482
rect 19340 20460 19392 20466
rect 19444 20460 19576 20466
rect 19444 20454 19524 20460
rect 19340 20402 19392 20408
rect 19524 20402 19576 20408
rect 19536 19718 19564 20402
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 18766 20024 20198
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19352 16590 19380 17274
rect 19444 16590 19472 17478
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 15570 19472 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19352 13530 19380 14758
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19444 13802 19472 14486
rect 19996 14414 20024 18566
rect 20272 18426 20300 18702
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20180 17610 20208 18226
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 20088 17338 20116 17478
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 20180 15026 20208 17546
rect 20364 16590 20392 22374
rect 20456 20262 20484 24006
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20640 20806 20668 20946
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20456 18086 20484 20198
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20456 17252 20484 18022
rect 20548 17354 20576 19654
rect 20640 17542 20668 20742
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20548 17326 20668 17354
rect 20456 17224 20576 17252
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19996 13326 20024 14214
rect 20088 13938 20116 14758
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19444 12646 19472 12786
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19444 12434 19472 12582
rect 19352 12406 19472 12434
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18616 7546 18644 7958
rect 18800 7750 18828 8570
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 16776 7398 16896 7426
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16592 4826 16620 5782
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16408 3738 16436 4014
rect 16776 4010 16804 7398
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 6254 16896 7278
rect 18156 6662 18184 7414
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16960 5914 16988 6122
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 18156 5574 18184 6598
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18616 5710 18644 6190
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18236 5636 18288 5642
rect 18236 5578 18288 5584
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16776 2922 16804 3946
rect 17604 3466 17632 5510
rect 18248 5370 18276 5578
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17592 3460 17644 3466
rect 17592 3402 17644 3408
rect 17604 3126 17632 3402
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 16684 2378 16712 2858
rect 17788 2446 17816 3878
rect 18616 3534 18644 5646
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 3126 18368 3334
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18616 3058 18644 3470
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18800 2582 18828 7686
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19168 6866 19196 7142
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19352 6202 19380 12406
rect 19812 12238 19840 12582
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19904 11150 19932 11494
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 20088 10674 20116 11698
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10062 19932 10406
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19444 8430 19472 9454
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19536 9042 19564 9318
rect 19628 9178 19656 9318
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 20088 8838 20116 10610
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19996 7886 20024 8774
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 20088 7426 20116 8774
rect 19996 7398 20116 7426
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19444 6322 19472 6598
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19260 6174 19380 6202
rect 19260 4282 19288 6174
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5302 19380 6054
rect 19812 5914 19840 6258
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19444 5114 19472 5646
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19352 5086 19472 5114
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 13372 800 13400 2314
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 2038 13584 2246
rect 13544 2032 13596 2038
rect 13544 1974 13596 1980
rect 14476 800 14504 2314
rect 15580 800 15608 2314
rect 16684 800 16712 2314
rect 17788 800 17816 2382
rect 18892 800 18920 2926
rect 19260 2774 19288 4218
rect 19352 3058 19380 5086
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19444 2922 19472 4082
rect 19536 3942 19564 4082
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19720 3534 19748 3878
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19996 3398 20024 7398
rect 20180 5710 20208 14962
rect 20456 14958 20484 16526
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20364 11694 20392 14418
rect 20456 12782 20484 14894
rect 20548 14482 20576 17224
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20548 13938 20576 14214
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20364 11354 20392 11630
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20456 10606 20484 12718
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20168 5160 20220 5166
rect 20168 5102 20220 5108
rect 20180 4826 20208 5102
rect 20272 5030 20300 5510
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20364 4842 20392 5306
rect 20456 5166 20484 5714
rect 20548 5370 20576 13874
rect 20640 12850 20668 17326
rect 21192 16794 21220 18634
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21468 17882 21496 18294
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21652 16794 21680 17614
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 21192 16658 21220 16730
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 22112 13870 22140 14554
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22204 14074 22232 14350
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22296 13938 22324 16390
rect 23492 14074 23520 17478
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22112 13530 22140 13806
rect 23492 13802 23520 14010
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22572 13530 22600 13670
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22572 12986 22600 13466
rect 23492 12986 23520 13738
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 22480 12442 22508 12922
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22664 12238 22692 12582
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22756 11762 22784 12786
rect 23492 12782 23520 12922
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 20732 10810 20760 11222
rect 21376 11014 21404 11494
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 22112 9450 22140 9930
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20640 6866 20668 8366
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20272 4814 20392 4842
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19168 2746 19288 2774
rect 19168 2514 19196 2746
rect 20088 2514 20116 3946
rect 20180 3534 20208 4422
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20272 2514 20300 4814
rect 20352 4072 20404 4078
rect 20456 4060 20484 5102
rect 20640 4078 20668 6802
rect 21560 6730 21588 7686
rect 21744 7342 21772 8298
rect 21928 8022 21956 8774
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 22112 6798 22140 7686
rect 22204 6866 22232 11154
rect 22572 11150 22600 11494
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22756 9926 22784 11698
rect 23112 11688 23164 11694
rect 23112 11630 23164 11636
rect 23124 11218 23152 11630
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 23388 10600 23440 10606
rect 23388 10542 23440 10548
rect 23400 10130 23428 10542
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22664 9586 22692 9862
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22480 7750 22508 8910
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22572 8498 22600 8774
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 21192 6390 21220 6598
rect 22112 6458 22140 6598
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 21180 6384 21232 6390
rect 21180 6326 21232 6332
rect 22204 6118 22232 6802
rect 22480 6730 22508 7686
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 20404 4032 20484 4060
rect 20628 4072 20680 4078
rect 20352 4014 20404 4020
rect 20628 4014 20680 4020
rect 20364 3602 20392 4014
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20456 2922 20484 3334
rect 20548 3058 20576 3334
rect 21376 3058 21404 4422
rect 22480 4214 22508 6666
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22572 6322 22600 6598
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22664 5914 22692 6054
rect 22652 5908 22704 5914
rect 22652 5850 22704 5856
rect 22468 4208 22520 4214
rect 22468 4150 22520 4156
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22112 3534 22140 3878
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22388 3058 22416 3334
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20088 2122 20116 2450
rect 19996 2094 20116 2122
rect 19996 800 20024 2094
rect 21100 800 21128 2994
rect 22480 2650 22508 4150
rect 22756 3398 22784 9862
rect 23400 9042 23428 10066
rect 23492 9178 23520 12718
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22848 6798 22876 7346
rect 23400 7342 23428 8978
rect 23492 8090 23520 9114
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23124 6798 23152 7142
rect 23492 7002 23520 8026
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 22848 6322 22876 6734
rect 23124 6322 23152 6734
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 22848 5574 22876 6258
rect 23124 6202 23152 6258
rect 23032 6174 23152 6202
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22848 5030 22876 5510
rect 22836 5024 22888 5030
rect 22836 4966 22888 4972
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22756 2650 22784 3334
rect 22848 3058 22876 4966
rect 23032 4486 23060 6174
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 23032 3058 23060 4422
rect 23204 4276 23256 4282
rect 23204 4218 23256 4224
rect 23216 4078 23244 4218
rect 23768 4078 23796 55830
rect 24780 55758 24808 56374
rect 24872 55826 24900 57190
rect 25056 56370 25084 57258
rect 25136 57248 25188 57254
rect 25136 57190 25188 57196
rect 25044 56364 25096 56370
rect 25044 56306 25096 56312
rect 24950 55856 25006 55865
rect 24860 55820 24912 55826
rect 24950 55791 25006 55800
rect 24860 55762 24912 55768
rect 23940 55752 23992 55758
rect 23940 55694 23992 55700
rect 24768 55752 24820 55758
rect 24768 55694 24820 55700
rect 23952 54194 23980 55694
rect 24780 54670 24808 55694
rect 24768 54664 24820 54670
rect 24768 54606 24820 54612
rect 24780 54330 24808 54606
rect 24768 54324 24820 54330
rect 24768 54266 24820 54272
rect 24964 54233 24992 55791
rect 25148 54738 25176 57190
rect 26252 57050 26280 57802
rect 26988 57594 27016 59200
rect 26976 57588 27028 57594
rect 26976 57530 27028 57536
rect 28184 57458 28212 59200
rect 29380 57594 29408 59200
rect 30288 57792 30340 57798
rect 30288 57734 30340 57740
rect 29368 57588 29420 57594
rect 29368 57530 29420 57536
rect 28172 57452 28224 57458
rect 28172 57394 28224 57400
rect 27160 57248 27212 57254
rect 27160 57190 27212 57196
rect 26240 57044 26292 57050
rect 26240 56986 26292 56992
rect 25964 56704 26016 56710
rect 25964 56646 26016 56652
rect 25596 56432 25648 56438
rect 25596 56374 25648 56380
rect 25608 56234 25636 56374
rect 25596 56228 25648 56234
rect 25596 56170 25648 56176
rect 25228 56160 25280 56166
rect 25228 56102 25280 56108
rect 25240 55758 25268 56102
rect 25608 55758 25636 56170
rect 25872 56160 25924 56166
rect 25872 56102 25924 56108
rect 25780 55888 25832 55894
rect 25780 55830 25832 55836
rect 25792 55758 25820 55830
rect 25884 55758 25912 56102
rect 25228 55752 25280 55758
rect 25228 55694 25280 55700
rect 25596 55752 25648 55758
rect 25596 55694 25648 55700
rect 25780 55752 25832 55758
rect 25780 55694 25832 55700
rect 25872 55752 25924 55758
rect 25872 55694 25924 55700
rect 25240 54874 25268 55694
rect 25228 54868 25280 54874
rect 25228 54810 25280 54816
rect 25136 54732 25188 54738
rect 25136 54674 25188 54680
rect 25044 54596 25096 54602
rect 25044 54538 25096 54544
rect 25056 54262 25084 54538
rect 25136 54528 25188 54534
rect 25136 54470 25188 54476
rect 25044 54256 25096 54262
rect 24950 54224 25006 54233
rect 23940 54188 23992 54194
rect 23940 54130 23992 54136
rect 24676 54188 24728 54194
rect 24676 54130 24728 54136
rect 24860 54188 24912 54194
rect 24912 54168 24950 54176
rect 25044 54198 25096 54204
rect 25148 54194 25176 54470
rect 24912 54159 25006 54168
rect 25136 54188 25188 54194
rect 24912 54148 24992 54159
rect 24860 54130 24912 54136
rect 24124 53984 24176 53990
rect 24124 53926 24176 53932
rect 24136 4146 24164 53926
rect 24688 53650 24716 54130
rect 24964 54099 24992 54148
rect 25136 54130 25188 54136
rect 25240 54058 25268 54810
rect 25608 54194 25636 55694
rect 25976 55690 26004 56646
rect 26252 56438 26280 56986
rect 26424 56908 26476 56914
rect 26424 56850 26476 56856
rect 26240 56432 26292 56438
rect 26240 56374 26292 56380
rect 26148 56364 26200 56370
rect 26148 56306 26200 56312
rect 26160 55962 26188 56306
rect 26148 55956 26200 55962
rect 26148 55898 26200 55904
rect 26054 55856 26110 55865
rect 26054 55791 26110 55800
rect 26068 55758 26096 55791
rect 26056 55752 26108 55758
rect 26056 55694 26108 55700
rect 25964 55684 26016 55690
rect 25964 55626 26016 55632
rect 26436 54262 26464 56850
rect 27068 55820 27120 55826
rect 27068 55762 27120 55768
rect 27080 55622 27108 55762
rect 27068 55616 27120 55622
rect 27068 55558 27120 55564
rect 26424 54256 26476 54262
rect 26424 54198 26476 54204
rect 27172 54194 27200 57190
rect 28184 57050 28212 57394
rect 28632 57384 28684 57390
rect 28632 57326 28684 57332
rect 28540 57248 28592 57254
rect 28540 57190 28592 57196
rect 28172 57044 28224 57050
rect 28172 56986 28224 56992
rect 28448 56840 28500 56846
rect 28448 56782 28500 56788
rect 28264 56772 28316 56778
rect 28264 56714 28316 56720
rect 27344 56364 27396 56370
rect 27344 56306 27396 56312
rect 27252 56160 27304 56166
rect 27252 56102 27304 56108
rect 25596 54188 25648 54194
rect 25596 54130 25648 54136
rect 27160 54188 27212 54194
rect 27160 54130 27212 54136
rect 25228 54052 25280 54058
rect 25228 53994 25280 54000
rect 27068 53984 27120 53990
rect 27068 53926 27120 53932
rect 24676 53644 24728 53650
rect 24676 53586 24728 53592
rect 27080 53582 27108 53926
rect 27068 53576 27120 53582
rect 27068 53518 27120 53524
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23216 3602 23244 4014
rect 23204 3596 23256 3602
rect 23204 3538 23256 3544
rect 23204 3460 23256 3466
rect 23204 3402 23256 3408
rect 23216 3194 23244 3402
rect 27264 3194 27292 56102
rect 27356 55826 27384 56306
rect 27344 55820 27396 55826
rect 27344 55762 27396 55768
rect 28276 55758 28304 56714
rect 28356 56364 28408 56370
rect 28356 56306 28408 56312
rect 28368 55962 28396 56306
rect 28460 55962 28488 56782
rect 28356 55956 28408 55962
rect 28356 55898 28408 55904
rect 28448 55956 28500 55962
rect 28448 55898 28500 55904
rect 28264 55752 28316 55758
rect 28264 55694 28316 55700
rect 27344 55276 27396 55282
rect 27344 55218 27396 55224
rect 27356 54233 27384 55218
rect 27896 54732 27948 54738
rect 27896 54674 27948 54680
rect 27908 54262 27936 54674
rect 28276 54330 28304 55694
rect 28264 54324 28316 54330
rect 28264 54266 28316 54272
rect 27896 54256 27948 54262
rect 27342 54224 27398 54233
rect 27896 54198 27948 54204
rect 27342 54159 27344 54168
rect 27396 54159 27398 54168
rect 27344 54130 27396 54136
rect 27344 54052 27396 54058
rect 27344 53994 27396 54000
rect 27356 53786 27384 53994
rect 27344 53780 27396 53786
rect 27344 53722 27396 53728
rect 28276 53242 28304 54266
rect 28460 53786 28488 55898
rect 28552 55826 28580 57190
rect 28644 56370 28672 57326
rect 29736 57248 29788 57254
rect 29736 57190 29788 57196
rect 28908 56976 28960 56982
rect 28908 56918 28960 56924
rect 28920 56506 28948 56918
rect 29748 56914 29776 57190
rect 29736 56908 29788 56914
rect 29736 56850 29788 56856
rect 30104 56704 30156 56710
rect 30104 56646 30156 56652
rect 28724 56500 28776 56506
rect 28724 56442 28776 56448
rect 28908 56500 28960 56506
rect 28908 56442 28960 56448
rect 28632 56364 28684 56370
rect 28632 56306 28684 56312
rect 28736 56234 28764 56442
rect 29828 56432 29880 56438
rect 29826 56400 29828 56409
rect 29880 56400 29882 56409
rect 29000 56364 29052 56370
rect 30116 56370 30144 56646
rect 30194 56536 30250 56545
rect 30194 56471 30250 56480
rect 30208 56438 30236 56471
rect 30196 56432 30248 56438
rect 30196 56374 30248 56380
rect 29826 56335 29882 56344
rect 30104 56364 30156 56370
rect 29000 56306 29052 56312
rect 30300 56352 30328 57734
rect 30576 57458 30604 59200
rect 31772 57458 31800 59200
rect 32968 57458 32996 59200
rect 34164 57594 34192 59200
rect 34152 57588 34204 57594
rect 34152 57530 34204 57536
rect 35360 57458 35388 59200
rect 36556 57458 36584 59200
rect 37752 57458 37780 59200
rect 38948 57458 38976 59200
rect 40144 57458 40172 59200
rect 41340 57458 41368 59200
rect 30564 57452 30616 57458
rect 30564 57394 30616 57400
rect 31760 57452 31812 57458
rect 31760 57394 31812 57400
rect 32128 57452 32180 57458
rect 32128 57394 32180 57400
rect 32956 57452 33008 57458
rect 32956 57394 33008 57400
rect 35348 57452 35400 57458
rect 35348 57394 35400 57400
rect 36544 57452 36596 57458
rect 36544 57394 36596 57400
rect 37740 57452 37792 57458
rect 37740 57394 37792 57400
rect 38936 57452 38988 57458
rect 38936 57394 38988 57400
rect 40132 57452 40184 57458
rect 40132 57394 40184 57400
rect 41328 57452 41380 57458
rect 42536 57440 42564 59200
rect 42892 57520 42944 57526
rect 42892 57462 42944 57468
rect 42800 57452 42852 57458
rect 42536 57412 42800 57440
rect 41328 57394 41380 57400
rect 42800 57394 42852 57400
rect 32140 57050 32168 57394
rect 33140 57316 33192 57322
rect 33140 57258 33192 57264
rect 32496 57248 32548 57254
rect 32496 57190 32548 57196
rect 32128 57044 32180 57050
rect 32128 56986 32180 56992
rect 30932 56500 30984 56506
rect 30932 56442 30984 56448
rect 30564 56364 30616 56370
rect 30300 56324 30564 56352
rect 30104 56306 30156 56312
rect 30944 56352 30972 56442
rect 32508 56438 32536 57190
rect 32496 56432 32548 56438
rect 32496 56374 32548 56380
rect 31116 56364 31168 56370
rect 30944 56324 31116 56352
rect 30564 56306 30616 56312
rect 31116 56306 31168 56312
rect 31300 56364 31352 56370
rect 31300 56306 31352 56312
rect 31484 56364 31536 56370
rect 31484 56306 31536 56312
rect 32956 56364 33008 56370
rect 32956 56306 33008 56312
rect 28724 56228 28776 56234
rect 28724 56170 28776 56176
rect 29012 55962 29040 56306
rect 29092 56296 29144 56302
rect 29092 56238 29144 56244
rect 29000 55956 29052 55962
rect 29000 55898 29052 55904
rect 28540 55820 28592 55826
rect 28540 55762 28592 55768
rect 29012 55282 29040 55898
rect 29000 55276 29052 55282
rect 29000 55218 29052 55224
rect 29104 54194 29132 56238
rect 30104 56228 30156 56234
rect 30104 56170 30156 56176
rect 29920 56160 29972 56166
rect 29920 56102 29972 56108
rect 29932 55758 29960 56102
rect 30116 55962 30144 56170
rect 30104 55956 30156 55962
rect 30104 55898 30156 55904
rect 29920 55752 29972 55758
rect 29920 55694 29972 55700
rect 29092 54188 29144 54194
rect 29092 54130 29144 54136
rect 28632 54120 28684 54126
rect 28632 54062 28684 54068
rect 28448 53780 28500 53786
rect 28448 53722 28500 53728
rect 28460 53446 28488 53722
rect 28644 53650 28672 54062
rect 29000 53984 29052 53990
rect 29000 53926 29052 53932
rect 29012 53802 29040 53926
rect 28920 53774 29040 53802
rect 28632 53644 28684 53650
rect 28632 53586 28684 53592
rect 28448 53440 28500 53446
rect 28448 53382 28500 53388
rect 28264 53236 28316 53242
rect 28264 53178 28316 53184
rect 27896 52896 27948 52902
rect 27896 52838 27948 52844
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22744 2644 22796 2650
rect 22744 2586 22796 2592
rect 22192 2372 22244 2378
rect 22192 2314 22244 2320
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21376 1902 21404 2246
rect 21364 1896 21416 1902
rect 21364 1838 21416 1844
rect 22204 800 22232 2314
rect 22848 2310 22876 2994
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 23032 2106 23060 2994
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 23492 2446 23520 2790
rect 23480 2440 23532 2446
rect 23308 2388 23480 2394
rect 23308 2382 23532 2388
rect 23308 2366 23520 2382
rect 24412 2378 24440 2790
rect 25516 2378 25544 2790
rect 24400 2372 24452 2378
rect 23020 2100 23072 2106
rect 23020 2042 23072 2048
rect 23308 800 23336 2366
rect 24400 2314 24452 2320
rect 25504 2372 25556 2378
rect 25504 2314 25556 2320
rect 24412 800 24440 2314
rect 25516 800 25544 2314
rect 26608 2304 26660 2310
rect 26608 2246 26660 2252
rect 26620 800 26648 2246
rect 27724 800 27752 2790
rect 27908 2514 27936 52838
rect 28644 2650 28672 53586
rect 28920 53582 28948 53774
rect 30116 53718 30144 55898
rect 30288 55888 30340 55894
rect 30288 55830 30340 55836
rect 30196 55752 30248 55758
rect 30196 55694 30248 55700
rect 30104 53712 30156 53718
rect 30104 53654 30156 53660
rect 28908 53576 28960 53582
rect 28908 53518 28960 53524
rect 29736 53576 29788 53582
rect 29736 53518 29788 53524
rect 30012 53576 30064 53582
rect 30012 53518 30064 53524
rect 28920 53106 28948 53518
rect 29748 53242 29776 53518
rect 29736 53236 29788 53242
rect 29736 53178 29788 53184
rect 30024 53106 30052 53518
rect 30208 53242 30236 55694
rect 30196 53236 30248 53242
rect 30196 53178 30248 53184
rect 28908 53100 28960 53106
rect 28908 53042 28960 53048
rect 30012 53100 30064 53106
rect 30012 53042 30064 53048
rect 28920 52902 28948 53042
rect 28908 52896 28960 52902
rect 28908 52838 28960 52844
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 28920 3194 28948 4014
rect 30024 3194 30052 4082
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 27896 2508 27948 2514
rect 27896 2450 27948 2456
rect 28920 2446 28948 3130
rect 30024 2446 30052 3130
rect 30300 3126 30328 55830
rect 31312 55622 31340 56306
rect 31496 55758 31524 56306
rect 32968 55962 32996 56306
rect 32956 55956 33008 55962
rect 32956 55898 33008 55904
rect 32968 55758 32996 55898
rect 33152 55758 33180 57258
rect 33232 57248 33284 57254
rect 33232 57190 33284 57196
rect 34796 57248 34848 57254
rect 34796 57190 34848 57196
rect 31484 55752 31536 55758
rect 31484 55694 31536 55700
rect 32956 55752 33008 55758
rect 32956 55694 33008 55700
rect 33140 55752 33192 55758
rect 33140 55694 33192 55700
rect 30840 55616 30892 55622
rect 30840 55558 30892 55564
rect 31300 55616 31352 55622
rect 31300 55558 31352 55564
rect 30852 55418 30880 55558
rect 30840 55412 30892 55418
rect 30840 55354 30892 55360
rect 32680 55276 32732 55282
rect 32680 55218 32732 55224
rect 31852 55208 31904 55214
rect 31852 55150 31904 55156
rect 31864 54194 31892 55150
rect 32404 55072 32456 55078
rect 32404 55014 32456 55020
rect 32416 54670 32444 55014
rect 32404 54664 32456 54670
rect 32404 54606 32456 54612
rect 32312 54528 32364 54534
rect 32312 54470 32364 54476
rect 32324 54330 32352 54470
rect 32312 54324 32364 54330
rect 32312 54266 32364 54272
rect 31852 54188 31904 54194
rect 31852 54130 31904 54136
rect 30472 54052 30524 54058
rect 30472 53994 30524 54000
rect 30484 53582 30512 53994
rect 31864 53582 31892 54130
rect 32324 54058 32352 54266
rect 32416 54058 32444 54606
rect 32312 54052 32364 54058
rect 32312 53994 32364 54000
rect 32404 54052 32456 54058
rect 32404 53994 32456 54000
rect 32416 53582 32444 53994
rect 32692 53990 32720 55218
rect 32772 54528 32824 54534
rect 32772 54470 32824 54476
rect 32784 54194 32812 54470
rect 32968 54194 32996 55694
rect 33244 54806 33272 57190
rect 33508 56364 33560 56370
rect 33508 56306 33560 56312
rect 33414 56264 33470 56273
rect 33414 56199 33416 56208
rect 33468 56199 33470 56208
rect 33416 56170 33468 56176
rect 33324 56160 33376 56166
rect 33324 56102 33376 56108
rect 33232 54800 33284 54806
rect 33232 54742 33284 54748
rect 32772 54188 32824 54194
rect 32772 54130 32824 54136
rect 32956 54188 33008 54194
rect 32956 54130 33008 54136
rect 32680 53984 32732 53990
rect 32680 53926 32732 53932
rect 32692 53650 32720 53926
rect 32680 53644 32732 53650
rect 32680 53586 32732 53592
rect 30472 53576 30524 53582
rect 30472 53518 30524 53524
rect 30564 53576 30616 53582
rect 30564 53518 30616 53524
rect 31852 53576 31904 53582
rect 31852 53518 31904 53524
rect 32404 53576 32456 53582
rect 32404 53518 32456 53524
rect 30484 52902 30512 53518
rect 30576 53174 30604 53518
rect 30932 53508 30984 53514
rect 30932 53450 30984 53456
rect 30564 53168 30616 53174
rect 30564 53110 30616 53116
rect 30472 52896 30524 52902
rect 30472 52838 30524 52844
rect 30944 3194 30972 53450
rect 31864 53106 31892 53518
rect 31944 53440 31996 53446
rect 31944 53382 31996 53388
rect 31956 53242 31984 53382
rect 31944 53236 31996 53242
rect 31944 53178 31996 53184
rect 31852 53100 31904 53106
rect 31852 53042 31904 53048
rect 33336 3194 33364 56102
rect 33520 55758 33548 56306
rect 33508 55752 33560 55758
rect 33508 55694 33560 55700
rect 34612 55752 34664 55758
rect 34612 55694 34664 55700
rect 34520 55616 34572 55622
rect 34520 55558 34572 55564
rect 34532 54738 34560 55558
rect 34520 54732 34572 54738
rect 34520 54674 34572 54680
rect 34624 54058 34652 55694
rect 34808 55690 34836 57190
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 35360 57050 35388 57394
rect 36556 57338 36584 57394
rect 36464 57310 36584 57338
rect 37648 57316 37700 57322
rect 35440 57248 35492 57254
rect 35440 57190 35492 57196
rect 35348 57044 35400 57050
rect 35348 56986 35400 56992
rect 35164 56500 35216 56506
rect 35164 56442 35216 56448
rect 35176 56409 35204 56442
rect 35452 56438 35480 57190
rect 36464 57050 36492 57310
rect 37648 57258 37700 57264
rect 36544 57248 36596 57254
rect 36544 57190 36596 57196
rect 37188 57248 37240 57254
rect 37188 57190 37240 57196
rect 36452 57044 36504 57050
rect 36452 56986 36504 56992
rect 35900 56704 35952 56710
rect 35900 56646 35952 56652
rect 35440 56432 35492 56438
rect 35162 56400 35218 56409
rect 35440 56374 35492 56380
rect 35806 56400 35862 56409
rect 35162 56335 35218 56344
rect 35348 56364 35400 56370
rect 35348 56306 35400 56312
rect 35532 56364 35584 56370
rect 35532 56306 35584 56312
rect 35716 56364 35768 56370
rect 35806 56335 35808 56344
rect 35716 56306 35768 56312
rect 35860 56335 35862 56344
rect 35808 56306 35860 56312
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 35072 55956 35124 55962
rect 35072 55898 35124 55904
rect 35084 55758 35112 55898
rect 35360 55758 35388 56306
rect 35072 55752 35124 55758
rect 35072 55694 35124 55700
rect 35348 55752 35400 55758
rect 35348 55694 35400 55700
rect 34796 55684 34848 55690
rect 34796 55626 34848 55632
rect 35256 55684 35308 55690
rect 35256 55626 35308 55632
rect 35268 55350 35296 55626
rect 35256 55344 35308 55350
rect 35256 55286 35308 55292
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 35360 54670 35388 55694
rect 35544 55622 35572 56306
rect 35728 56166 35756 56306
rect 35716 56160 35768 56166
rect 35716 56102 35768 56108
rect 35820 55758 35848 56306
rect 35808 55752 35860 55758
rect 35808 55694 35860 55700
rect 35532 55616 35584 55622
rect 35532 55558 35584 55564
rect 35820 54670 35848 55694
rect 35912 55690 35940 56646
rect 36266 56536 36322 56545
rect 36266 56471 36322 56480
rect 36280 56234 36308 56471
rect 36556 56438 36584 57190
rect 36544 56432 36596 56438
rect 36544 56374 36596 56380
rect 36910 56400 36966 56409
rect 36452 56364 36504 56370
rect 36452 56306 36504 56312
rect 36636 56364 36688 56370
rect 36910 56335 36912 56344
rect 36636 56306 36688 56312
rect 36964 56335 36966 56344
rect 36912 56306 36964 56312
rect 36268 56228 36320 56234
rect 36268 56170 36320 56176
rect 36464 55962 36492 56306
rect 36648 56234 36676 56306
rect 36728 56296 36780 56302
rect 36728 56238 36780 56244
rect 36636 56228 36688 56234
rect 36636 56170 36688 56176
rect 36452 55956 36504 55962
rect 36452 55898 36504 55904
rect 36740 55758 36768 56238
rect 37200 55826 37228 57190
rect 37188 55820 37240 55826
rect 37188 55762 37240 55768
rect 36544 55752 36596 55758
rect 36544 55694 36596 55700
rect 36728 55752 36780 55758
rect 36728 55694 36780 55700
rect 36820 55752 36872 55758
rect 36820 55694 36872 55700
rect 35900 55684 35952 55690
rect 35900 55626 35952 55632
rect 36556 55282 36584 55694
rect 36544 55276 36596 55282
rect 36544 55218 36596 55224
rect 35348 54664 35400 54670
rect 35348 54606 35400 54612
rect 35716 54664 35768 54670
rect 35716 54606 35768 54612
rect 35808 54664 35860 54670
rect 35808 54606 35860 54612
rect 35728 54330 35756 54606
rect 35716 54324 35768 54330
rect 35716 54266 35768 54272
rect 35820 54058 35848 54606
rect 36452 54528 36504 54534
rect 36452 54470 36504 54476
rect 36464 54194 36492 54470
rect 36740 54262 36768 55694
rect 36832 55078 36860 55694
rect 36820 55072 36872 55078
rect 36820 55014 36872 55020
rect 36832 54262 36860 55014
rect 36728 54256 36780 54262
rect 36728 54198 36780 54204
rect 36820 54256 36872 54262
rect 36820 54198 36872 54204
rect 36452 54188 36504 54194
rect 36452 54130 36504 54136
rect 36740 54126 36768 54198
rect 37660 54194 37688 57258
rect 38948 57050 38976 57394
rect 40040 57384 40092 57390
rect 40040 57326 40092 57332
rect 39028 57248 39080 57254
rect 39028 57190 39080 57196
rect 38936 57044 38988 57050
rect 38936 56986 38988 56992
rect 38660 56772 38712 56778
rect 38660 56714 38712 56720
rect 38384 56500 38436 56506
rect 38384 56442 38436 56448
rect 38200 56432 38252 56438
rect 38200 56374 38252 56380
rect 38212 55962 38240 56374
rect 38396 56273 38424 56442
rect 38672 56370 38700 56714
rect 39040 56438 39068 57190
rect 39212 56840 39264 56846
rect 39212 56782 39264 56788
rect 39304 56840 39356 56846
rect 39304 56782 39356 56788
rect 39224 56438 39252 56782
rect 39028 56432 39080 56438
rect 39028 56374 39080 56380
rect 39212 56432 39264 56438
rect 39212 56374 39264 56380
rect 39316 56370 39344 56782
rect 39580 56772 39632 56778
rect 39580 56714 39632 56720
rect 39592 56370 39620 56714
rect 38660 56364 38712 56370
rect 38660 56306 38712 56312
rect 38844 56364 38896 56370
rect 38844 56306 38896 56312
rect 39304 56364 39356 56370
rect 39304 56306 39356 56312
rect 39580 56364 39632 56370
rect 39580 56306 39632 56312
rect 38382 56264 38438 56273
rect 38382 56199 38438 56208
rect 38200 55956 38252 55962
rect 38200 55898 38252 55904
rect 37924 55616 37976 55622
rect 37924 55558 37976 55564
rect 37740 55276 37792 55282
rect 37740 55218 37792 55224
rect 37752 54330 37780 55218
rect 37936 54534 37964 55558
rect 38672 55282 38700 56306
rect 38752 55752 38804 55758
rect 38752 55694 38804 55700
rect 38764 55622 38792 55694
rect 38752 55616 38804 55622
rect 38752 55558 38804 55564
rect 38856 55604 38884 56306
rect 38936 56296 38988 56302
rect 38936 56238 38988 56244
rect 38948 55736 38976 56238
rect 40052 55826 40080 57326
rect 40500 57316 40552 57322
rect 40500 57258 40552 57264
rect 40512 56370 40540 57258
rect 41340 57050 41368 57394
rect 41420 57248 41472 57254
rect 41420 57190 41472 57196
rect 42800 57248 42852 57254
rect 42800 57190 42852 57196
rect 41328 57044 41380 57050
rect 41328 56986 41380 56992
rect 41432 56914 41460 57190
rect 42708 56976 42760 56982
rect 42708 56918 42760 56924
rect 41420 56908 41472 56914
rect 41420 56850 41472 56856
rect 40500 56364 40552 56370
rect 40500 56306 40552 56312
rect 41696 56364 41748 56370
rect 41696 56306 41748 56312
rect 42156 56364 42208 56370
rect 42156 56306 42208 56312
rect 41512 56296 41564 56302
rect 41512 56238 41564 56244
rect 41708 56250 41736 56306
rect 41236 56160 41288 56166
rect 41236 56102 41288 56108
rect 41248 55894 41276 56102
rect 41236 55888 41288 55894
rect 41236 55830 41288 55836
rect 40040 55820 40092 55826
rect 40040 55762 40092 55768
rect 41524 55758 41552 56238
rect 41708 56222 41920 56250
rect 41892 55894 41920 56222
rect 42168 55962 42196 56306
rect 42156 55956 42208 55962
rect 42156 55898 42208 55904
rect 41880 55888 41932 55894
rect 41880 55830 41932 55836
rect 39028 55752 39080 55758
rect 38936 55730 38988 55736
rect 39028 55694 39080 55700
rect 41512 55752 41564 55758
rect 41512 55694 41564 55700
rect 38936 55672 38988 55678
rect 39040 55604 39068 55694
rect 38856 55576 39068 55604
rect 38660 55276 38712 55282
rect 38660 55218 38712 55224
rect 37924 54528 37976 54534
rect 37924 54470 37976 54476
rect 38568 54528 38620 54534
rect 38568 54470 38620 54476
rect 37740 54324 37792 54330
rect 37740 54266 37792 54272
rect 37752 54194 37780 54266
rect 38580 54194 38608 54470
rect 38660 54256 38712 54262
rect 38856 54244 38884 55576
rect 41052 55412 41104 55418
rect 41052 55354 41104 55360
rect 40040 55276 40092 55282
rect 40040 55218 40092 55224
rect 40052 54670 40080 55218
rect 40316 55072 40368 55078
rect 40316 55014 40368 55020
rect 40868 55072 40920 55078
rect 40868 55014 40920 55020
rect 40328 54874 40356 55014
rect 40316 54868 40368 54874
rect 40316 54810 40368 54816
rect 40040 54664 40092 54670
rect 40040 54606 40092 54612
rect 39396 54528 39448 54534
rect 39396 54470 39448 54476
rect 39408 54262 39436 54470
rect 38712 54216 38884 54244
rect 39396 54256 39448 54262
rect 38660 54198 38712 54204
rect 39396 54198 39448 54204
rect 37648 54188 37700 54194
rect 37648 54130 37700 54136
rect 37740 54188 37792 54194
rect 37740 54130 37792 54136
rect 38568 54188 38620 54194
rect 38568 54130 38620 54136
rect 36728 54120 36780 54126
rect 36728 54062 36780 54068
rect 34612 54052 34664 54058
rect 34612 53994 34664 54000
rect 35808 54052 35860 54058
rect 35808 53994 35860 54000
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 36740 53786 36768 54062
rect 38672 53786 38700 54198
rect 36728 53780 36780 53786
rect 36728 53722 36780 53728
rect 38660 53780 38712 53786
rect 38660 53722 38712 53728
rect 39408 53582 39436 54198
rect 40052 53990 40080 54606
rect 40328 54194 40356 54810
rect 40880 54602 40908 55014
rect 41064 54874 41092 55354
rect 41524 54874 41552 55694
rect 41892 55690 41920 55830
rect 42168 55758 42196 55898
rect 42156 55752 42208 55758
rect 42156 55694 42208 55700
rect 41880 55684 41932 55690
rect 41880 55626 41932 55632
rect 41052 54868 41104 54874
rect 41052 54810 41104 54816
rect 41328 54868 41380 54874
rect 41328 54810 41380 54816
rect 41512 54868 41564 54874
rect 41512 54810 41564 54816
rect 40868 54596 40920 54602
rect 40868 54538 40920 54544
rect 41064 54534 41092 54810
rect 41052 54528 41104 54534
rect 41052 54470 41104 54476
rect 40316 54188 40368 54194
rect 40316 54130 40368 54136
rect 40040 53984 40092 53990
rect 40040 53926 40092 53932
rect 39396 53576 39448 53582
rect 39396 53518 39448 53524
rect 40052 53514 40080 53926
rect 40328 53786 40356 54130
rect 41340 53990 41368 54810
rect 41892 54330 41920 55626
rect 42168 54806 42196 55694
rect 42720 55622 42748 56918
rect 42812 56302 42840 57190
rect 42800 56296 42852 56302
rect 42800 56238 42852 56244
rect 42904 55690 42932 57462
rect 43732 57458 43760 59200
rect 44928 57458 44956 59200
rect 45468 57588 45520 57594
rect 45468 57530 45520 57536
rect 43720 57452 43772 57458
rect 43720 57394 43772 57400
rect 44916 57452 44968 57458
rect 44916 57394 44968 57400
rect 44272 57384 44324 57390
rect 44272 57326 44324 57332
rect 44180 57316 44232 57322
rect 44180 57258 44232 57264
rect 43536 56840 43588 56846
rect 43536 56782 43588 56788
rect 44088 56840 44140 56846
rect 44088 56782 44140 56788
rect 43444 56704 43496 56710
rect 43444 56646 43496 56652
rect 43456 56506 43484 56646
rect 43444 56500 43496 56506
rect 43444 56442 43496 56448
rect 43548 56386 43576 56782
rect 43812 56772 43864 56778
rect 43812 56714 43864 56720
rect 43824 56386 43852 56714
rect 43456 56370 43576 56386
rect 43640 56370 43852 56386
rect 44100 56370 44128 56782
rect 43444 56364 43576 56370
rect 43496 56358 43576 56364
rect 43628 56364 43852 56370
rect 43444 56306 43496 56312
rect 43680 56358 43852 56364
rect 43904 56364 43956 56370
rect 43628 56306 43680 56312
rect 43904 56306 43956 56312
rect 44088 56364 44140 56370
rect 44088 56306 44140 56312
rect 43456 55758 43484 56306
rect 43640 55894 43668 56306
rect 43916 55962 43944 56306
rect 43904 55956 43956 55962
rect 43904 55898 43956 55904
rect 43628 55888 43680 55894
rect 43628 55830 43680 55836
rect 43444 55752 43496 55758
rect 43444 55694 43496 55700
rect 42892 55684 42944 55690
rect 42892 55626 42944 55632
rect 42708 55616 42760 55622
rect 42708 55558 42760 55564
rect 43260 55616 43312 55622
rect 43260 55558 43312 55564
rect 42156 54800 42208 54806
rect 42156 54742 42208 54748
rect 43272 54670 43300 55558
rect 43456 55282 43484 55694
rect 43640 55298 43668 55830
rect 43916 55758 43944 55898
rect 43904 55752 43956 55758
rect 43956 55700 44036 55706
rect 43904 55694 44036 55700
rect 43916 55678 44036 55694
rect 43640 55282 43760 55298
rect 44008 55282 44036 55678
rect 44192 55282 44220 57258
rect 44284 56234 44312 57326
rect 44928 57050 44956 57394
rect 44916 57044 44968 57050
rect 44916 56986 44968 56992
rect 44272 56228 44324 56234
rect 44272 56170 44324 56176
rect 45480 55826 45508 57530
rect 46124 57458 46152 59200
rect 47320 57458 47348 59200
rect 48516 57458 48544 59200
rect 49712 57458 49740 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50436 57588 50488 57594
rect 50436 57530 50488 57536
rect 46112 57452 46164 57458
rect 46112 57394 46164 57400
rect 47308 57452 47360 57458
rect 47308 57394 47360 57400
rect 48504 57452 48556 57458
rect 48504 57394 48556 57400
rect 49700 57452 49752 57458
rect 49700 57394 49752 57400
rect 50344 57452 50396 57458
rect 50344 57394 50396 57400
rect 46204 57248 46256 57254
rect 46204 57190 46256 57196
rect 46216 56914 46244 57190
rect 47320 57050 47348 57394
rect 50356 57050 50384 57394
rect 47308 57044 47360 57050
rect 47308 56986 47360 56992
rect 50344 57044 50396 57050
rect 50344 56986 50396 56992
rect 50448 56982 50476 57530
rect 50908 57474 50936 59200
rect 50908 57458 51120 57474
rect 52104 57458 52132 59200
rect 53300 57458 53328 59200
rect 54496 57458 54524 59200
rect 55692 57458 55720 59200
rect 56888 57458 56916 59200
rect 57518 58984 57574 58993
rect 57518 58919 57574 58928
rect 50908 57452 51132 57458
rect 50908 57446 51080 57452
rect 51080 57394 51132 57400
rect 52092 57452 52144 57458
rect 52092 57394 52144 57400
rect 53288 57452 53340 57458
rect 53288 57394 53340 57400
rect 54484 57452 54536 57458
rect 54484 57394 54536 57400
rect 55680 57452 55732 57458
rect 55680 57394 55732 57400
rect 56876 57452 56928 57458
rect 56876 57394 56928 57400
rect 52104 57050 52132 57394
rect 52184 57248 52236 57254
rect 52184 57190 52236 57196
rect 53380 57248 53432 57254
rect 53380 57190 53432 57196
rect 52092 57044 52144 57050
rect 52092 56986 52144 56992
rect 50436 56976 50488 56982
rect 50436 56918 50488 56924
rect 46204 56908 46256 56914
rect 46204 56850 46256 56856
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 52196 56438 52224 57190
rect 53392 56710 53420 57190
rect 54496 57050 54524 57394
rect 54576 57248 54628 57254
rect 54576 57190 54628 57196
rect 54668 57248 54720 57254
rect 54668 57190 54720 57196
rect 54484 57044 54536 57050
rect 54484 56986 54536 56992
rect 53380 56704 53432 56710
rect 53380 56646 53432 56652
rect 52184 56432 52236 56438
rect 52184 56374 52236 56380
rect 45468 55820 45520 55826
rect 45468 55762 45520 55768
rect 54588 55622 54616 57190
rect 54576 55616 54628 55622
rect 54576 55558 54628 55564
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 54680 55350 54708 57190
rect 56888 57050 56916 57394
rect 57058 57352 57114 57361
rect 57058 57287 57114 57296
rect 56876 57044 56928 57050
rect 56876 56986 56928 56992
rect 57072 56846 57100 57287
rect 57532 56846 57560 58919
rect 58084 57458 58112 59200
rect 58438 58168 58494 58177
rect 58438 58103 58494 58112
rect 58072 57452 58124 57458
rect 58072 57394 58124 57400
rect 57060 56840 57112 56846
rect 57060 56782 57112 56788
rect 57520 56840 57572 56846
rect 58084 56794 58112 57394
rect 58164 57248 58216 57254
rect 58164 57190 58216 57196
rect 57520 56782 57572 56788
rect 56784 56704 56836 56710
rect 56784 56646 56836 56652
rect 54668 55344 54720 55350
rect 54668 55286 54720 55292
rect 43444 55276 43496 55282
rect 43640 55276 43772 55282
rect 43640 55270 43720 55276
rect 43444 55218 43496 55224
rect 43720 55218 43772 55224
rect 43996 55276 44048 55282
rect 43996 55218 44048 55224
rect 44180 55276 44232 55282
rect 44180 55218 44232 55224
rect 43260 54664 43312 54670
rect 43260 54606 43312 54612
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 41880 54324 41932 54330
rect 41880 54266 41932 54272
rect 41328 53984 41380 53990
rect 41328 53926 41380 53932
rect 40316 53780 40368 53786
rect 40316 53722 40368 53728
rect 38384 53508 38436 53514
rect 38384 53450 38436 53456
rect 40040 53508 40092 53514
rect 40040 53450 40092 53456
rect 38396 52902 38424 53450
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 38384 52896 38436 52902
rect 38384 52838 38436 52844
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 30932 3188 30984 3194
rect 30932 3130 30984 3136
rect 33324 3188 33376 3194
rect 33324 3130 33376 3136
rect 30288 3120 30340 3126
rect 30288 3062 30340 3068
rect 30944 2446 30972 3130
rect 32312 3120 32364 3126
rect 32312 3062 32364 3068
rect 32324 2446 32352 3062
rect 33336 2446 33364 3130
rect 37740 3120 37792 3126
rect 37740 3062 37792 3068
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 36004 2446 36032 2790
rect 37752 2446 37780 3062
rect 38396 2582 38424 52838
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 55956 47456 56008 47462
rect 55956 47398 56008 47404
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 55680 39296 55732 39302
rect 55680 39238 55732 39244
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 55496 38548 55548 38554
rect 55496 38490 55548 38496
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 55508 37874 55536 38490
rect 55496 37868 55548 37874
rect 55496 37810 55548 37816
rect 54668 37664 54720 37670
rect 54668 37606 54720 37612
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 53932 35284 53984 35290
rect 53932 35226 53984 35232
rect 52368 35012 52420 35018
rect 52368 34954 52420 34960
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 52380 34610 52408 34954
rect 53944 34746 53972 35226
rect 54576 35080 54628 35086
rect 54576 35022 54628 35028
rect 53932 34740 53984 34746
rect 53932 34682 53984 34688
rect 52368 34604 52420 34610
rect 52368 34546 52420 34552
rect 51448 34536 51500 34542
rect 51448 34478 51500 34484
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 49056 32360 49108 32366
rect 49056 32302 49108 32308
rect 44364 26240 44416 26246
rect 44364 26182 44416 26188
rect 40868 9716 40920 9722
rect 40868 9658 40920 9664
rect 40880 3738 40908 9658
rect 40868 3732 40920 3738
rect 40868 3674 40920 3680
rect 40880 3534 40908 3674
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 40316 3392 40368 3398
rect 40316 3334 40368 3340
rect 38660 2984 38712 2990
rect 38660 2926 38712 2932
rect 38384 2576 38436 2582
rect 38384 2518 38436 2524
rect 38672 2446 38700 2926
rect 39212 2916 39264 2922
rect 39212 2858 39264 2864
rect 39224 2446 39252 2858
rect 40328 2446 40356 3334
rect 44376 3194 44404 26182
rect 45836 18624 45888 18630
rect 45836 18566 45888 18572
rect 44824 6180 44876 6186
rect 44824 6122 44876 6128
rect 44836 3194 44864 6122
rect 45848 3194 45876 18566
rect 48044 3392 48096 3398
rect 48044 3334 48096 3340
rect 43628 3188 43680 3194
rect 43628 3130 43680 3136
rect 44364 3188 44416 3194
rect 44364 3130 44416 3136
rect 44824 3188 44876 3194
rect 44824 3130 44876 3136
rect 45836 3188 45888 3194
rect 45836 3130 45888 3136
rect 43640 2446 43668 3130
rect 44836 2446 44864 3130
rect 45848 2446 45876 3130
rect 48056 2446 48084 3334
rect 49068 2446 49096 32302
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50160 9920 50212 9926
rect 50160 9862 50212 9868
rect 50172 9722 50200 9862
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50160 9716 50212 9722
rect 50160 9658 50212 9664
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 51460 3194 51488 34478
rect 53104 23112 53156 23118
rect 53104 23054 53156 23060
rect 51724 10464 51776 10470
rect 51724 10406 51776 10412
rect 51448 3188 51500 3194
rect 51448 3130 51500 3136
rect 50620 2848 50672 2854
rect 50620 2790 50672 2796
rect 50632 2446 50660 2790
rect 51460 2446 51488 3130
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 33324 2440 33376 2446
rect 35992 2440 36044 2446
rect 33324 2382 33376 2388
rect 35820 2400 35992 2428
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 29920 2304 29972 2310
rect 29920 2246 29972 2252
rect 31024 2304 31076 2310
rect 31024 2246 31076 2252
rect 32128 2304 32180 2310
rect 32128 2246 32180 2252
rect 33232 2304 33284 2310
rect 33232 2246 33284 2252
rect 34336 2304 34388 2310
rect 34336 2246 34388 2252
rect 28828 800 28856 2246
rect 29932 800 29960 2246
rect 31036 800 31064 2246
rect 32140 800 32168 2246
rect 33244 800 33272 2246
rect 34348 800 34376 2246
rect 35452 870 35572 898
rect 35452 800 35480 870
rect 2318 0 2374 800
rect 3422 0 3478 800
rect 4526 0 4582 800
rect 5630 0 5686 800
rect 6734 0 6790 800
rect 7838 0 7894 800
rect 8942 0 8998 800
rect 10046 0 10102 800
rect 11150 0 11206 800
rect 12254 0 12310 800
rect 13358 0 13414 800
rect 14462 0 14518 800
rect 15566 0 15622 800
rect 16670 0 16726 800
rect 17774 0 17830 800
rect 18878 0 18934 800
rect 19982 0 20038 800
rect 21086 0 21142 800
rect 22190 0 22246 800
rect 23294 0 23350 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26606 0 26662 800
rect 27710 0 27766 800
rect 28814 0 28870 800
rect 29918 0 29974 800
rect 31022 0 31078 800
rect 32126 0 32182 800
rect 33230 0 33286 800
rect 34334 0 34390 800
rect 35438 0 35494 800
rect 35544 762 35572 870
rect 35820 762 35848 2400
rect 35992 2382 36044 2388
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 39212 2440 39264 2446
rect 39212 2382 39264 2388
rect 40316 2440 40368 2446
rect 40316 2382 40368 2388
rect 43628 2440 43680 2446
rect 43628 2382 43680 2388
rect 44824 2440 44876 2446
rect 44824 2382 44876 2388
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 48044 2440 48096 2446
rect 48044 2382 48096 2388
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 50620 2440 50672 2446
rect 50620 2382 50672 2388
rect 51448 2440 51500 2446
rect 51448 2382 51500 2388
rect 36360 2372 36412 2378
rect 36360 2314 36412 2320
rect 36372 2106 36400 2314
rect 36544 2304 36596 2310
rect 36544 2246 36596 2252
rect 37648 2304 37700 2310
rect 37648 2246 37700 2252
rect 38752 2304 38804 2310
rect 38752 2246 38804 2252
rect 39856 2304 39908 2310
rect 39856 2246 39908 2252
rect 40960 2304 41012 2310
rect 40960 2246 41012 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 42064 2304 42116 2310
rect 42064 2246 42116 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 44272 2304 44324 2310
rect 44272 2246 44324 2252
rect 45376 2304 45428 2310
rect 45376 2246 45428 2252
rect 46480 2304 46532 2310
rect 46480 2246 46532 2252
rect 47584 2304 47636 2310
rect 47584 2246 47636 2252
rect 48688 2304 48740 2310
rect 48688 2246 48740 2252
rect 49792 2304 49844 2310
rect 49792 2246 49844 2252
rect 50896 2304 50948 2310
rect 50896 2246 50948 2252
rect 36360 2100 36412 2106
rect 36360 2042 36412 2048
rect 36556 800 36584 2246
rect 37660 800 37688 2246
rect 38764 800 38792 2246
rect 39868 800 39896 2246
rect 40972 800 41000 2246
rect 41892 2038 41920 2246
rect 41880 2032 41932 2038
rect 41880 1974 41932 1980
rect 42076 800 42104 2246
rect 43180 800 43208 2246
rect 44284 800 44312 2246
rect 45388 800 45416 2246
rect 46492 800 46520 2246
rect 47596 800 47624 2246
rect 48700 800 48728 2246
rect 49804 800 49832 2246
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50908 800 50936 2246
rect 51736 2038 51764 10406
rect 53116 6186 53144 23054
rect 53104 6180 53156 6186
rect 53104 6122 53156 6128
rect 53380 4004 53432 4010
rect 53380 3946 53432 3952
rect 53392 2446 53420 3946
rect 53748 3664 53800 3670
rect 53748 3606 53800 3612
rect 53760 3194 53788 3606
rect 54484 3392 54536 3398
rect 54484 3334 54536 3340
rect 53748 3188 53800 3194
rect 53748 3130 53800 3136
rect 54496 2446 54524 3334
rect 54588 2854 54616 35022
rect 54680 3534 54708 37606
rect 54760 35080 54812 35086
rect 54760 35022 54812 35028
rect 54772 34746 54800 35022
rect 54760 34740 54812 34746
rect 54760 34682 54812 34688
rect 55220 34740 55272 34746
rect 55220 34682 55272 34688
rect 55232 34610 55260 34682
rect 55220 34604 55272 34610
rect 55220 34546 55272 34552
rect 55588 34468 55640 34474
rect 55588 34410 55640 34416
rect 55600 34202 55628 34410
rect 55588 34196 55640 34202
rect 55588 34138 55640 34144
rect 55312 11552 55364 11558
rect 55312 11494 55364 11500
rect 55324 10674 55352 11494
rect 55312 10668 55364 10674
rect 55312 10610 55364 10616
rect 55404 9648 55456 9654
rect 55404 9590 55456 9596
rect 55312 3596 55364 3602
rect 55312 3538 55364 3544
rect 54668 3528 54720 3534
rect 54668 3470 54720 3476
rect 54680 3194 54708 3470
rect 54668 3188 54720 3194
rect 54668 3130 54720 3136
rect 54576 2848 54628 2854
rect 54576 2790 54628 2796
rect 55324 2689 55352 3538
rect 55310 2680 55366 2689
rect 55310 2615 55366 2624
rect 53380 2440 53432 2446
rect 53380 2382 53432 2388
rect 54484 2440 54536 2446
rect 54484 2382 54536 2388
rect 52000 2304 52052 2310
rect 52000 2246 52052 2252
rect 53104 2304 53156 2310
rect 53104 2246 53156 2252
rect 54208 2304 54260 2310
rect 54208 2246 54260 2252
rect 55312 2304 55364 2310
rect 55312 2246 55364 2252
rect 51724 2032 51776 2038
rect 51724 1974 51776 1980
rect 52012 800 52040 2246
rect 53116 800 53144 2246
rect 54220 800 54248 2246
rect 55324 800 55352 2246
rect 55416 2106 55444 9590
rect 55588 6656 55640 6662
rect 55588 6598 55640 6604
rect 55600 3602 55628 6598
rect 55692 4146 55720 39238
rect 55968 38010 55996 47398
rect 56692 39500 56744 39506
rect 56692 39442 56744 39448
rect 56232 39432 56284 39438
rect 56232 39374 56284 39380
rect 56140 39364 56192 39370
rect 56140 39306 56192 39312
rect 56152 39098 56180 39306
rect 56140 39092 56192 39098
rect 56140 39034 56192 39040
rect 56244 38554 56272 39374
rect 56704 38758 56732 39442
rect 56692 38752 56744 38758
rect 56692 38694 56744 38700
rect 56232 38548 56284 38554
rect 56232 38490 56284 38496
rect 55772 38004 55824 38010
rect 55772 37946 55824 37952
rect 55956 38004 56008 38010
rect 55956 37946 56008 37952
rect 55784 37754 55812 37946
rect 55784 37726 55904 37754
rect 55876 37670 55904 37726
rect 55864 37664 55916 37670
rect 55864 37606 55916 37612
rect 56244 37466 56272 38490
rect 56704 38418 56732 38694
rect 56692 38412 56744 38418
rect 56692 38354 56744 38360
rect 56600 38208 56652 38214
rect 56600 38150 56652 38156
rect 56232 37460 56284 37466
rect 56232 37402 56284 37408
rect 56244 37194 56272 37402
rect 56232 37188 56284 37194
rect 56232 37130 56284 37136
rect 56244 35290 56272 37130
rect 56612 35986 56640 38150
rect 56704 37806 56732 38354
rect 56796 38010 56824 56646
rect 57072 56506 57100 56782
rect 57060 56500 57112 56506
rect 57060 56442 57112 56448
rect 57532 56438 57560 56782
rect 57992 56766 58112 56794
rect 57888 56704 57940 56710
rect 57888 56646 57940 56652
rect 57520 56432 57572 56438
rect 57520 56374 57572 56380
rect 57900 45554 57928 56646
rect 57992 56370 58020 56766
rect 58072 56704 58124 56710
rect 58072 56646 58124 56652
rect 57980 56364 58032 56370
rect 57980 56306 58032 56312
rect 57980 55276 58032 55282
rect 57980 55218 58032 55224
rect 57992 54913 58020 55218
rect 57978 54904 58034 54913
rect 57978 54839 58034 54848
rect 57808 45526 57928 45554
rect 57244 45280 57296 45286
rect 57244 45222 57296 45228
rect 56968 42560 57020 42566
rect 56968 42502 57020 42508
rect 56980 41414 57008 42502
rect 56888 41386 57008 41414
rect 56784 38004 56836 38010
rect 56784 37946 56836 37952
rect 56796 37874 56824 37946
rect 56784 37868 56836 37874
rect 56784 37810 56836 37816
rect 56692 37800 56744 37806
rect 56692 37742 56744 37748
rect 56704 37330 56732 37742
rect 56692 37324 56744 37330
rect 56692 37266 56744 37272
rect 56704 36922 56732 37266
rect 56692 36916 56744 36922
rect 56692 36858 56744 36864
rect 56428 35958 56640 35986
rect 56232 35284 56284 35290
rect 56232 35226 56284 35232
rect 56048 34536 56100 34542
rect 56048 34478 56100 34484
rect 55864 32768 55916 32774
rect 55864 32710 55916 32716
rect 55876 32434 55904 32710
rect 55864 32428 55916 32434
rect 55864 32370 55916 32376
rect 55956 32224 56008 32230
rect 55956 32166 56008 32172
rect 55772 11552 55824 11558
rect 55772 11494 55824 11500
rect 55784 6662 55812 11494
rect 55772 6656 55824 6662
rect 55772 6598 55824 6604
rect 55680 4140 55732 4146
rect 55680 4082 55732 4088
rect 55588 3596 55640 3602
rect 55588 3538 55640 3544
rect 55692 3534 55720 4082
rect 55968 3738 55996 32166
rect 56060 26042 56088 34478
rect 56244 33658 56272 35226
rect 56232 33652 56284 33658
rect 56232 33594 56284 33600
rect 56140 33108 56192 33114
rect 56140 33050 56192 33056
rect 56048 26036 56100 26042
rect 56048 25978 56100 25984
rect 56152 16574 56180 33050
rect 56244 32978 56272 33594
rect 56232 32972 56284 32978
rect 56232 32914 56284 32920
rect 56244 32434 56272 32914
rect 56232 32428 56284 32434
rect 56232 32370 56284 32376
rect 56244 32026 56272 32370
rect 56232 32020 56284 32026
rect 56232 31962 56284 31968
rect 56060 16546 56180 16574
rect 56060 13870 56088 16546
rect 56048 13864 56100 13870
rect 56048 13806 56100 13812
rect 55956 3732 56008 3738
rect 55956 3674 56008 3680
rect 55680 3528 55732 3534
rect 55680 3470 55732 3476
rect 55496 3392 55548 3398
rect 55496 3334 55548 3340
rect 55508 2446 55536 3334
rect 56060 3210 56088 13806
rect 56140 13184 56192 13190
rect 56140 13126 56192 13132
rect 56152 4078 56180 13126
rect 56244 9654 56272 31962
rect 56428 16574 56456 35958
rect 56704 35834 56732 36858
rect 56692 35828 56744 35834
rect 56692 35770 56744 35776
rect 56704 34474 56732 35770
rect 56692 34468 56744 34474
rect 56692 34410 56744 34416
rect 56600 34128 56652 34134
rect 56600 34070 56652 34076
rect 56612 32502 56640 34070
rect 56704 33658 56732 34410
rect 56692 33652 56744 33658
rect 56692 33594 56744 33600
rect 56704 33114 56732 33594
rect 56692 33108 56744 33114
rect 56692 33050 56744 33056
rect 56600 32496 56652 32502
rect 56600 32438 56652 32444
rect 56704 32366 56732 33050
rect 56692 32360 56744 32366
rect 56692 32302 56744 32308
rect 56888 30954 56916 41386
rect 56968 37392 57020 37398
rect 56968 37334 57020 37340
rect 56980 34474 57008 37334
rect 57152 35284 57204 35290
rect 57152 35226 57204 35232
rect 57164 35154 57192 35226
rect 57152 35148 57204 35154
rect 57152 35090 57204 35096
rect 57256 34746 57284 45222
rect 57336 40384 57388 40390
rect 57336 40326 57388 40332
rect 57244 34740 57296 34746
rect 57244 34682 57296 34688
rect 56968 34468 57020 34474
rect 56968 34410 57020 34416
rect 56968 32564 57020 32570
rect 56968 32506 57020 32512
rect 56980 31754 57008 32506
rect 56980 31726 57192 31754
rect 56888 30926 57008 30954
rect 56980 30598 57008 30926
rect 57060 30660 57112 30666
rect 57060 30602 57112 30608
rect 56784 30592 56836 30598
rect 56784 30534 56836 30540
rect 56968 30592 57020 30598
rect 56968 30534 57020 30540
rect 56692 24676 56744 24682
rect 56692 24618 56744 24624
rect 56600 19508 56652 19514
rect 56600 19450 56652 19456
rect 56428 16546 56548 16574
rect 56324 11892 56376 11898
rect 56324 11834 56376 11840
rect 56336 11762 56364 11834
rect 56324 11756 56376 11762
rect 56324 11698 56376 11704
rect 56232 9648 56284 9654
rect 56232 9590 56284 9596
rect 56324 6996 56376 7002
rect 56324 6938 56376 6944
rect 56336 6866 56364 6938
rect 56324 6860 56376 6866
rect 56324 6802 56376 6808
rect 56416 6792 56468 6798
rect 56416 6734 56468 6740
rect 56428 6662 56456 6734
rect 56416 6656 56468 6662
rect 56416 6598 56468 6604
rect 56520 4826 56548 16546
rect 56612 11762 56640 19450
rect 56704 14006 56732 24618
rect 56796 22778 56824 30534
rect 56876 30048 56928 30054
rect 56876 29990 56928 29996
rect 56888 29714 56916 29990
rect 56876 29708 56928 29714
rect 56876 29650 56928 29656
rect 56888 28422 56916 29650
rect 56876 28416 56928 28422
rect 56876 28358 56928 28364
rect 56784 22772 56836 22778
rect 56784 22714 56836 22720
rect 57072 22094 57100 30602
rect 57164 28506 57192 31726
rect 57244 30660 57296 30666
rect 57244 30602 57296 30608
rect 57256 30054 57284 30602
rect 57244 30048 57296 30054
rect 57244 29990 57296 29996
rect 57244 29640 57296 29646
rect 57244 29582 57296 29588
rect 57256 29102 57284 29582
rect 57244 29096 57296 29102
rect 57244 29038 57296 29044
rect 57164 28478 57284 28506
rect 57152 28416 57204 28422
rect 57152 28358 57204 28364
rect 57164 26790 57192 28358
rect 57152 26784 57204 26790
rect 57152 26726 57204 26732
rect 57164 26382 57192 26726
rect 57152 26376 57204 26382
rect 57152 26318 57204 26324
rect 57164 25294 57192 26318
rect 57152 25288 57204 25294
rect 57152 25230 57204 25236
rect 57164 24614 57192 25230
rect 57152 24608 57204 24614
rect 57152 24550 57204 24556
rect 57256 24342 57284 28478
rect 57348 26450 57376 40326
rect 57428 39296 57480 39302
rect 57428 39238 57480 39244
rect 57612 39296 57664 39302
rect 57612 39238 57664 39244
rect 57440 37346 57468 39238
rect 57520 38752 57572 38758
rect 57520 38694 57572 38700
rect 57532 37874 57560 38694
rect 57624 38350 57652 39238
rect 57808 38842 57836 45526
rect 57980 44328 58032 44334
rect 57980 44270 58032 44276
rect 57888 39840 57940 39846
rect 57888 39782 57940 39788
rect 57900 38962 57928 39782
rect 57992 39642 58020 44270
rect 57980 39636 58032 39642
rect 57980 39578 58032 39584
rect 57888 38956 57940 38962
rect 57888 38898 57940 38904
rect 57808 38814 57928 38842
rect 57900 38350 57928 38814
rect 57612 38344 57664 38350
rect 57612 38286 57664 38292
rect 57888 38344 57940 38350
rect 57888 38286 57940 38292
rect 57980 38276 58032 38282
rect 57980 38218 58032 38224
rect 57888 38004 57940 38010
rect 57888 37946 57940 37952
rect 57520 37868 57572 37874
rect 57520 37810 57572 37816
rect 57440 37318 57836 37346
rect 57428 37188 57480 37194
rect 57428 37130 57480 37136
rect 57440 36922 57468 37130
rect 57428 36916 57480 36922
rect 57428 36858 57480 36864
rect 57704 36032 57756 36038
rect 57704 35974 57756 35980
rect 57428 35828 57480 35834
rect 57428 35770 57480 35776
rect 57440 35170 57468 35770
rect 57716 35698 57744 35974
rect 57704 35692 57756 35698
rect 57704 35634 57756 35640
rect 57612 35488 57664 35494
rect 57612 35430 57664 35436
rect 57440 35154 57560 35170
rect 57440 35148 57572 35154
rect 57440 35142 57520 35148
rect 57520 35090 57572 35096
rect 57624 34678 57652 35430
rect 57612 34672 57664 34678
rect 57612 34614 57664 34620
rect 57520 34468 57572 34474
rect 57520 34410 57572 34416
rect 57428 33652 57480 33658
rect 57428 33594 57480 33600
rect 57440 32910 57468 33594
rect 57428 32904 57480 32910
rect 57428 32846 57480 32852
rect 57532 31754 57560 34410
rect 57704 33108 57756 33114
rect 57704 33050 57756 33056
rect 57716 32978 57744 33050
rect 57704 32972 57756 32978
rect 57704 32914 57756 32920
rect 57532 31726 57744 31754
rect 57612 30796 57664 30802
rect 57612 30738 57664 30744
rect 57624 30054 57652 30738
rect 57612 30048 57664 30054
rect 57612 29990 57664 29996
rect 57624 29714 57652 29990
rect 57520 29708 57572 29714
rect 57520 29650 57572 29656
rect 57612 29708 57664 29714
rect 57612 29650 57664 29656
rect 57428 29504 57480 29510
rect 57428 29446 57480 29452
rect 57336 26444 57388 26450
rect 57336 26386 57388 26392
rect 57334 26208 57390 26217
rect 57334 26143 57390 26152
rect 57348 25362 57376 26143
rect 57336 25356 57388 25362
rect 57336 25298 57388 25304
rect 57336 24608 57388 24614
rect 57336 24550 57388 24556
rect 57244 24336 57296 24342
rect 57244 24278 57296 24284
rect 57072 22066 57192 22094
rect 57164 16574 57192 22066
rect 57244 19304 57296 19310
rect 57244 19246 57296 19252
rect 57256 18630 57284 19246
rect 57244 18624 57296 18630
rect 57244 18566 57296 18572
rect 56980 16546 57192 16574
rect 56784 16448 56836 16454
rect 56784 16390 56836 16396
rect 56692 14000 56744 14006
rect 56692 13942 56744 13948
rect 56600 11756 56652 11762
rect 56600 11698 56652 11704
rect 56692 11280 56744 11286
rect 56692 11222 56744 11228
rect 56600 7880 56652 7886
rect 56600 7822 56652 7828
rect 56612 7546 56640 7822
rect 56600 7540 56652 7546
rect 56600 7482 56652 7488
rect 56704 5914 56732 11222
rect 56796 6866 56824 16390
rect 56876 14000 56928 14006
rect 56876 13942 56928 13948
rect 56888 11626 56916 13942
rect 56876 11620 56928 11626
rect 56876 11562 56928 11568
rect 56888 11218 56916 11562
rect 56876 11212 56928 11218
rect 56876 11154 56928 11160
rect 56888 10130 56916 11154
rect 56876 10124 56928 10130
rect 56876 10066 56928 10072
rect 56888 9586 56916 10066
rect 56876 9580 56928 9586
rect 56876 9522 56928 9528
rect 56888 8022 56916 9522
rect 56980 8922 57008 16546
rect 57348 14906 57376 24550
rect 57440 22094 57468 29446
rect 57532 29238 57560 29650
rect 57520 29232 57572 29238
rect 57520 29174 57572 29180
rect 57624 29050 57652 29650
rect 57532 29034 57652 29050
rect 57520 29028 57652 29034
rect 57572 29022 57652 29028
rect 57520 28970 57572 28976
rect 57532 26790 57560 28970
rect 57520 26784 57572 26790
rect 57520 26726 57572 26732
rect 57520 25900 57572 25906
rect 57520 25842 57572 25848
rect 57532 25537 57560 25842
rect 57518 25528 57574 25537
rect 57518 25463 57574 25472
rect 57716 22094 57744 31726
rect 57808 28762 57836 37318
rect 57900 37262 57928 37946
rect 57888 37256 57940 37262
rect 57888 37198 57940 37204
rect 57992 37194 58020 38218
rect 58084 38010 58112 56646
rect 58176 56302 58204 57190
rect 58348 56840 58400 56846
rect 58348 56782 58400 56788
rect 58360 56545 58388 56782
rect 58346 56536 58402 56545
rect 58346 56471 58402 56480
rect 58452 56370 58480 58103
rect 58440 56364 58492 56370
rect 58440 56306 58492 56312
rect 58164 56296 58216 56302
rect 58164 56238 58216 56244
rect 58164 56160 58216 56166
rect 58164 56102 58216 56108
rect 58176 50386 58204 56102
rect 58452 55962 58480 56306
rect 58440 55956 58492 55962
rect 58440 55898 58492 55904
rect 58348 55752 58400 55758
rect 58346 55720 58348 55729
rect 58400 55720 58402 55729
rect 58346 55655 58402 55664
rect 58532 55616 58584 55622
rect 58532 55558 58584 55564
rect 58348 55412 58400 55418
rect 58348 55354 58400 55360
rect 58360 55214 58388 55354
rect 58268 55186 58388 55214
rect 58164 50380 58216 50386
rect 58164 50322 58216 50328
rect 58164 40928 58216 40934
rect 58164 40870 58216 40876
rect 58176 40089 58204 40870
rect 58162 40080 58218 40089
rect 58162 40015 58218 40024
rect 58268 38434 58296 55186
rect 58348 54528 58400 54534
rect 58348 54470 58400 54476
rect 58360 54194 58388 54470
rect 58348 54188 58400 54194
rect 58348 54130 58400 54136
rect 58360 54097 58388 54130
rect 58346 54088 58402 54097
rect 58346 54023 58402 54032
rect 58348 53576 58400 53582
rect 58348 53518 58400 53524
rect 58360 53281 58388 53518
rect 58346 53272 58402 53281
rect 58346 53207 58402 53216
rect 58348 52488 58400 52494
rect 58346 52456 58348 52465
rect 58400 52456 58402 52465
rect 58346 52391 58402 52400
rect 58348 52012 58400 52018
rect 58348 51954 58400 51960
rect 58360 51649 58388 51954
rect 58346 51640 58402 51649
rect 58346 51575 58402 51584
rect 58348 51264 58400 51270
rect 58348 51206 58400 51212
rect 58360 50930 58388 51206
rect 58348 50924 58400 50930
rect 58348 50866 58400 50872
rect 58360 50833 58388 50866
rect 58346 50824 58402 50833
rect 58346 50759 58402 50768
rect 58348 50312 58400 50318
rect 58348 50254 58400 50260
rect 58360 50017 58388 50254
rect 58346 50008 58402 50017
rect 58346 49943 58402 49952
rect 58348 49224 58400 49230
rect 58346 49192 58348 49201
rect 58400 49192 58402 49201
rect 58346 49127 58402 49136
rect 58348 48748 58400 48754
rect 58348 48690 58400 48696
rect 58360 48385 58388 48690
rect 58346 48376 58402 48385
rect 58346 48311 58402 48320
rect 58348 48000 58400 48006
rect 58348 47942 58400 47948
rect 58360 47666 58388 47942
rect 58348 47660 58400 47666
rect 58348 47602 58400 47608
rect 58360 47569 58388 47602
rect 58346 47560 58402 47569
rect 58346 47495 58402 47504
rect 58348 47048 58400 47054
rect 58348 46990 58400 46996
rect 58360 46753 58388 46990
rect 58346 46744 58402 46753
rect 58346 46679 58402 46688
rect 58348 45960 58400 45966
rect 58346 45928 58348 45937
rect 58400 45928 58402 45937
rect 58346 45863 58402 45872
rect 58348 45484 58400 45490
rect 58348 45426 58400 45432
rect 58360 45121 58388 45426
rect 58346 45112 58402 45121
rect 58346 45047 58402 45056
rect 58348 44736 58400 44742
rect 58348 44678 58400 44684
rect 58360 44402 58388 44678
rect 58348 44396 58400 44402
rect 58348 44338 58400 44344
rect 58360 44305 58388 44338
rect 58346 44296 58402 44305
rect 58346 44231 58402 44240
rect 58348 43784 58400 43790
rect 58348 43726 58400 43732
rect 58360 43489 58388 43726
rect 58346 43480 58402 43489
rect 58346 43415 58402 43424
rect 58348 42696 58400 42702
rect 58346 42664 58348 42673
rect 58400 42664 58402 42673
rect 58346 42599 58402 42608
rect 58348 42220 58400 42226
rect 58348 42162 58400 42168
rect 58360 41857 58388 42162
rect 58346 41848 58402 41857
rect 58346 41783 58402 41792
rect 58348 41472 58400 41478
rect 58348 41414 58400 41420
rect 58360 41138 58388 41414
rect 58348 41132 58400 41138
rect 58348 41074 58400 41080
rect 58360 41041 58388 41074
rect 58346 41032 58402 41041
rect 58346 40967 58402 40976
rect 58348 40520 58400 40526
rect 58348 40462 58400 40468
rect 58360 40225 58388 40462
rect 58346 40216 58402 40225
rect 58346 40151 58402 40160
rect 58348 39908 58400 39914
rect 58348 39850 58400 39856
rect 58360 39438 58388 39850
rect 58348 39432 58400 39438
rect 58346 39400 58348 39409
rect 58400 39400 58402 39409
rect 58346 39335 58402 39344
rect 58348 38956 58400 38962
rect 58348 38898 58400 38904
rect 58360 38593 58388 38898
rect 58346 38584 58402 38593
rect 58346 38519 58402 38528
rect 58268 38406 58480 38434
rect 58256 38344 58308 38350
rect 58256 38286 58308 38292
rect 58072 38004 58124 38010
rect 58072 37946 58124 37952
rect 57980 37188 58032 37194
rect 57980 37130 58032 37136
rect 58072 37120 58124 37126
rect 58072 37062 58124 37068
rect 57980 35828 58032 35834
rect 57980 35770 58032 35776
rect 57992 35222 58020 35770
rect 57980 35216 58032 35222
rect 57980 35158 58032 35164
rect 57888 34604 57940 34610
rect 57888 34546 57940 34552
rect 57900 34513 57928 34546
rect 57886 34504 57942 34513
rect 57886 34439 57942 34448
rect 57888 33856 57940 33862
rect 57888 33798 57940 33804
rect 57900 33522 57928 33798
rect 57888 33516 57940 33522
rect 57888 33458 57940 33464
rect 57900 32881 57928 33458
rect 57980 33312 58032 33318
rect 57980 33254 58032 33260
rect 57886 32872 57942 32881
rect 57886 32807 57942 32816
rect 57992 30734 58020 33254
rect 57980 30728 58032 30734
rect 57980 30670 58032 30676
rect 57886 29608 57942 29617
rect 57886 29543 57942 29552
rect 57900 29170 57928 29543
rect 57888 29164 57940 29170
rect 57888 29106 57940 29112
rect 57796 28756 57848 28762
rect 57796 28698 57848 28704
rect 57900 28694 57928 29106
rect 57888 28688 57940 28694
rect 57888 28630 57940 28636
rect 58084 27606 58112 37062
rect 58164 36032 58216 36038
rect 58164 35974 58216 35980
rect 58176 35154 58204 35974
rect 58164 35148 58216 35154
rect 58164 35090 58216 35096
rect 58268 33658 58296 38286
rect 58348 37868 58400 37874
rect 58348 37810 58400 37816
rect 58360 37777 58388 37810
rect 58346 37768 58402 37777
rect 58346 37703 58402 37712
rect 58346 36952 58402 36961
rect 58346 36887 58402 36896
rect 58360 36786 58388 36887
rect 58348 36780 58400 36786
rect 58348 36722 58400 36728
rect 58348 36168 58400 36174
rect 58346 36136 58348 36145
rect 58400 36136 58402 36145
rect 58346 36071 58402 36080
rect 58348 35692 58400 35698
rect 58348 35634 58400 35640
rect 58360 35329 58388 35634
rect 58346 35320 58402 35329
rect 58346 35255 58402 35264
rect 58452 34542 58480 38406
rect 58544 35834 58572 55558
rect 59176 53984 59228 53990
rect 59176 53926 59228 53932
rect 58992 51808 59044 51814
rect 58992 51750 59044 51756
rect 58900 50720 58952 50726
rect 58900 50662 58952 50668
rect 58624 50380 58676 50386
rect 58624 50322 58676 50328
rect 58636 44334 58664 50322
rect 58808 49088 58860 49094
rect 58808 49030 58860 49036
rect 58716 45824 58768 45830
rect 58716 45766 58768 45772
rect 58624 44328 58676 44334
rect 58624 44270 58676 44276
rect 58624 44192 58676 44198
rect 58624 44134 58676 44140
rect 58532 35828 58584 35834
rect 58532 35770 58584 35776
rect 58440 34536 58492 34542
rect 58440 34478 58492 34484
rect 58348 34400 58400 34406
rect 58348 34342 58400 34348
rect 58256 33652 58308 33658
rect 58256 33594 58308 33600
rect 58360 32978 58388 34342
rect 58440 33992 58492 33998
rect 58440 33934 58492 33940
rect 58452 33697 58480 33934
rect 58438 33688 58494 33697
rect 58438 33623 58494 33632
rect 58636 33046 58664 44134
rect 58728 35290 58756 45766
rect 58820 38282 58848 49030
rect 58808 38276 58860 38282
rect 58808 38218 58860 38224
rect 58716 35284 58768 35290
rect 58716 35226 58768 35232
rect 58808 35080 58860 35086
rect 58808 35022 58860 35028
rect 58624 33040 58676 33046
rect 58624 32982 58676 32988
rect 58348 32972 58400 32978
rect 58348 32914 58400 32920
rect 58624 32904 58676 32910
rect 58624 32846 58676 32852
rect 58164 32428 58216 32434
rect 58164 32370 58216 32376
rect 58348 32428 58400 32434
rect 58348 32370 58400 32376
rect 58176 31958 58204 32370
rect 58256 32224 58308 32230
rect 58256 32166 58308 32172
rect 58164 31952 58216 31958
rect 58164 31894 58216 31900
rect 58164 31340 58216 31346
rect 58164 31282 58216 31288
rect 58176 31249 58204 31282
rect 58162 31240 58218 31249
rect 58162 31175 58218 31184
rect 58162 30424 58218 30433
rect 58162 30359 58218 30368
rect 58176 30258 58204 30359
rect 58164 30252 58216 30258
rect 58164 30194 58216 30200
rect 58268 29714 58296 32166
rect 58360 32065 58388 32370
rect 58346 32056 58402 32065
rect 58346 31991 58348 32000
rect 58400 31991 58402 32000
rect 58348 31962 58400 31968
rect 58440 31476 58492 31482
rect 58440 31418 58492 31424
rect 58348 31136 58400 31142
rect 58348 31078 58400 31084
rect 58256 29708 58308 29714
rect 58256 29650 58308 29656
rect 58360 28914 58388 31078
rect 58452 30666 58480 31418
rect 58440 30660 58492 30666
rect 58440 30602 58492 30608
rect 58440 30048 58492 30054
rect 58440 29990 58492 29996
rect 58268 28886 58388 28914
rect 58072 27600 58124 27606
rect 58072 27542 58124 27548
rect 57980 27532 58032 27538
rect 57980 27474 58032 27480
rect 57796 26784 57848 26790
rect 57796 26726 57848 26732
rect 57808 26450 57836 26726
rect 57992 26518 58020 27474
rect 57980 26512 58032 26518
rect 57980 26454 58032 26460
rect 57796 26444 57848 26450
rect 57796 26386 57848 26392
rect 57808 25362 57836 26386
rect 58268 25362 58296 28886
rect 58346 28792 58402 28801
rect 58346 28727 58402 28736
rect 58360 28558 58388 28727
rect 58348 28552 58400 28558
rect 58348 28494 58400 28500
rect 58360 28218 58388 28494
rect 58348 28212 58400 28218
rect 58348 28154 58400 28160
rect 58348 28076 58400 28082
rect 58348 28018 58400 28024
rect 58360 27985 58388 28018
rect 58346 27976 58402 27985
rect 58346 27911 58402 27920
rect 58360 27674 58388 27911
rect 58348 27668 58400 27674
rect 58348 27610 58400 27616
rect 58348 27464 58400 27470
rect 58348 27406 58400 27412
rect 58360 27169 58388 27406
rect 58346 27160 58402 27169
rect 58346 27095 58348 27104
rect 58400 27095 58402 27104
rect 58348 27066 58400 27072
rect 58452 26450 58480 29990
rect 58440 26444 58492 26450
rect 58440 26386 58492 26392
rect 58346 26344 58402 26353
rect 58346 26279 58402 26288
rect 58440 26308 58492 26314
rect 58360 25906 58388 26279
rect 58440 26250 58492 26256
rect 58348 25900 58400 25906
rect 58348 25842 58400 25848
rect 57796 25356 57848 25362
rect 57796 25298 57848 25304
rect 58256 25356 58308 25362
rect 58256 25298 58308 25304
rect 57808 24682 57836 25298
rect 58164 25288 58216 25294
rect 58164 25230 58216 25236
rect 57980 25152 58032 25158
rect 57980 25094 58032 25100
rect 57796 24676 57848 24682
rect 57796 24618 57848 24624
rect 57992 23186 58020 25094
rect 57980 23180 58032 23186
rect 57980 23122 58032 23128
rect 57440 22066 57560 22094
rect 57716 22066 57928 22094
rect 57532 19310 57560 22066
rect 57520 19304 57572 19310
rect 57520 19246 57572 19252
rect 57428 18080 57480 18086
rect 57428 18022 57480 18028
rect 57164 14878 57376 14906
rect 57164 13394 57192 14878
rect 57336 14816 57388 14822
rect 57336 14758 57388 14764
rect 57348 13394 57376 14758
rect 57152 13388 57204 13394
rect 57152 13330 57204 13336
rect 57336 13388 57388 13394
rect 57336 13330 57388 13336
rect 57164 12986 57192 13330
rect 57152 12980 57204 12986
rect 57152 12922 57204 12928
rect 57164 11898 57192 12922
rect 57152 11892 57204 11898
rect 57152 11834 57204 11840
rect 57164 11354 57192 11834
rect 57152 11348 57204 11354
rect 57152 11290 57204 11296
rect 57164 10146 57192 11290
rect 57072 10118 57192 10146
rect 57072 9994 57100 10118
rect 57060 9988 57112 9994
rect 57060 9930 57112 9936
rect 57072 9654 57100 9930
rect 57440 9926 57468 18022
rect 57796 15904 57848 15910
rect 57796 15846 57848 15852
rect 57704 14000 57756 14006
rect 57704 13942 57756 13948
rect 57716 13394 57744 13942
rect 57704 13388 57756 13394
rect 57704 13330 57756 13336
rect 57704 12844 57756 12850
rect 57704 12786 57756 12792
rect 57716 12442 57744 12786
rect 57704 12436 57756 12442
rect 57704 12378 57756 12384
rect 57612 12096 57664 12102
rect 57612 12038 57664 12044
rect 57518 10840 57574 10849
rect 57518 10775 57520 10784
rect 57572 10775 57574 10784
rect 57520 10746 57572 10752
rect 57336 9920 57388 9926
rect 57336 9862 57388 9868
rect 57428 9920 57480 9926
rect 57428 9862 57480 9868
rect 57060 9648 57112 9654
rect 57060 9590 57112 9596
rect 57072 9110 57100 9590
rect 57060 9104 57112 9110
rect 57060 9046 57112 9052
rect 56980 8894 57284 8922
rect 56876 8016 56928 8022
rect 56876 7958 56928 7964
rect 57152 8016 57204 8022
rect 57152 7958 57204 7964
rect 56876 7880 56928 7886
rect 56876 7822 56928 7828
rect 56784 6860 56836 6866
rect 56784 6802 56836 6808
rect 56784 6180 56836 6186
rect 56784 6122 56836 6128
rect 56692 5908 56744 5914
rect 56692 5850 56744 5856
rect 56796 5846 56824 6122
rect 56784 5840 56836 5846
rect 56784 5782 56836 5788
rect 56692 5704 56744 5710
rect 56692 5646 56744 5652
rect 56508 4820 56560 4826
rect 56508 4762 56560 4768
rect 56520 4162 56548 4762
rect 56520 4134 56640 4162
rect 56140 4072 56192 4078
rect 56140 4014 56192 4020
rect 56508 3936 56560 3942
rect 56508 3878 56560 3884
rect 56140 3392 56192 3398
rect 56140 3334 56192 3340
rect 55600 3182 56088 3210
rect 55600 2446 55628 3182
rect 55956 3052 56008 3058
rect 55956 2994 56008 3000
rect 56048 3052 56100 3058
rect 56048 2994 56100 3000
rect 55680 2644 55732 2650
rect 55680 2586 55732 2592
rect 55496 2440 55548 2446
rect 55496 2382 55548 2388
rect 55588 2440 55640 2446
rect 55588 2382 55640 2388
rect 55692 2378 55720 2586
rect 55968 2446 55996 2994
rect 56060 2854 56088 2994
rect 56152 2990 56180 3334
rect 56520 3058 56548 3878
rect 56612 3534 56640 4134
rect 56600 3528 56652 3534
rect 56600 3470 56652 3476
rect 56704 3194 56732 5646
rect 56784 3392 56836 3398
rect 56784 3334 56836 3340
rect 56692 3188 56744 3194
rect 56692 3130 56744 3136
rect 56508 3052 56560 3058
rect 56508 2994 56560 3000
rect 56140 2984 56192 2990
rect 56140 2926 56192 2932
rect 56048 2848 56100 2854
rect 56048 2790 56100 2796
rect 55956 2440 56008 2446
rect 55956 2382 56008 2388
rect 55680 2372 55732 2378
rect 55680 2314 55732 2320
rect 55404 2100 55456 2106
rect 55404 2042 55456 2048
rect 56060 1873 56088 2790
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 56046 1864 56102 1873
rect 56046 1799 56102 1808
rect 56428 800 56456 2382
rect 56520 1057 56548 2994
rect 56796 2514 56824 3334
rect 56784 2508 56836 2514
rect 56784 2450 56836 2456
rect 56888 2310 56916 7822
rect 56968 7472 57020 7478
rect 56968 7414 57020 7420
rect 56980 7002 57008 7414
rect 57164 7342 57192 7958
rect 57152 7336 57204 7342
rect 57152 7278 57204 7284
rect 56968 6996 57020 7002
rect 56968 6938 57020 6944
rect 56980 6458 57008 6938
rect 57164 6934 57192 7278
rect 57152 6928 57204 6934
rect 57152 6870 57204 6876
rect 57152 6792 57204 6798
rect 57152 6734 57204 6740
rect 56968 6452 57020 6458
rect 56968 6394 57020 6400
rect 56980 5574 57008 6394
rect 57060 6112 57112 6118
rect 57060 6054 57112 6060
rect 57072 5778 57100 6054
rect 57060 5772 57112 5778
rect 57060 5714 57112 5720
rect 56968 5568 57020 5574
rect 56968 5510 57020 5516
rect 56980 5370 57008 5510
rect 56968 5364 57020 5370
rect 56968 5306 57020 5312
rect 57164 2854 57192 6734
rect 57256 5930 57284 8894
rect 57348 8378 57376 9862
rect 57348 8350 57560 8378
rect 57428 8288 57480 8294
rect 57428 8230 57480 8236
rect 57336 6928 57388 6934
rect 57336 6870 57388 6876
rect 57348 6458 57376 6870
rect 57336 6452 57388 6458
rect 57336 6394 57388 6400
rect 57348 6186 57376 6394
rect 57336 6180 57388 6186
rect 57336 6122 57388 6128
rect 57256 5902 57376 5930
rect 57244 5840 57296 5846
rect 57244 5782 57296 5788
rect 57256 5370 57284 5782
rect 57244 5364 57296 5370
rect 57244 5306 57296 5312
rect 57348 3670 57376 5902
rect 57440 5778 57468 8230
rect 57428 5772 57480 5778
rect 57428 5714 57480 5720
rect 57532 4826 57560 8350
rect 57624 7954 57652 12038
rect 57808 10146 57836 15846
rect 57716 10118 57836 10146
rect 57716 8294 57744 10118
rect 57794 10024 57850 10033
rect 57794 9959 57850 9968
rect 57808 9586 57836 9959
rect 57796 9580 57848 9586
rect 57796 9522 57848 9528
rect 57808 9178 57836 9522
rect 57796 9172 57848 9178
rect 57796 9114 57848 9120
rect 57796 9036 57848 9042
rect 57796 8978 57848 8984
rect 57704 8288 57756 8294
rect 57704 8230 57756 8236
rect 57808 8106 57836 8978
rect 57716 8078 57836 8106
rect 57716 7954 57744 8078
rect 57612 7948 57664 7954
rect 57612 7890 57664 7896
rect 57704 7948 57756 7954
rect 57704 7890 57756 7896
rect 57716 7478 57744 7890
rect 57704 7472 57756 7478
rect 57704 7414 57756 7420
rect 57900 6914 57928 22066
rect 58176 21690 58204 25230
rect 58348 24812 58400 24818
rect 58348 24754 58400 24760
rect 58360 24721 58388 24754
rect 58346 24712 58402 24721
rect 58346 24647 58402 24656
rect 58360 24410 58388 24647
rect 58348 24404 58400 24410
rect 58348 24346 58400 24352
rect 58452 24290 58480 26250
rect 58636 24682 58664 32846
rect 58716 29640 58768 29646
rect 58716 29582 58768 29588
rect 58624 24676 58676 24682
rect 58624 24618 58676 24624
rect 58268 24262 58480 24290
rect 58164 21684 58216 21690
rect 58164 21626 58216 21632
rect 58268 21146 58296 24262
rect 58348 24200 58400 24206
rect 58348 24142 58400 24148
rect 58360 23905 58388 24142
rect 58346 23896 58402 23905
rect 58346 23831 58402 23840
rect 58346 23080 58402 23089
rect 58346 23015 58402 23024
rect 58360 22642 58388 23015
rect 58348 22636 58400 22642
rect 58348 22578 58400 22584
rect 58346 22264 58402 22273
rect 58346 22199 58402 22208
rect 58360 22030 58388 22199
rect 58348 22024 58400 22030
rect 58348 21966 58400 21972
rect 58728 21894 58756 29582
rect 58820 26042 58848 35022
rect 58808 26036 58860 26042
rect 58808 25978 58860 25984
rect 58912 25430 58940 50662
rect 59004 36582 59032 51750
rect 59084 50176 59136 50182
rect 59084 50118 59136 50124
rect 58992 36576 59044 36582
rect 58992 36518 59044 36524
rect 59096 35154 59124 50118
rect 59188 38350 59216 53926
rect 59636 53440 59688 53446
rect 59636 53382 59688 53388
rect 59268 52624 59320 52630
rect 59268 52566 59320 52572
rect 59176 38344 59228 38350
rect 59176 38286 59228 38292
rect 59176 38208 59228 38214
rect 59176 38150 59228 38156
rect 59084 35148 59136 35154
rect 59084 35090 59136 35096
rect 59188 35034 59216 38150
rect 59004 35006 59216 35034
rect 59004 29306 59032 35006
rect 59084 34944 59136 34950
rect 59084 34886 59136 34892
rect 58992 29300 59044 29306
rect 58992 29242 59044 29248
rect 59096 27538 59124 34886
rect 59280 31482 59308 52566
rect 59544 47184 59596 47190
rect 59544 47126 59596 47132
rect 59452 42016 59504 42022
rect 59452 41958 59504 41964
rect 59360 36576 59412 36582
rect 59360 36518 59412 36524
rect 59268 31476 59320 31482
rect 59268 31418 59320 31424
rect 59372 29238 59400 36518
rect 59360 29232 59412 29238
rect 59360 29174 59412 29180
rect 59464 29102 59492 41958
rect 59556 37194 59584 47126
rect 59544 37188 59596 37194
rect 59544 37130 59596 37136
rect 59648 31958 59676 53382
rect 59820 48544 59872 48550
rect 59820 48486 59872 48492
rect 59728 43648 59780 43654
rect 59728 43590 59780 43596
rect 59740 32570 59768 43590
rect 59832 39370 59860 48486
rect 59820 39364 59872 39370
rect 59820 39306 59872 39312
rect 59820 37664 59872 37670
rect 59820 37606 59872 37612
rect 59728 32564 59780 32570
rect 59728 32506 59780 32512
rect 59636 31952 59688 31958
rect 59636 31894 59688 31900
rect 59452 29096 59504 29102
rect 59452 29038 59504 29044
rect 59832 27946 59860 37606
rect 59820 27940 59872 27946
rect 59820 27882 59872 27888
rect 59084 27532 59136 27538
rect 59084 27474 59136 27480
rect 58900 25424 58952 25430
rect 58900 25366 58952 25372
rect 58912 23866 58940 25366
rect 58900 23860 58952 23866
rect 58900 23802 58952 23808
rect 58716 21888 58768 21894
rect 58716 21830 58768 21836
rect 58348 21548 58400 21554
rect 58348 21490 58400 21496
rect 58360 21457 58388 21490
rect 58346 21448 58402 21457
rect 58346 21383 58402 21392
rect 58256 21140 58308 21146
rect 58256 21082 58308 21088
rect 58348 20936 58400 20942
rect 58348 20878 58400 20884
rect 58360 20641 58388 20878
rect 58346 20632 58402 20641
rect 58346 20567 58402 20576
rect 58348 19848 58400 19854
rect 58346 19816 58348 19825
rect 58400 19816 58402 19825
rect 58346 19751 58402 19760
rect 58072 19712 58124 19718
rect 58072 19654 58124 19660
rect 57980 14272 58032 14278
rect 57980 14214 58032 14220
rect 57992 11762 58020 14214
rect 58084 13462 58112 19654
rect 58348 19372 58400 19378
rect 58348 19314 58400 19320
rect 58360 19009 58388 19314
rect 58346 19000 58402 19009
rect 58346 18935 58348 18944
rect 58400 18935 58402 18944
rect 58348 18906 58400 18912
rect 58348 18284 58400 18290
rect 58348 18226 58400 18232
rect 58360 18193 58388 18226
rect 58346 18184 58402 18193
rect 58346 18119 58402 18128
rect 58348 17672 58400 17678
rect 58348 17614 58400 17620
rect 58360 17377 58388 17614
rect 58716 17536 58768 17542
rect 58716 17478 58768 17484
rect 58346 17368 58402 17377
rect 58346 17303 58402 17312
rect 58348 16584 58400 16590
rect 58346 16552 58348 16561
rect 58400 16552 58402 16561
rect 58346 16487 58402 16496
rect 58348 16108 58400 16114
rect 58348 16050 58400 16056
rect 58360 15745 58388 16050
rect 58346 15736 58402 15745
rect 58346 15671 58348 15680
rect 58400 15671 58402 15680
rect 58348 15642 58400 15648
rect 58348 15020 58400 15026
rect 58348 14962 58400 14968
rect 58360 14929 58388 14962
rect 58346 14920 58402 14929
rect 58346 14855 58402 14864
rect 58348 14408 58400 14414
rect 58348 14350 58400 14356
rect 58360 14113 58388 14350
rect 58346 14104 58402 14113
rect 58346 14039 58402 14048
rect 58072 13456 58124 13462
rect 58072 13398 58124 13404
rect 58532 13388 58584 13394
rect 58532 13330 58584 13336
rect 58256 13320 58308 13326
rect 58256 13262 58308 13268
rect 58346 13288 58402 13297
rect 58164 12640 58216 12646
rect 58164 12582 58216 12588
rect 57980 11756 58032 11762
rect 57980 11698 58032 11704
rect 58072 11688 58124 11694
rect 58072 11630 58124 11636
rect 57980 11620 58032 11626
rect 57980 11562 58032 11568
rect 57992 10198 58020 11562
rect 57980 10192 58032 10198
rect 57980 10134 58032 10140
rect 57980 10056 58032 10062
rect 57980 9998 58032 10004
rect 57992 8362 58020 9998
rect 58084 9178 58112 11630
rect 58176 9994 58204 12582
rect 58164 9988 58216 9994
rect 58164 9930 58216 9936
rect 58268 9450 58296 13262
rect 58346 13223 58402 13232
rect 58360 12850 58388 13223
rect 58348 12844 58400 12850
rect 58348 12786 58400 12792
rect 58346 12472 58402 12481
rect 58346 12407 58402 12416
rect 58360 12238 58388 12407
rect 58348 12232 58400 12238
rect 58348 12174 58400 12180
rect 58348 11756 58400 11762
rect 58348 11698 58400 11704
rect 58360 11665 58388 11698
rect 58346 11656 58402 11665
rect 58346 11591 58402 11600
rect 58360 10810 58388 11591
rect 58440 11144 58492 11150
rect 58440 11086 58492 11092
rect 58452 10849 58480 11086
rect 58438 10840 58494 10849
rect 58348 10804 58400 10810
rect 58438 10775 58494 10784
rect 58348 10746 58400 10752
rect 58348 10192 58400 10198
rect 58348 10134 58400 10140
rect 58256 9444 58308 9450
rect 58256 9386 58308 9392
rect 58360 9330 58388 10134
rect 58176 9302 58388 9330
rect 58072 9172 58124 9178
rect 58072 9114 58124 9120
rect 57980 8356 58032 8362
rect 57980 8298 58032 8304
rect 57808 6886 57928 6914
rect 57612 5908 57664 5914
rect 57612 5850 57664 5856
rect 57624 5778 57652 5850
rect 57612 5772 57664 5778
rect 57612 5714 57664 5720
rect 57704 5704 57756 5710
rect 57704 5646 57756 5652
rect 57716 5574 57744 5646
rect 57704 5568 57756 5574
rect 57704 5510 57756 5516
rect 57520 4820 57572 4826
rect 57520 4762 57572 4768
rect 57704 4616 57756 4622
rect 57704 4558 57756 4564
rect 57336 3664 57388 3670
rect 57336 3606 57388 3612
rect 57348 3058 57376 3606
rect 57428 3528 57480 3534
rect 57716 3505 57744 4558
rect 57808 4146 57836 6886
rect 58176 4826 58204 9302
rect 58346 9208 58402 9217
rect 58346 9143 58402 9152
rect 58360 8974 58388 9143
rect 58348 8968 58400 8974
rect 58348 8910 58400 8916
rect 58360 8634 58388 8910
rect 58348 8628 58400 8634
rect 58348 8570 58400 8576
rect 58348 8492 58400 8498
rect 58348 8434 58400 8440
rect 58360 8401 58388 8434
rect 58346 8392 58402 8401
rect 58346 8327 58402 8336
rect 58440 7744 58492 7750
rect 58440 7686 58492 7692
rect 58346 7576 58402 7585
rect 58346 7511 58402 7520
rect 58360 7410 58388 7511
rect 58348 7404 58400 7410
rect 58348 7346 58400 7352
rect 58348 6792 58400 6798
rect 58346 6760 58348 6769
rect 58400 6760 58402 6769
rect 58346 6695 58402 6704
rect 58360 6458 58388 6695
rect 58348 6452 58400 6458
rect 58348 6394 58400 6400
rect 58348 6316 58400 6322
rect 58348 6258 58400 6264
rect 58360 5953 58388 6258
rect 58346 5944 58402 5953
rect 58346 5879 58402 5888
rect 58256 5568 58308 5574
rect 58256 5510 58308 5516
rect 58164 4820 58216 4826
rect 58164 4762 58216 4768
rect 57796 4140 57848 4146
rect 57796 4082 57848 4088
rect 58164 3936 58216 3942
rect 58164 3878 58216 3884
rect 57428 3470 57480 3476
rect 57702 3496 57758 3505
rect 57336 3052 57388 3058
rect 57336 2994 57388 3000
rect 57152 2848 57204 2854
rect 57152 2790 57204 2796
rect 57336 2848 57388 2854
rect 57336 2790 57388 2796
rect 57348 2582 57376 2790
rect 57440 2650 57468 3470
rect 57702 3431 57758 3440
rect 57980 3392 58032 3398
rect 57980 3334 58032 3340
rect 58072 3392 58124 3398
rect 58072 3334 58124 3340
rect 57518 2680 57574 2689
rect 57428 2644 57480 2650
rect 57518 2615 57574 2624
rect 57428 2586 57480 2592
rect 57336 2576 57388 2582
rect 57336 2518 57388 2524
rect 57532 2446 57560 2615
rect 57992 2446 58020 3334
rect 58084 3126 58112 3334
rect 58072 3120 58124 3126
rect 58072 3062 58124 3068
rect 57520 2440 57572 2446
rect 57520 2382 57572 2388
rect 57980 2440 58032 2446
rect 57980 2382 58032 2388
rect 58176 2378 58204 3878
rect 58268 3534 58296 5510
rect 58348 5228 58400 5234
rect 58348 5170 58400 5176
rect 58360 5137 58388 5170
rect 58346 5128 58402 5137
rect 58346 5063 58402 5072
rect 58348 4616 58400 4622
rect 58348 4558 58400 4564
rect 58360 4321 58388 4558
rect 58346 4312 58402 4321
rect 58346 4247 58402 4256
rect 58256 3528 58308 3534
rect 58256 3470 58308 3476
rect 58452 3058 58480 7686
rect 58544 5370 58572 13330
rect 58728 8090 58756 17478
rect 58716 8084 58768 8090
rect 58716 8026 58768 8032
rect 58532 5364 58584 5370
rect 58532 5306 58584 5312
rect 58440 3052 58492 3058
rect 58440 2994 58492 3000
rect 58164 2372 58216 2378
rect 58164 2314 58216 2320
rect 56876 2304 56928 2310
rect 56876 2246 56928 2252
rect 57520 2304 57572 2310
rect 57520 2246 57572 2252
rect 56506 1048 56562 1057
rect 56506 983 56562 992
rect 57532 800 57560 2246
rect 35544 734 35848 762
rect 36542 0 36598 800
rect 37646 0 37702 800
rect 38750 0 38806 800
rect 39854 0 39910 800
rect 40958 0 41014 800
rect 42062 0 42118 800
rect 43166 0 43222 800
rect 44270 0 44326 800
rect 45374 0 45430 800
rect 46478 0 46534 800
rect 47582 0 47638 800
rect 48686 0 48742 800
rect 49790 0 49846 800
rect 50894 0 50950 800
rect 51998 0 52054 800
rect 53102 0 53158 800
rect 54206 0 54262 800
rect 55310 0 55366 800
rect 56414 0 56470 800
rect 57518 0 57574 800
<< via2 >>
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 1674 55664 1730 55720
rect 1674 54848 1730 54904
rect 1674 54052 1730 54088
rect 1674 54032 1676 54052
rect 1676 54032 1728 54052
rect 1728 54032 1730 54052
rect 1674 53216 1730 53272
rect 1674 52400 1730 52456
rect 1674 51584 1730 51640
rect 1674 50788 1730 50824
rect 1674 50768 1676 50788
rect 1676 50768 1728 50788
rect 1728 50768 1730 50788
rect 1674 49952 1730 50008
rect 1674 49136 1730 49192
rect 1674 48320 1730 48376
rect 1674 47524 1730 47560
rect 1674 47504 1676 47524
rect 1676 47504 1728 47524
rect 1728 47504 1730 47524
rect 1674 46688 1730 46744
rect 1674 45872 1730 45928
rect 1674 45056 1730 45112
rect 1674 44260 1730 44296
rect 1674 44240 1676 44260
rect 1676 44240 1728 44260
rect 1728 44240 1730 44260
rect 1674 43424 1730 43480
rect 1674 42608 1730 42664
rect 1674 41792 1730 41848
rect 1674 40996 1730 41032
rect 1674 40976 1676 40996
rect 1676 40976 1728 40996
rect 1728 40976 1730 40996
rect 1674 40160 1730 40216
rect 1674 39344 1730 39400
rect 1674 38528 1730 38584
rect 1674 37732 1730 37768
rect 1674 37712 1676 37732
rect 1676 37712 1728 37732
rect 1728 37712 1730 37732
rect 1674 36896 1730 36952
rect 1674 36080 1730 36136
rect 1674 35264 1730 35320
rect 1674 34468 1730 34504
rect 1674 34448 1676 34468
rect 1676 34448 1728 34468
rect 1728 34448 1730 34468
rect 1674 33632 1730 33688
rect 1674 32816 1730 32872
rect 1674 32000 1730 32056
rect 1674 31204 1730 31240
rect 1674 31184 1676 31204
rect 1676 31184 1728 31204
rect 1728 31184 1730 31204
rect 1674 30368 1730 30424
rect 1674 29552 1730 29608
rect 1674 28736 1730 28792
rect 1674 27940 1730 27976
rect 1674 27920 1676 27940
rect 1676 27920 1728 27940
rect 1728 27920 1730 27940
rect 1674 27104 1730 27160
rect 1674 26288 1730 26344
rect 1674 25492 1730 25528
rect 1674 25472 1676 25492
rect 1676 25472 1728 25492
rect 1728 25472 1730 25492
rect 1674 24676 1730 24712
rect 1674 24656 1676 24676
rect 1676 24656 1728 24676
rect 1728 24656 1730 24676
rect 1674 23840 1730 23896
rect 1674 23024 1730 23080
rect 1674 22228 1730 22264
rect 1674 22208 1676 22228
rect 1676 22208 1728 22228
rect 1728 22208 1730 22228
rect 1674 21412 1730 21448
rect 1674 21392 1676 21412
rect 1676 21392 1728 21412
rect 1728 21392 1730 21412
rect 1674 20596 1730 20632
rect 1674 20576 1676 20596
rect 1676 20576 1728 20596
rect 1728 20576 1730 20596
rect 1674 19760 1730 19816
rect 1674 18944 1730 19000
rect 1674 18128 1730 18184
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 1674 17332 1730 17368
rect 1674 17312 1676 17332
rect 1676 17312 1728 17332
rect 1728 17312 1730 17332
rect 1674 16496 1730 16552
rect 1674 15680 1730 15736
rect 1674 14884 1730 14920
rect 1674 14864 1676 14884
rect 1676 14864 1728 14884
rect 1728 14864 1730 14884
rect 1674 14068 1730 14104
rect 1674 14048 1676 14068
rect 1676 14048 1728 14068
rect 1728 14048 1730 14068
rect 1674 13232 1730 13288
rect 1674 12416 1730 12472
rect 1674 11600 1730 11656
rect 1674 10804 1730 10840
rect 1674 10784 1676 10804
rect 1676 10784 1728 10804
rect 1728 10784 1730 10804
rect 1674 9968 1730 10024
rect 1674 9152 1730 9208
rect 1674 8336 1730 8392
rect 1674 6704 1730 6760
rect 1674 5908 1730 5944
rect 1674 5888 1676 5908
rect 1676 5888 1728 5908
rect 1728 5888 1730 5908
rect 1674 5092 1730 5128
rect 1674 5072 1676 5092
rect 1676 5072 1728 5092
rect 1728 5072 1730 5092
rect 1674 4256 1730 4312
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 2410 7520 2466 7576
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 23478 55800 23534 55856
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 24950 55800 25006 55856
rect 24950 54168 25006 54224
rect 26054 55800 26110 55856
rect 27342 54188 27398 54224
rect 27342 54168 27344 54188
rect 27344 54168 27396 54188
rect 27396 54168 27398 54188
rect 29826 56380 29828 56400
rect 29828 56380 29880 56400
rect 29880 56380 29882 56400
rect 29826 56344 29882 56380
rect 30194 56480 30250 56536
rect 33414 56228 33470 56264
rect 33414 56208 33416 56228
rect 33416 56208 33468 56228
rect 33468 56208 33470 56228
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 35162 56344 35218 56400
rect 35806 56364 35862 56400
rect 35806 56344 35808 56364
rect 35808 56344 35860 56364
rect 35860 56344 35862 56364
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 36266 56480 36322 56536
rect 36910 56364 36966 56400
rect 36910 56344 36912 56364
rect 36912 56344 36964 56364
rect 36964 56344 36966 56364
rect 38382 56208 38438 56264
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 57518 58928 57574 58984
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 57058 57296 57114 57352
rect 58438 58112 58494 58168
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 55310 2624 55366 2680
rect 57978 54848 58034 54904
rect 57334 26152 57390 26208
rect 57518 25472 57574 25528
rect 58346 56480 58402 56536
rect 58346 55700 58348 55720
rect 58348 55700 58400 55720
rect 58400 55700 58402 55720
rect 58346 55664 58402 55700
rect 58162 40024 58218 40080
rect 58346 54032 58402 54088
rect 58346 53216 58402 53272
rect 58346 52436 58348 52456
rect 58348 52436 58400 52456
rect 58400 52436 58402 52456
rect 58346 52400 58402 52436
rect 58346 51584 58402 51640
rect 58346 50768 58402 50824
rect 58346 49952 58402 50008
rect 58346 49172 58348 49192
rect 58348 49172 58400 49192
rect 58400 49172 58402 49192
rect 58346 49136 58402 49172
rect 58346 48320 58402 48376
rect 58346 47504 58402 47560
rect 58346 46688 58402 46744
rect 58346 45908 58348 45928
rect 58348 45908 58400 45928
rect 58400 45908 58402 45928
rect 58346 45872 58402 45908
rect 58346 45056 58402 45112
rect 58346 44240 58402 44296
rect 58346 43424 58402 43480
rect 58346 42644 58348 42664
rect 58348 42644 58400 42664
rect 58400 42644 58402 42664
rect 58346 42608 58402 42644
rect 58346 41792 58402 41848
rect 58346 40976 58402 41032
rect 58346 40160 58402 40216
rect 58346 39380 58348 39400
rect 58348 39380 58400 39400
rect 58400 39380 58402 39400
rect 58346 39344 58402 39380
rect 58346 38528 58402 38584
rect 57886 34448 57942 34504
rect 57886 32816 57942 32872
rect 57886 29552 57942 29608
rect 58346 37712 58402 37768
rect 58346 36896 58402 36952
rect 58346 36116 58348 36136
rect 58348 36116 58400 36136
rect 58400 36116 58402 36136
rect 58346 36080 58402 36116
rect 58346 35264 58402 35320
rect 58438 33632 58494 33688
rect 58162 31184 58218 31240
rect 58162 30368 58218 30424
rect 58346 32020 58402 32056
rect 58346 32000 58348 32020
rect 58348 32000 58400 32020
rect 58400 32000 58402 32020
rect 58346 28736 58402 28792
rect 58346 27920 58402 27976
rect 58346 27124 58402 27160
rect 58346 27104 58348 27124
rect 58348 27104 58400 27124
rect 58400 27104 58402 27124
rect 58346 26288 58402 26344
rect 57518 10804 57574 10840
rect 57518 10784 57520 10804
rect 57520 10784 57572 10804
rect 57572 10784 57574 10804
rect 56046 1808 56102 1864
rect 57794 9968 57850 10024
rect 58346 24656 58402 24712
rect 58346 23840 58402 23896
rect 58346 23024 58402 23080
rect 58346 22208 58402 22264
rect 58346 21392 58402 21448
rect 58346 20576 58402 20632
rect 58346 19796 58348 19816
rect 58348 19796 58400 19816
rect 58400 19796 58402 19816
rect 58346 19760 58402 19796
rect 58346 18964 58402 19000
rect 58346 18944 58348 18964
rect 58348 18944 58400 18964
rect 58400 18944 58402 18964
rect 58346 18128 58402 18184
rect 58346 17312 58402 17368
rect 58346 16532 58348 16552
rect 58348 16532 58400 16552
rect 58400 16532 58402 16552
rect 58346 16496 58402 16532
rect 58346 15700 58402 15736
rect 58346 15680 58348 15700
rect 58348 15680 58400 15700
rect 58400 15680 58402 15700
rect 58346 14864 58402 14920
rect 58346 14048 58402 14104
rect 58346 13232 58402 13288
rect 58346 12416 58402 12472
rect 58346 11600 58402 11656
rect 58438 10784 58494 10840
rect 58346 9152 58402 9208
rect 58346 8336 58402 8392
rect 58346 7520 58402 7576
rect 58346 6740 58348 6760
rect 58348 6740 58400 6760
rect 58400 6740 58402 6760
rect 58346 6704 58402 6740
rect 58346 5888 58402 5944
rect 57702 3440 57758 3496
rect 57518 2624 57574 2680
rect 58346 5072 58402 5128
rect 58346 4256 58402 4312
rect 56506 992 56562 1048
<< metal3 >>
rect 57513 58986 57579 58989
rect 59200 58986 60000 59016
rect 57513 58984 60000 58986
rect 57513 58928 57518 58984
rect 57574 58928 60000 58984
rect 57513 58926 60000 58928
rect 57513 58923 57579 58926
rect 59200 58896 60000 58926
rect 58433 58170 58499 58173
rect 59200 58170 60000 58200
rect 58433 58168 60000 58170
rect 58433 58112 58438 58168
rect 58494 58112 60000 58168
rect 58433 58110 60000 58112
rect 58433 58107 58499 58110
rect 59200 58080 60000 58110
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 57053 57354 57119 57357
rect 59200 57354 60000 57384
rect 57053 57352 60000 57354
rect 57053 57296 57058 57352
rect 57114 57296 60000 57352
rect 57053 57294 60000 57296
rect 57053 57291 57119 57294
rect 59200 57264 60000 57294
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 30189 56538 30255 56541
rect 36261 56538 36327 56541
rect 30189 56536 36327 56538
rect 30189 56480 30194 56536
rect 30250 56480 36266 56536
rect 36322 56480 36327 56536
rect 30189 56478 36327 56480
rect 30189 56475 30255 56478
rect 36261 56475 36327 56478
rect 58341 56538 58407 56541
rect 59200 56538 60000 56568
rect 58341 56536 60000 56538
rect 58341 56480 58346 56536
rect 58402 56480 60000 56536
rect 58341 56478 60000 56480
rect 58341 56475 58407 56478
rect 59200 56448 60000 56478
rect 29821 56402 29887 56405
rect 35157 56402 35223 56405
rect 29821 56400 35223 56402
rect 29821 56344 29826 56400
rect 29882 56344 35162 56400
rect 35218 56344 35223 56400
rect 29821 56342 35223 56344
rect 29821 56339 29887 56342
rect 35157 56339 35223 56342
rect 35801 56402 35867 56405
rect 36905 56402 36971 56405
rect 35801 56400 36971 56402
rect 35801 56344 35806 56400
rect 35862 56344 36910 56400
rect 36966 56344 36971 56400
rect 35801 56342 36971 56344
rect 35801 56339 35867 56342
rect 36905 56339 36971 56342
rect 33409 56266 33475 56269
rect 38377 56266 38443 56269
rect 33409 56264 38443 56266
rect 33409 56208 33414 56264
rect 33470 56208 38382 56264
rect 38438 56208 38443 56264
rect 33409 56206 38443 56208
rect 33409 56203 33475 56206
rect 38377 56203 38443 56206
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 23473 55858 23539 55861
rect 24945 55858 25011 55861
rect 26049 55858 26115 55861
rect 23473 55856 26115 55858
rect 23473 55800 23478 55856
rect 23534 55800 24950 55856
rect 25006 55800 26054 55856
rect 26110 55800 26115 55856
rect 23473 55798 26115 55800
rect 23473 55795 23539 55798
rect 24945 55795 25011 55798
rect 26049 55795 26115 55798
rect 0 55722 800 55752
rect 1669 55722 1735 55725
rect 0 55720 1735 55722
rect 0 55664 1674 55720
rect 1730 55664 1735 55720
rect 0 55662 1735 55664
rect 0 55632 800 55662
rect 1669 55659 1735 55662
rect 58341 55722 58407 55725
rect 59200 55722 60000 55752
rect 58341 55720 60000 55722
rect 58341 55664 58346 55720
rect 58402 55664 60000 55720
rect 58341 55662 60000 55664
rect 58341 55659 58407 55662
rect 59200 55632 60000 55662
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 0 54906 800 54936
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 1669 54906 1735 54909
rect 0 54904 1735 54906
rect 0 54848 1674 54904
rect 1730 54848 1735 54904
rect 0 54846 1735 54848
rect 0 54816 800 54846
rect 1669 54843 1735 54846
rect 57973 54906 58039 54909
rect 59200 54906 60000 54936
rect 57973 54904 60000 54906
rect 57973 54848 57978 54904
rect 58034 54848 60000 54904
rect 57973 54846 60000 54848
rect 57973 54843 58039 54846
rect 59200 54816 60000 54846
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 24945 54226 25011 54229
rect 27337 54226 27403 54229
rect 24945 54224 27403 54226
rect 24945 54168 24950 54224
rect 25006 54168 27342 54224
rect 27398 54168 27403 54224
rect 24945 54166 27403 54168
rect 24945 54163 25011 54166
rect 27337 54163 27403 54166
rect 0 54090 800 54120
rect 1669 54090 1735 54093
rect 0 54088 1735 54090
rect 0 54032 1674 54088
rect 1730 54032 1735 54088
rect 0 54030 1735 54032
rect 0 54000 800 54030
rect 1669 54027 1735 54030
rect 58341 54090 58407 54093
rect 59200 54090 60000 54120
rect 58341 54088 60000 54090
rect 58341 54032 58346 54088
rect 58402 54032 60000 54088
rect 58341 54030 60000 54032
rect 58341 54027 58407 54030
rect 59200 54000 60000 54030
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 0 53274 800 53304
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 1669 53274 1735 53277
rect 0 53272 1735 53274
rect 0 53216 1674 53272
rect 1730 53216 1735 53272
rect 0 53214 1735 53216
rect 0 53184 800 53214
rect 1669 53211 1735 53214
rect 58341 53274 58407 53277
rect 59200 53274 60000 53304
rect 58341 53272 60000 53274
rect 58341 53216 58346 53272
rect 58402 53216 60000 53272
rect 58341 53214 60000 53216
rect 58341 53211 58407 53214
rect 59200 53184 60000 53214
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 0 52458 800 52488
rect 1669 52458 1735 52461
rect 0 52456 1735 52458
rect 0 52400 1674 52456
rect 1730 52400 1735 52456
rect 0 52398 1735 52400
rect 0 52368 800 52398
rect 1669 52395 1735 52398
rect 58341 52458 58407 52461
rect 59200 52458 60000 52488
rect 58341 52456 60000 52458
rect 58341 52400 58346 52456
rect 58402 52400 60000 52456
rect 58341 52398 60000 52400
rect 58341 52395 58407 52398
rect 59200 52368 60000 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51642 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 1669 51642 1735 51645
rect 0 51640 1735 51642
rect 0 51584 1674 51640
rect 1730 51584 1735 51640
rect 0 51582 1735 51584
rect 0 51552 800 51582
rect 1669 51579 1735 51582
rect 58341 51642 58407 51645
rect 59200 51642 60000 51672
rect 58341 51640 60000 51642
rect 58341 51584 58346 51640
rect 58402 51584 60000 51640
rect 58341 51582 60000 51584
rect 58341 51579 58407 51582
rect 59200 51552 60000 51582
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 0 50826 800 50856
rect 1669 50826 1735 50829
rect 0 50824 1735 50826
rect 0 50768 1674 50824
rect 1730 50768 1735 50824
rect 0 50766 1735 50768
rect 0 50736 800 50766
rect 1669 50763 1735 50766
rect 58341 50826 58407 50829
rect 59200 50826 60000 50856
rect 58341 50824 60000 50826
rect 58341 50768 58346 50824
rect 58402 50768 60000 50824
rect 58341 50766 60000 50768
rect 58341 50763 58407 50766
rect 59200 50736 60000 50766
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 0 50010 800 50040
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 1669 50010 1735 50013
rect 0 50008 1735 50010
rect 0 49952 1674 50008
rect 1730 49952 1735 50008
rect 0 49950 1735 49952
rect 0 49920 800 49950
rect 1669 49947 1735 49950
rect 58341 50010 58407 50013
rect 59200 50010 60000 50040
rect 58341 50008 60000 50010
rect 58341 49952 58346 50008
rect 58402 49952 60000 50008
rect 58341 49950 60000 49952
rect 58341 49947 58407 49950
rect 59200 49920 60000 49950
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 0 49194 800 49224
rect 1669 49194 1735 49197
rect 0 49192 1735 49194
rect 0 49136 1674 49192
rect 1730 49136 1735 49192
rect 0 49134 1735 49136
rect 0 49104 800 49134
rect 1669 49131 1735 49134
rect 58341 49194 58407 49197
rect 59200 49194 60000 49224
rect 58341 49192 60000 49194
rect 58341 49136 58346 49192
rect 58402 49136 60000 49192
rect 58341 49134 60000 49136
rect 58341 49131 58407 49134
rect 59200 49104 60000 49134
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 0 48378 800 48408
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 1669 48378 1735 48381
rect 0 48376 1735 48378
rect 0 48320 1674 48376
rect 1730 48320 1735 48376
rect 0 48318 1735 48320
rect 0 48288 800 48318
rect 1669 48315 1735 48318
rect 58341 48378 58407 48381
rect 59200 48378 60000 48408
rect 58341 48376 60000 48378
rect 58341 48320 58346 48376
rect 58402 48320 60000 48376
rect 58341 48318 60000 48320
rect 58341 48315 58407 48318
rect 59200 48288 60000 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 0 47562 800 47592
rect 1669 47562 1735 47565
rect 0 47560 1735 47562
rect 0 47504 1674 47560
rect 1730 47504 1735 47560
rect 0 47502 1735 47504
rect 0 47472 800 47502
rect 1669 47499 1735 47502
rect 58341 47562 58407 47565
rect 59200 47562 60000 47592
rect 58341 47560 60000 47562
rect 58341 47504 58346 47560
rect 58402 47504 60000 47560
rect 58341 47502 60000 47504
rect 58341 47499 58407 47502
rect 59200 47472 60000 47502
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 0 46746 800 46776
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 1669 46746 1735 46749
rect 0 46744 1735 46746
rect 0 46688 1674 46744
rect 1730 46688 1735 46744
rect 0 46686 1735 46688
rect 0 46656 800 46686
rect 1669 46683 1735 46686
rect 58341 46746 58407 46749
rect 59200 46746 60000 46776
rect 58341 46744 60000 46746
rect 58341 46688 58346 46744
rect 58402 46688 60000 46744
rect 58341 46686 60000 46688
rect 58341 46683 58407 46686
rect 59200 46656 60000 46686
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 0 45930 800 45960
rect 1669 45930 1735 45933
rect 0 45928 1735 45930
rect 0 45872 1674 45928
rect 1730 45872 1735 45928
rect 0 45870 1735 45872
rect 0 45840 800 45870
rect 1669 45867 1735 45870
rect 58341 45930 58407 45933
rect 59200 45930 60000 45960
rect 58341 45928 60000 45930
rect 58341 45872 58346 45928
rect 58402 45872 60000 45928
rect 58341 45870 60000 45872
rect 58341 45867 58407 45870
rect 59200 45840 60000 45870
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 0 45114 800 45144
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 1669 45114 1735 45117
rect 0 45112 1735 45114
rect 0 45056 1674 45112
rect 1730 45056 1735 45112
rect 0 45054 1735 45056
rect 0 45024 800 45054
rect 1669 45051 1735 45054
rect 58341 45114 58407 45117
rect 59200 45114 60000 45144
rect 58341 45112 60000 45114
rect 58341 45056 58346 45112
rect 58402 45056 60000 45112
rect 58341 45054 60000 45056
rect 58341 45051 58407 45054
rect 59200 45024 60000 45054
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 0 44298 800 44328
rect 1669 44298 1735 44301
rect 0 44296 1735 44298
rect 0 44240 1674 44296
rect 1730 44240 1735 44296
rect 0 44238 1735 44240
rect 0 44208 800 44238
rect 1669 44235 1735 44238
rect 58341 44298 58407 44301
rect 59200 44298 60000 44328
rect 58341 44296 60000 44298
rect 58341 44240 58346 44296
rect 58402 44240 60000 44296
rect 58341 44238 60000 44240
rect 58341 44235 58407 44238
rect 59200 44208 60000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 0 43482 800 43512
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 1669 43482 1735 43485
rect 0 43480 1735 43482
rect 0 43424 1674 43480
rect 1730 43424 1735 43480
rect 0 43422 1735 43424
rect 0 43392 800 43422
rect 1669 43419 1735 43422
rect 58341 43482 58407 43485
rect 59200 43482 60000 43512
rect 58341 43480 60000 43482
rect 58341 43424 58346 43480
rect 58402 43424 60000 43480
rect 58341 43422 60000 43424
rect 58341 43419 58407 43422
rect 59200 43392 60000 43422
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 0 42666 800 42696
rect 1669 42666 1735 42669
rect 0 42664 1735 42666
rect 0 42608 1674 42664
rect 1730 42608 1735 42664
rect 0 42606 1735 42608
rect 0 42576 800 42606
rect 1669 42603 1735 42606
rect 58341 42666 58407 42669
rect 59200 42666 60000 42696
rect 58341 42664 60000 42666
rect 58341 42608 58346 42664
rect 58402 42608 60000 42664
rect 58341 42606 60000 42608
rect 58341 42603 58407 42606
rect 59200 42576 60000 42606
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 0 41850 800 41880
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 1669 41850 1735 41853
rect 0 41848 1735 41850
rect 0 41792 1674 41848
rect 1730 41792 1735 41848
rect 0 41790 1735 41792
rect 0 41760 800 41790
rect 1669 41787 1735 41790
rect 58341 41850 58407 41853
rect 59200 41850 60000 41880
rect 58341 41848 60000 41850
rect 58341 41792 58346 41848
rect 58402 41792 60000 41848
rect 58341 41790 60000 41792
rect 58341 41787 58407 41790
rect 59200 41760 60000 41790
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41034 800 41064
rect 1669 41034 1735 41037
rect 0 41032 1735 41034
rect 0 40976 1674 41032
rect 1730 40976 1735 41032
rect 0 40974 1735 40976
rect 0 40944 800 40974
rect 1669 40971 1735 40974
rect 58341 41034 58407 41037
rect 59200 41034 60000 41064
rect 58341 41032 60000 41034
rect 58341 40976 58346 41032
rect 58402 40976 60000 41032
rect 58341 40974 60000 40976
rect 58341 40971 58407 40974
rect 59200 40944 60000 40974
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 0 40218 800 40248
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 1669 40218 1735 40221
rect 0 40216 1735 40218
rect 0 40160 1674 40216
rect 1730 40160 1735 40216
rect 0 40158 1735 40160
rect 0 40128 800 40158
rect 1669 40155 1735 40158
rect 58341 40218 58407 40221
rect 59200 40218 60000 40248
rect 58341 40216 60000 40218
rect 58341 40160 58346 40216
rect 58402 40160 60000 40216
rect 58341 40158 60000 40160
rect 58341 40155 58407 40158
rect 59200 40128 60000 40158
rect 57278 40020 57284 40084
rect 57348 40082 57354 40084
rect 58157 40082 58223 40085
rect 57348 40080 58223 40082
rect 57348 40024 58162 40080
rect 58218 40024 58223 40080
rect 57348 40022 58223 40024
rect 57348 40020 57354 40022
rect 58157 40019 58223 40022
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39402 800 39432
rect 1669 39402 1735 39405
rect 0 39400 1735 39402
rect 0 39344 1674 39400
rect 1730 39344 1735 39400
rect 0 39342 1735 39344
rect 0 39312 800 39342
rect 1669 39339 1735 39342
rect 58341 39402 58407 39405
rect 59200 39402 60000 39432
rect 58341 39400 60000 39402
rect 58341 39344 58346 39400
rect 58402 39344 60000 39400
rect 58341 39342 60000 39344
rect 58341 39339 58407 39342
rect 59200 39312 60000 39342
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 0 38586 800 38616
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 1669 38586 1735 38589
rect 0 38584 1735 38586
rect 0 38528 1674 38584
rect 1730 38528 1735 38584
rect 0 38526 1735 38528
rect 0 38496 800 38526
rect 1669 38523 1735 38526
rect 58341 38586 58407 38589
rect 59200 38586 60000 38616
rect 58341 38584 60000 38586
rect 58341 38528 58346 38584
rect 58402 38528 60000 38584
rect 58341 38526 60000 38528
rect 58341 38523 58407 38526
rect 59200 38496 60000 38526
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 0 37770 800 37800
rect 1669 37770 1735 37773
rect 0 37768 1735 37770
rect 0 37712 1674 37768
rect 1730 37712 1735 37768
rect 0 37710 1735 37712
rect 0 37680 800 37710
rect 1669 37707 1735 37710
rect 58341 37770 58407 37773
rect 59200 37770 60000 37800
rect 58341 37768 60000 37770
rect 58341 37712 58346 37768
rect 58402 37712 60000 37768
rect 58341 37710 60000 37712
rect 58341 37707 58407 37710
rect 59200 37680 60000 37710
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 0 36954 800 36984
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 1669 36954 1735 36957
rect 0 36952 1735 36954
rect 0 36896 1674 36952
rect 1730 36896 1735 36952
rect 0 36894 1735 36896
rect 0 36864 800 36894
rect 1669 36891 1735 36894
rect 58341 36954 58407 36957
rect 59200 36954 60000 36984
rect 58341 36952 60000 36954
rect 58341 36896 58346 36952
rect 58402 36896 60000 36952
rect 58341 36894 60000 36896
rect 58341 36891 58407 36894
rect 59200 36864 60000 36894
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 36138 800 36168
rect 1669 36138 1735 36141
rect 0 36136 1735 36138
rect 0 36080 1674 36136
rect 1730 36080 1735 36136
rect 0 36078 1735 36080
rect 0 36048 800 36078
rect 1669 36075 1735 36078
rect 58341 36138 58407 36141
rect 59200 36138 60000 36168
rect 58341 36136 60000 36138
rect 58341 36080 58346 36136
rect 58402 36080 60000 36136
rect 58341 36078 60000 36080
rect 58341 36075 58407 36078
rect 59200 36048 60000 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 0 35322 800 35352
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 1669 35322 1735 35325
rect 0 35320 1735 35322
rect 0 35264 1674 35320
rect 1730 35264 1735 35320
rect 0 35262 1735 35264
rect 0 35232 800 35262
rect 1669 35259 1735 35262
rect 58341 35322 58407 35325
rect 59200 35322 60000 35352
rect 58341 35320 60000 35322
rect 58341 35264 58346 35320
rect 58402 35264 60000 35320
rect 58341 35262 60000 35264
rect 58341 35259 58407 35262
rect 59200 35232 60000 35262
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 0 34506 800 34536
rect 1669 34506 1735 34509
rect 0 34504 1735 34506
rect 0 34448 1674 34504
rect 1730 34448 1735 34504
rect 0 34446 1735 34448
rect 0 34416 800 34446
rect 1669 34443 1735 34446
rect 57881 34506 57947 34509
rect 59200 34506 60000 34536
rect 57881 34504 60000 34506
rect 57881 34448 57886 34504
rect 57942 34448 60000 34504
rect 57881 34446 60000 34448
rect 57881 34443 57947 34446
rect 59200 34416 60000 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 0 33690 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 1669 33690 1735 33693
rect 0 33688 1735 33690
rect 0 33632 1674 33688
rect 1730 33632 1735 33688
rect 0 33630 1735 33632
rect 0 33600 800 33630
rect 1669 33627 1735 33630
rect 58433 33690 58499 33693
rect 59200 33690 60000 33720
rect 58433 33688 60000 33690
rect 58433 33632 58438 33688
rect 58494 33632 60000 33688
rect 58433 33630 60000 33632
rect 58433 33627 58499 33630
rect 59200 33600 60000 33630
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 0 32874 800 32904
rect 1669 32874 1735 32877
rect 0 32872 1735 32874
rect 0 32816 1674 32872
rect 1730 32816 1735 32872
rect 0 32814 1735 32816
rect 0 32784 800 32814
rect 1669 32811 1735 32814
rect 57881 32874 57947 32877
rect 59200 32874 60000 32904
rect 57881 32872 60000 32874
rect 57881 32816 57886 32872
rect 57942 32816 60000 32872
rect 57881 32814 60000 32816
rect 57881 32811 57947 32814
rect 59200 32784 60000 32814
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1669 32058 1735 32061
rect 0 32056 1735 32058
rect 0 32000 1674 32056
rect 1730 32000 1735 32056
rect 0 31998 1735 32000
rect 0 31968 800 31998
rect 1669 31995 1735 31998
rect 58341 32058 58407 32061
rect 59200 32058 60000 32088
rect 58341 32056 60000 32058
rect 58341 32000 58346 32056
rect 58402 32000 60000 32056
rect 58341 31998 60000 32000
rect 58341 31995 58407 31998
rect 59200 31968 60000 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 0 31242 800 31272
rect 1669 31242 1735 31245
rect 0 31240 1735 31242
rect 0 31184 1674 31240
rect 1730 31184 1735 31240
rect 0 31182 1735 31184
rect 0 31152 800 31182
rect 1669 31179 1735 31182
rect 58157 31242 58223 31245
rect 59200 31242 60000 31272
rect 58157 31240 60000 31242
rect 58157 31184 58162 31240
rect 58218 31184 60000 31240
rect 58157 31182 60000 31184
rect 58157 31179 58223 31182
rect 59200 31152 60000 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 0 30426 800 30456
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 1669 30426 1735 30429
rect 0 30424 1735 30426
rect 0 30368 1674 30424
rect 1730 30368 1735 30424
rect 0 30366 1735 30368
rect 0 30336 800 30366
rect 1669 30363 1735 30366
rect 58157 30426 58223 30429
rect 59200 30426 60000 30456
rect 58157 30424 60000 30426
rect 58157 30368 58162 30424
rect 58218 30368 60000 30424
rect 58157 30366 60000 30368
rect 58157 30363 58223 30366
rect 59200 30336 60000 30366
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 0 29610 800 29640
rect 1669 29610 1735 29613
rect 0 29608 1735 29610
rect 0 29552 1674 29608
rect 1730 29552 1735 29608
rect 0 29550 1735 29552
rect 0 29520 800 29550
rect 1669 29547 1735 29550
rect 57881 29610 57947 29613
rect 59200 29610 60000 29640
rect 57881 29608 60000 29610
rect 57881 29552 57886 29608
rect 57942 29552 60000 29608
rect 57881 29550 60000 29552
rect 57881 29547 57947 29550
rect 59200 29520 60000 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 0 28794 800 28824
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 1669 28794 1735 28797
rect 0 28792 1735 28794
rect 0 28736 1674 28792
rect 1730 28736 1735 28792
rect 0 28734 1735 28736
rect 0 28704 800 28734
rect 1669 28731 1735 28734
rect 58341 28794 58407 28797
rect 59200 28794 60000 28824
rect 58341 28792 60000 28794
rect 58341 28736 58346 28792
rect 58402 28736 60000 28792
rect 58341 28734 60000 28736
rect 58341 28731 58407 28734
rect 59200 28704 60000 28734
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 0 27978 800 28008
rect 1669 27978 1735 27981
rect 0 27976 1735 27978
rect 0 27920 1674 27976
rect 1730 27920 1735 27976
rect 0 27918 1735 27920
rect 0 27888 800 27918
rect 1669 27915 1735 27918
rect 58341 27978 58407 27981
rect 59200 27978 60000 28008
rect 58341 27976 60000 27978
rect 58341 27920 58346 27976
rect 58402 27920 60000 27976
rect 58341 27918 60000 27920
rect 58341 27915 58407 27918
rect 59200 27888 60000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 0 27162 800 27192
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 1669 27162 1735 27165
rect 0 27160 1735 27162
rect 0 27104 1674 27160
rect 1730 27104 1735 27160
rect 0 27102 1735 27104
rect 0 27072 800 27102
rect 1669 27099 1735 27102
rect 58341 27162 58407 27165
rect 59200 27162 60000 27192
rect 58341 27160 60000 27162
rect 58341 27104 58346 27160
rect 58402 27104 60000 27160
rect 58341 27102 60000 27104
rect 58341 27099 58407 27102
rect 59200 27072 60000 27102
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 0 26346 800 26376
rect 1669 26346 1735 26349
rect 0 26344 1735 26346
rect 0 26288 1674 26344
rect 1730 26288 1735 26344
rect 0 26286 1735 26288
rect 0 26256 800 26286
rect 1669 26283 1735 26286
rect 58341 26346 58407 26349
rect 59200 26346 60000 26376
rect 58341 26344 60000 26346
rect 58341 26288 58346 26344
rect 58402 26288 60000 26344
rect 58341 26286 60000 26288
rect 58341 26283 58407 26286
rect 59200 26256 60000 26286
rect 57329 26212 57395 26213
rect 57278 26210 57284 26212
rect 57238 26150 57284 26210
rect 57348 26208 57395 26212
rect 57390 26152 57395 26208
rect 57278 26148 57284 26150
rect 57348 26148 57395 26152
rect 57329 26147 57395 26148
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 0 25530 800 25560
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 1669 25530 1735 25533
rect 0 25528 1735 25530
rect 0 25472 1674 25528
rect 1730 25472 1735 25528
rect 0 25470 1735 25472
rect 0 25440 800 25470
rect 1669 25467 1735 25470
rect 57513 25530 57579 25533
rect 59200 25530 60000 25560
rect 57513 25528 60000 25530
rect 57513 25472 57518 25528
rect 57574 25472 60000 25528
rect 57513 25470 60000 25472
rect 57513 25467 57579 25470
rect 59200 25440 60000 25470
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 0 24714 800 24744
rect 1669 24714 1735 24717
rect 0 24712 1735 24714
rect 0 24656 1674 24712
rect 1730 24656 1735 24712
rect 0 24654 1735 24656
rect 0 24624 800 24654
rect 1669 24651 1735 24654
rect 58341 24714 58407 24717
rect 59200 24714 60000 24744
rect 58341 24712 60000 24714
rect 58341 24656 58346 24712
rect 58402 24656 60000 24712
rect 58341 24654 60000 24656
rect 58341 24651 58407 24654
rect 59200 24624 60000 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 0 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 1669 23898 1735 23901
rect 0 23896 1735 23898
rect 0 23840 1674 23896
rect 1730 23840 1735 23896
rect 0 23838 1735 23840
rect 0 23808 800 23838
rect 1669 23835 1735 23838
rect 58341 23898 58407 23901
rect 59200 23898 60000 23928
rect 58341 23896 60000 23898
rect 58341 23840 58346 23896
rect 58402 23840 60000 23896
rect 58341 23838 60000 23840
rect 58341 23835 58407 23838
rect 59200 23808 60000 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23082 800 23112
rect 1669 23082 1735 23085
rect 0 23080 1735 23082
rect 0 23024 1674 23080
rect 1730 23024 1735 23080
rect 0 23022 1735 23024
rect 0 22992 800 23022
rect 1669 23019 1735 23022
rect 58341 23082 58407 23085
rect 59200 23082 60000 23112
rect 58341 23080 60000 23082
rect 58341 23024 58346 23080
rect 58402 23024 60000 23080
rect 58341 23022 60000 23024
rect 58341 23019 58407 23022
rect 59200 22992 60000 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4210 22336 4526 22337
rect 0 22266 800 22296
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 1669 22266 1735 22269
rect 0 22264 1735 22266
rect 0 22208 1674 22264
rect 1730 22208 1735 22264
rect 0 22206 1735 22208
rect 0 22176 800 22206
rect 1669 22203 1735 22206
rect 58341 22266 58407 22269
rect 59200 22266 60000 22296
rect 58341 22264 60000 22266
rect 58341 22208 58346 22264
rect 58402 22208 60000 22264
rect 58341 22206 60000 22208
rect 58341 22203 58407 22206
rect 59200 22176 60000 22206
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 0 21450 800 21480
rect 1669 21450 1735 21453
rect 0 21448 1735 21450
rect 0 21392 1674 21448
rect 1730 21392 1735 21448
rect 0 21390 1735 21392
rect 0 21360 800 21390
rect 1669 21387 1735 21390
rect 58341 21450 58407 21453
rect 59200 21450 60000 21480
rect 58341 21448 60000 21450
rect 58341 21392 58346 21448
rect 58402 21392 60000 21448
rect 58341 21390 60000 21392
rect 58341 21387 58407 21390
rect 59200 21360 60000 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 0 20634 800 20664
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 1669 20634 1735 20637
rect 0 20632 1735 20634
rect 0 20576 1674 20632
rect 1730 20576 1735 20632
rect 0 20574 1735 20576
rect 0 20544 800 20574
rect 1669 20571 1735 20574
rect 58341 20634 58407 20637
rect 59200 20634 60000 20664
rect 58341 20632 60000 20634
rect 58341 20576 58346 20632
rect 58402 20576 60000 20632
rect 58341 20574 60000 20576
rect 58341 20571 58407 20574
rect 59200 20544 60000 20574
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 0 19818 800 19848
rect 1669 19818 1735 19821
rect 0 19816 1735 19818
rect 0 19760 1674 19816
rect 1730 19760 1735 19816
rect 0 19758 1735 19760
rect 0 19728 800 19758
rect 1669 19755 1735 19758
rect 58341 19818 58407 19821
rect 59200 19818 60000 19848
rect 58341 19816 60000 19818
rect 58341 19760 58346 19816
rect 58402 19760 60000 19816
rect 58341 19758 60000 19760
rect 58341 19755 58407 19758
rect 59200 19728 60000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 0 19002 800 19032
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 1669 19002 1735 19005
rect 0 19000 1735 19002
rect 0 18944 1674 19000
rect 1730 18944 1735 19000
rect 0 18942 1735 18944
rect 0 18912 800 18942
rect 1669 18939 1735 18942
rect 58341 19002 58407 19005
rect 59200 19002 60000 19032
rect 58341 19000 60000 19002
rect 58341 18944 58346 19000
rect 58402 18944 60000 19000
rect 58341 18942 60000 18944
rect 58341 18939 58407 18942
rect 59200 18912 60000 18942
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 0 18186 800 18216
rect 1669 18186 1735 18189
rect 0 18184 1735 18186
rect 0 18128 1674 18184
rect 1730 18128 1735 18184
rect 0 18126 1735 18128
rect 0 18096 800 18126
rect 1669 18123 1735 18126
rect 58341 18186 58407 18189
rect 59200 18186 60000 18216
rect 58341 18184 60000 18186
rect 58341 18128 58346 18184
rect 58402 18128 60000 18184
rect 58341 18126 60000 18128
rect 58341 18123 58407 18126
rect 59200 18096 60000 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 0 17370 800 17400
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 1669 17370 1735 17373
rect 0 17368 1735 17370
rect 0 17312 1674 17368
rect 1730 17312 1735 17368
rect 0 17310 1735 17312
rect 0 17280 800 17310
rect 1669 17307 1735 17310
rect 58341 17370 58407 17373
rect 59200 17370 60000 17400
rect 58341 17368 60000 17370
rect 58341 17312 58346 17368
rect 58402 17312 60000 17368
rect 58341 17310 60000 17312
rect 58341 17307 58407 17310
rect 59200 17280 60000 17310
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 0 16554 800 16584
rect 1669 16554 1735 16557
rect 0 16552 1735 16554
rect 0 16496 1674 16552
rect 1730 16496 1735 16552
rect 0 16494 1735 16496
rect 0 16464 800 16494
rect 1669 16491 1735 16494
rect 58341 16554 58407 16557
rect 59200 16554 60000 16584
rect 58341 16552 60000 16554
rect 58341 16496 58346 16552
rect 58402 16496 60000 16552
rect 58341 16494 60000 16496
rect 58341 16491 58407 16494
rect 59200 16464 60000 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 0 15736 1735 15738
rect 0 15680 1674 15736
rect 1730 15680 1735 15736
rect 0 15678 1735 15680
rect 0 15648 800 15678
rect 1669 15675 1735 15678
rect 58341 15738 58407 15741
rect 59200 15738 60000 15768
rect 58341 15736 60000 15738
rect 58341 15680 58346 15736
rect 58402 15680 60000 15736
rect 58341 15678 60000 15680
rect 58341 15675 58407 15678
rect 59200 15648 60000 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 0 14922 800 14952
rect 1669 14922 1735 14925
rect 0 14920 1735 14922
rect 0 14864 1674 14920
rect 1730 14864 1735 14920
rect 0 14862 1735 14864
rect 0 14832 800 14862
rect 1669 14859 1735 14862
rect 58341 14922 58407 14925
rect 59200 14922 60000 14952
rect 58341 14920 60000 14922
rect 58341 14864 58346 14920
rect 58402 14864 60000 14920
rect 58341 14862 60000 14864
rect 58341 14859 58407 14862
rect 59200 14832 60000 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 0 14106 800 14136
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 1669 14106 1735 14109
rect 0 14104 1735 14106
rect 0 14048 1674 14104
rect 1730 14048 1735 14104
rect 0 14046 1735 14048
rect 0 14016 800 14046
rect 1669 14043 1735 14046
rect 58341 14106 58407 14109
rect 59200 14106 60000 14136
rect 58341 14104 60000 14106
rect 58341 14048 58346 14104
rect 58402 14048 60000 14104
rect 58341 14046 60000 14048
rect 58341 14043 58407 14046
rect 59200 14016 60000 14046
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 0 13290 800 13320
rect 1669 13290 1735 13293
rect 0 13288 1735 13290
rect 0 13232 1674 13288
rect 1730 13232 1735 13288
rect 0 13230 1735 13232
rect 0 13200 800 13230
rect 1669 13227 1735 13230
rect 58341 13290 58407 13293
rect 59200 13290 60000 13320
rect 58341 13288 60000 13290
rect 58341 13232 58346 13288
rect 58402 13232 60000 13288
rect 58341 13230 60000 13232
rect 58341 13227 58407 13230
rect 59200 13200 60000 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 0 12474 800 12504
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 1669 12474 1735 12477
rect 0 12472 1735 12474
rect 0 12416 1674 12472
rect 1730 12416 1735 12472
rect 0 12414 1735 12416
rect 0 12384 800 12414
rect 1669 12411 1735 12414
rect 58341 12474 58407 12477
rect 59200 12474 60000 12504
rect 58341 12472 60000 12474
rect 58341 12416 58346 12472
rect 58402 12416 60000 12472
rect 58341 12414 60000 12416
rect 58341 12411 58407 12414
rect 59200 12384 60000 12414
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 0 11658 800 11688
rect 1669 11658 1735 11661
rect 0 11656 1735 11658
rect 0 11600 1674 11656
rect 1730 11600 1735 11656
rect 0 11598 1735 11600
rect 0 11568 800 11598
rect 1669 11595 1735 11598
rect 58341 11658 58407 11661
rect 59200 11658 60000 11688
rect 58341 11656 60000 11658
rect 58341 11600 58346 11656
rect 58402 11600 60000 11656
rect 58341 11598 60000 11600
rect 58341 11595 58407 11598
rect 59200 11568 60000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 0 10842 800 10872
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 1669 10842 1735 10845
rect 0 10840 1735 10842
rect 0 10784 1674 10840
rect 1730 10784 1735 10840
rect 0 10782 1735 10784
rect 0 10752 800 10782
rect 1669 10779 1735 10782
rect 57513 10842 57579 10845
rect 58433 10842 58499 10845
rect 59200 10842 60000 10872
rect 57513 10840 60000 10842
rect 57513 10784 57518 10840
rect 57574 10784 58438 10840
rect 58494 10784 60000 10840
rect 57513 10782 60000 10784
rect 57513 10779 57579 10782
rect 58433 10779 58499 10782
rect 59200 10752 60000 10782
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 0 10026 800 10056
rect 1669 10026 1735 10029
rect 0 10024 1735 10026
rect 0 9968 1674 10024
rect 1730 9968 1735 10024
rect 0 9966 1735 9968
rect 0 9936 800 9966
rect 1669 9963 1735 9966
rect 57789 10026 57855 10029
rect 59200 10026 60000 10056
rect 57789 10024 60000 10026
rect 57789 9968 57794 10024
rect 57850 9968 60000 10024
rect 57789 9966 60000 9968
rect 57789 9963 57855 9966
rect 59200 9936 60000 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 0 9210 800 9240
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 1669 9210 1735 9213
rect 0 9208 1735 9210
rect 0 9152 1674 9208
rect 1730 9152 1735 9208
rect 0 9150 1735 9152
rect 0 9120 800 9150
rect 1669 9147 1735 9150
rect 58341 9210 58407 9213
rect 59200 9210 60000 9240
rect 58341 9208 60000 9210
rect 58341 9152 58346 9208
rect 58402 9152 60000 9208
rect 58341 9150 60000 9152
rect 58341 9147 58407 9150
rect 59200 9120 60000 9150
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 0 8394 800 8424
rect 1669 8394 1735 8397
rect 0 8392 1735 8394
rect 0 8336 1674 8392
rect 1730 8336 1735 8392
rect 0 8334 1735 8336
rect 0 8304 800 8334
rect 1669 8331 1735 8334
rect 58341 8394 58407 8397
rect 59200 8394 60000 8424
rect 58341 8392 60000 8394
rect 58341 8336 58346 8392
rect 58402 8336 60000 8392
rect 58341 8334 60000 8336
rect 58341 8331 58407 8334
rect 59200 8304 60000 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 2405 7578 2471 7581
rect 0 7576 2471 7578
rect 0 7520 2410 7576
rect 2466 7520 2471 7576
rect 0 7518 2471 7520
rect 0 7488 800 7518
rect 2405 7515 2471 7518
rect 58341 7578 58407 7581
rect 59200 7578 60000 7608
rect 58341 7576 60000 7578
rect 58341 7520 58346 7576
rect 58402 7520 60000 7576
rect 58341 7518 60000 7520
rect 58341 7515 58407 7518
rect 59200 7488 60000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6762 800 6792
rect 1669 6762 1735 6765
rect 0 6760 1735 6762
rect 0 6704 1674 6760
rect 1730 6704 1735 6760
rect 0 6702 1735 6704
rect 0 6672 800 6702
rect 1669 6699 1735 6702
rect 58341 6762 58407 6765
rect 59200 6762 60000 6792
rect 58341 6760 60000 6762
rect 58341 6704 58346 6760
rect 58402 6704 60000 6760
rect 58341 6702 60000 6704
rect 58341 6699 58407 6702
rect 59200 6672 60000 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 0 5946 800 5976
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 1669 5946 1735 5949
rect 0 5944 1735 5946
rect 0 5888 1674 5944
rect 1730 5888 1735 5944
rect 0 5886 1735 5888
rect 0 5856 800 5886
rect 1669 5883 1735 5886
rect 58341 5946 58407 5949
rect 59200 5946 60000 5976
rect 58341 5944 60000 5946
rect 58341 5888 58346 5944
rect 58402 5888 60000 5944
rect 58341 5886 60000 5888
rect 58341 5883 58407 5886
rect 59200 5856 60000 5886
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 0 5130 800 5160
rect 1669 5130 1735 5133
rect 0 5128 1735 5130
rect 0 5072 1674 5128
rect 1730 5072 1735 5128
rect 0 5070 1735 5072
rect 0 5040 800 5070
rect 1669 5067 1735 5070
rect 58341 5130 58407 5133
rect 59200 5130 60000 5160
rect 58341 5128 60000 5130
rect 58341 5072 58346 5128
rect 58402 5072 60000 5128
rect 58341 5070 60000 5072
rect 58341 5067 58407 5070
rect 59200 5040 60000 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 0 4314 800 4344
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 800 4254
rect 1669 4251 1735 4254
rect 58341 4314 58407 4317
rect 59200 4314 60000 4344
rect 58341 4312 60000 4314
rect 58341 4256 58346 4312
rect 58402 4256 60000 4312
rect 58341 4254 60000 4256
rect 58341 4251 58407 4254
rect 59200 4224 60000 4254
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 57697 3498 57763 3501
rect 59200 3498 60000 3528
rect 57697 3496 60000 3498
rect 57697 3440 57702 3496
rect 57758 3440 60000 3496
rect 57697 3438 60000 3440
rect 57697 3435 57763 3438
rect 59200 3408 60000 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 55305 2682 55371 2685
rect 57513 2682 57579 2685
rect 59200 2682 60000 2712
rect 55305 2680 60000 2682
rect 55305 2624 55310 2680
rect 55366 2624 57518 2680
rect 57574 2624 60000 2680
rect 55305 2622 60000 2624
rect 55305 2619 55371 2622
rect 57513 2619 57579 2622
rect 59200 2592 60000 2622
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 56041 1866 56107 1869
rect 59200 1866 60000 1896
rect 56041 1864 60000 1866
rect 56041 1808 56046 1864
rect 56102 1808 60000 1864
rect 56041 1806 60000 1808
rect 56041 1803 56107 1806
rect 59200 1776 60000 1806
rect 56501 1050 56567 1053
rect 59200 1050 60000 1080
rect 56501 1048 60000 1050
rect 56501 992 56506 1048
rect 56562 992 60000 1048
rect 56501 990 60000 992
rect 56501 987 56567 990
rect 59200 960 60000 990
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 57284 40020 57348 40084
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 57284 26208 57348 26212
rect 57284 26152 57334 26208
rect 57334 26152 57348 26208
rect 57284 26148 57348 26152
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 57283 40084 57349 40085
rect 57283 40020 57284 40084
rect 57348 40020 57349 40084
rect 57283 40019 57349 40020
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 57286 26213 57346 40019
rect 57283 26212 57349 26213
rect 57283 26148 57284 26212
rect 57348 26148 57349 26212
rect 57283 26147 57349 26148
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 3128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__S
timestamp 1670032574
transform 1 0 2760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A0
timestamp 1670032574
transform 1 0 12420 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A1
timestamp 1670032574
transform 1 0 14260 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__S
timestamp 1670032574
transform 1 0 13800 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A0
timestamp 1670032574
transform 1 0 8280 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A1
timestamp 1670032574
transform 1 0 7728 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__S
timestamp 1670032574
transform 1 0 7360 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A0
timestamp 1670032574
transform -1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A1
timestamp 1670032574
transform 1 0 11592 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__S
timestamp 1670032574
transform 1 0 11224 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A0
timestamp 1670032574
transform 1 0 15732 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A1
timestamp 1670032574
transform 1 0 13616 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__S
timestamp 1670032574
transform 1 0 15180 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A0
timestamp 1670032574
transform -1 0 17112 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A1
timestamp 1670032574
transform 1 0 15272 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__S
timestamp 1670032574
transform 1 0 17480 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A0
timestamp 1670032574
transform -1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1670032574
transform 1 0 18216 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__S
timestamp 1670032574
transform 1 0 20608 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1
timestamp 1670032574
transform 1 0 19412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__S
timestamp 1670032574
transform 1 0 20792 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A1
timestamp 1670032574
transform -1 0 22172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__S
timestamp 1670032574
transform 1 0 23368 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A1
timestamp 1670032574
transform 1 0 19504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__S
timestamp 1670032574
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A1
timestamp 1670032574
transform 1 0 21528 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__S
timestamp 1670032574
transform 1 0 23276 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A1
timestamp 1670032574
transform 1 0 22540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__S
timestamp 1670032574
transform -1 0 23828 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1670032574
transform 1 0 38088 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1670032574
transform 1 0 38272 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A
timestamp 1670032574
transform 1 0 31372 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1670032574
transform 1 0 29532 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1670032574
transform 1 0 28244 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__C_N
timestamp 1670032574
transform 1 0 28060 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A
timestamp 1670032574
transform 1 0 28980 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A_N
timestamp 1670032574
transform 1 0 32844 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__B
timestamp 1670032574
transform 1 0 33396 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1670032574
transform 1 0 36616 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1670032574
transform 1 0 40848 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__B
timestamp 1670032574
transform 1 0 41216 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__C
timestamp 1670032574
transform -1 0 41584 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A_N
timestamp 1670032574
transform 1 0 40572 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__B
timestamp 1670032574
transform 1 0 40020 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__C
timestamp 1670032574
transform 1 0 39652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A_N
timestamp 1670032574
transform -1 0 39928 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__B
timestamp 1670032574
transform 1 0 40296 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__C
timestamp 1670032574
transform 1 0 39376 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__C
timestamp 1670032574
transform 1 0 33948 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A
timestamp 1670032574
transform 1 0 31648 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1670032574
transform 1 0 25760 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A1
timestamp 1670032574
transform 1 0 22540 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A1
timestamp 1670032574
transform -1 0 23184 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A1
timestamp 1670032574
transform 1 0 26312 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A1
timestamp 1670032574
transform 1 0 29072 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A1
timestamp 1670032574
transform -1 0 38088 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A1
timestamp 1670032574
transform -1 0 31004 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1670032574
transform 1 0 55936 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1670032574
transform 1 0 55568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__S0
timestamp 1670032574
transform -1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__S1
timestamp 1670032574
transform -1 0 57040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__S0
timestamp 1670032574
transform 1 0 57408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__S1
timestamp 1670032574
transform 1 0 56856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__S0
timestamp 1670032574
transform 1 0 57408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__S1
timestamp 1670032574
transform 1 0 56856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__S0
timestamp 1670032574
transform 1 0 57408 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__S1
timestamp 1670032574
transform 1 0 57592 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1670032574
transform 1 0 40848 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__S0
timestamp 1670032574
transform 1 0 57592 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__S1
timestamp 1670032574
transform 1 0 57040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__S0
timestamp 1670032574
transform -1 0 58420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__S1
timestamp 1670032574
transform 1 0 57408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A3
timestamp 1670032574
transform -1 0 57224 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__S0
timestamp 1670032574
transform 1 0 57408 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__S1
timestamp 1670032574
transform 1 0 56856 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A3
timestamp 1670032574
transform -1 0 58420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__S0
timestamp 1670032574
transform 1 0 57408 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__S1
timestamp 1670032574
transform 1 0 56856 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A3
timestamp 1670032574
transform -1 0 57040 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__S0
timestamp 1670032574
transform 1 0 57408 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__S1
timestamp 1670032574
transform 1 0 57592 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A3
timestamp 1670032574
transform -1 0 57040 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__S0
timestamp 1670032574
transform 1 0 57408 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__S1
timestamp 1670032574
transform 1 0 56856 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A
timestamp 1670032574
transform -1 0 53820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A3
timestamp 1670032574
transform -1 0 57776 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__S0
timestamp 1670032574
transform 1 0 55752 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__S1
timestamp 1670032574
transform 1 0 55568 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1670032574
transform 1 0 48576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A3
timestamp 1670032574
transform 1 0 57408 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__S0
timestamp 1670032574
transform 1 0 56672 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__S1
timestamp 1670032574
transform 1 0 56120 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A3
timestamp 1670032574
transform 1 0 56672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__S0
timestamp 1670032574
transform 1 0 54188 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__S1
timestamp 1670032574
transform 1 0 53820 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A3
timestamp 1670032574
transform 1 0 57408 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__S0
timestamp 1670032574
transform 1 0 56120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__S1
timestamp 1670032574
transform 1 0 55752 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A3
timestamp 1670032574
transform 1 0 57408 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__S0
timestamp 1670032574
transform 1 0 56580 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__S1
timestamp 1670032574
transform 1 0 56212 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 1670032574
transform -1 0 56948 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A3
timestamp 1670032574
transform -1 0 56672 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__S0
timestamp 1670032574
transform 1 0 54280 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__S1
timestamp 1670032574
transform 1 0 53912 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1670032574
transform -1 0 54924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A3
timestamp 1670032574
transform 1 0 57500 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__S0
timestamp 1670032574
transform 1 0 55292 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__S1
timestamp 1670032574
transform -1 0 55016 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 1670032574
transform 1 0 55752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A3
timestamp 1670032574
transform -1 0 55844 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__S0
timestamp 1670032574
transform 1 0 56580 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__S1
timestamp 1670032574
transform 1 0 56212 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 1670032574
transform -1 0 56580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1670032574
transform 1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__B
timestamp 1670032574
transform 1 0 22632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 1670032574
transform -1 0 20516 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A0
timestamp 1670032574
transform -1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A1
timestamp 1670032574
transform 1 0 5888 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__S
timestamp 1670032574
transform 1 0 5336 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A0
timestamp 1670032574
transform 1 0 7176 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A1
timestamp 1670032574
transform 1 0 8004 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__S
timestamp 1670032574
transform 1 0 6992 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A0
timestamp 1670032574
transform -1 0 10028 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A1
timestamp 1670032574
transform -1 0 10212 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__S
timestamp 1670032574
transform 1 0 10396 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A0
timestamp 1670032574
transform 1 0 8464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A1
timestamp 1670032574
transform 1 0 9108 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__S
timestamp 1670032574
transform 1 0 8464 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A0
timestamp 1670032574
transform 1 0 7360 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A1
timestamp 1670032574
transform 1 0 7544 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__S
timestamp 1670032574
transform 1 0 6624 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A0
timestamp 1670032574
transform -1 0 10120 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A1
timestamp 1670032574
transform 1 0 10120 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__S
timestamp 1670032574
transform -1 0 10672 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A0
timestamp 1670032574
transform 1 0 11592 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A1
timestamp 1670032574
transform -1 0 11224 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__S
timestamp 1670032574
transform 1 0 10672 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A0
timestamp 1670032574
transform -1 0 14996 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A1
timestamp 1670032574
transform -1 0 14444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__S
timestamp 1670032574
transform 1 0 14352 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A0
timestamp 1670032574
transform -1 0 13248 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A1
timestamp 1670032574
transform 1 0 12512 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__S
timestamp 1670032574
transform 1 0 15364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A0
timestamp 1670032574
transform 1 0 17480 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A1
timestamp 1670032574
transform 1 0 16744 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__S
timestamp 1670032574
transform 1 0 18308 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A0
timestamp 1670032574
transform 1 0 19412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A1
timestamp 1670032574
transform 1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__S
timestamp 1670032574
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A1
timestamp 1670032574
transform -1 0 19136 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__S
timestamp 1670032574
transform 1 0 20700 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A1
timestamp 1670032574
transform 1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__S
timestamp 1670032574
transform 1 0 21068 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A1
timestamp 1670032574
transform -1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__S
timestamp 1670032574
transform 1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A1
timestamp 1670032574
transform -1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__S
timestamp 1670032574
transform -1 0 22816 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A1
timestamp 1670032574
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__S
timestamp 1670032574
transform -1 0 23828 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1670032574
transform 1 0 22632 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__B
timestamp 1670032574
transform 1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A0
timestamp 1670032574
transform -1 0 1840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__S
timestamp 1670032574
transform -1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A0
timestamp 1670032574
transform 1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__S
timestamp 1670032574
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A0
timestamp 1670032574
transform -1 0 1840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__S
timestamp 1670032574
transform 1 0 4600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A0
timestamp 1670032574
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__S
timestamp 1670032574
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A0
timestamp 1670032574
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__S
timestamp 1670032574
transform 1 0 3036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A0
timestamp 1670032574
transform 1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__S
timestamp 1670032574
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A0
timestamp 1670032574
transform 1 0 3956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__S
timestamp 1670032574
transform -1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A0
timestamp 1670032574
transform 1 0 10304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__S
timestamp 1670032574
transform 1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A0
timestamp 1670032574
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A1
timestamp 1670032574
transform 1 0 19136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__S
timestamp 1670032574
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A0
timestamp 1670032574
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A1
timestamp 1670032574
transform -1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__S
timestamp 1670032574
transform 1 0 20516 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A0
timestamp 1670032574
transform 1 0 19136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A1
timestamp 1670032574
transform 1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A1
timestamp 1670032574
transform -1 0 21160 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A1
timestamp 1670032574
transform -1 0 19872 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A1
timestamp 1670032574
transform -1 0 20424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A1
timestamp 1670032574
transform 1 0 21988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A1
timestamp 1670032574
transform 1 0 21344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A_N
timestamp 1670032574
transform 1 0 21988 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__B
timestamp 1670032574
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A0
timestamp 1670032574
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__S
timestamp 1670032574
transform 1 0 2944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A0
timestamp 1670032574
transform 1 0 2944 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__S
timestamp 1670032574
transform 1 0 3956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A0
timestamp 1670032574
transform 1 0 3128 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__S
timestamp 1670032574
transform 1 0 2944 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A0
timestamp 1670032574
transform 1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__S
timestamp 1670032574
transform 1 0 2760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A0
timestamp 1670032574
transform 1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__S
timestamp 1670032574
transform 1 0 2944 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A0
timestamp 1670032574
transform 1 0 3036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__S
timestamp 1670032574
transform -1 0 2668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A0
timestamp 1670032574
transform 1 0 3128 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__S
timestamp 1670032574
transform 1 0 2760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A0
timestamp 1670032574
transform 1 0 11132 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A1
timestamp 1670032574
transform -1 0 11868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__S
timestamp 1670032574
transform 1 0 11684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A0
timestamp 1670032574
transform 1 0 15548 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A1
timestamp 1670032574
transform -1 0 15180 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__S
timestamp 1670032574
transform 1 0 14444 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A0
timestamp 1670032574
transform 1 0 18584 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A1
timestamp 1670032574
transform 1 0 18400 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__S
timestamp 1670032574
transform 1 0 19964 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A0
timestamp 1670032574
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A1
timestamp 1670032574
transform 1 0 18676 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A1
timestamp 1670032574
transform 1 0 19228 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A1
timestamp 1670032574
transform 1 0 21160 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A1
timestamp 1670032574
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A1
timestamp 1670032574
transform 1 0 21896 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A1
timestamp 1670032574
transform 1 0 21988 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A_N
timestamp 1670032574
transform -1 0 24748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__B
timestamp 1670032574
transform 1 0 23184 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1670032574
transform 1 0 20056 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A0
timestamp 1670032574
transform 1 0 3036 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__S
timestamp 1670032574
transform 1 0 2852 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A0
timestamp 1670032574
transform 1 0 5152 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__S
timestamp 1670032574
transform 1 0 4784 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A0
timestamp 1670032574
transform 1 0 3680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__S
timestamp 1670032574
transform 1 0 4232 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A0
timestamp 1670032574
transform 1 0 3128 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__S
timestamp 1670032574
transform 1 0 2852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_reg_wr_i_A
timestamp 1670032574
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout235_A
timestamp 1670032574
transform 1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout236_A
timestamp 1670032574
transform 1 0 7268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout237_A
timestamp 1670032574
transform 1 0 13616 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout238_A
timestamp 1670032574
transform 1 0 11960 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout239_A
timestamp 1670032574
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout240_A
timestamp 1670032574
transform -1 0 6532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout241_A
timestamp 1670032574
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout242_A
timestamp 1670032574
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1670032574
transform -1 0 54372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1670032574
transform -1 0 1932 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1670032574
transform -1 0 3220 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1670032574
transform -1 0 4324 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1670032574
transform -1 0 6164 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1670032574
transform -1 0 6716 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1670032574
transform -1 0 8648 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1670032574
transform -1 0 9292 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1670032574
transform -1 0 9936 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1670032574
transform -1 0 11224 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1670032574
transform -1 0 12696 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1670032574
transform -1 0 13800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1670032574
transform -1 0 15088 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1670032574
transform -1 0 16376 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1670032574
transform -1 0 17480 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1670032574
transform -1 0 18308 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1670032574
transform -1 0 19872 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1670032574
transform -1 0 20700 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1670032574
transform -1 0 22264 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1670032574
transform -1 0 23092 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1670032574
transform -1 0 24748 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1670032574
transform -1 0 25484 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1670032574
transform -1 0 26680 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1670032574
transform -1 0 28244 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1670032574
transform -1 0 29256 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1670032574
transform -1 0 31464 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1670032574
transform -1 0 32292 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1670032574
transform -1 0 33856 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1670032574
transform -1 0 34408 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1670032574
transform -1 0 35512 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1670032574
transform -1 0 36616 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1670032574
transform -1 0 38640 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1670032574
transform -1 0 38364 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1670032574
transform -1 0 41032 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1670032574
transform -1 0 41400 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1670032574
transform -1 0 43424 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1670032574
transform -1 0 44620 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1670032574
transform -1 0 45356 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1670032574
transform -1 0 47012 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1670032574
transform -1 0 47748 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1670032574
transform -1 0 49404 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1670032574
transform -1 0 50508 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1670032574
transform -1 0 51796 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1670032574
transform -1 0 52164 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1670032574
transform -1 0 54188 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1670032574
transform -1 0 54556 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1670032574
transform -1 0 56580 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1670032574
transform -1 0 56488 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1670032574
transform -1 0 56212 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1670032574
transform -1 0 24564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1670032574
transform -1 0 25576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1670032574
transform -1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1670032574
transform -1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1670032574
transform -1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1670032574
transform -1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1670032574
transform -1 0 17664 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1670032574
transform -1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1670032574
transform -1 0 18216 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1670032574
transform -1 0 21160 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1670032574
transform -1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1670032574
transform -1 0 23828 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1670032574
transform -1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1670032574
transform -1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1670032574
transform -1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1670032574
transform -1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1670032574
transform -1 0 12144 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1670032574
transform -1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1670032574
transform -1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1670032574
transform -1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1670032574
transform -1 0 15824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1670032574
transform -1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1670032574
transform -1 0 55384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1670032574
transform -1 0 55660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1670032574
transform -1 0 54096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1670032574
transform -1 0 57132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1670032574
transform -1 0 56028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1670032574
transform -1 0 56488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1670032574
transform -1 0 57776 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1670032574
transform -1 0 57592 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1670032574
transform -1 0 57224 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1670032574
transform -1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1670032574
transform -1 0 57776 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1670032574
transform -1 0 57592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1670032574
transform -1 0 57224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1670032574
transform -1 0 57776 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1670032574
transform -1 0 56948 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1670032574
transform -1 0 56396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1670032574
transform -1 0 58420 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1670032574
transform -1 0 57776 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1670032574
transform -1 0 55936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1670032574
transform -1 0 56488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1670032574
transform -1 0 56488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1670032574
transform -1 0 57040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1670032574
transform -1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1670032574
transform -1 0 57224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1670032574
transform -1 0 56488 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1670032574
transform -1 0 58420 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1670032574
transform -1 0 57592 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1670032574
transform -1 0 57592 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1670032574
transform -1 0 58420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1670032574
transform -1 0 57776 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1670032574
transform -1 0 57224 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1670032574
transform -1 0 57592 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1670032574
transform -1 0 57776 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1670032574
transform -1 0 57224 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1670032574
transform -1 0 57592 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1670032574
transform -1 0 57592 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1670032574
transform -1 0 57592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1670032574
transform -1 0 58420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1670032574
transform -1 0 57224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1670032574
transform -1 0 57776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1670032574
transform -1 0 57776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1670032574
transform -1 0 57592 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1670032574
transform -1 0 57776 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1670032574
transform -1 0 57592 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1670032574
transform -1 0 57776 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1670032574
transform -1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1670032574
transform -1 0 57592 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1670032574
transform -1 0 57776 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1670032574
transform -1 0 57776 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1670032574
transform -1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1670032574
transform -1 0 57592 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1670032574
transform -1 0 57776 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1670032574
transform -1 0 57776 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1670032574
transform -1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1670032574
transform -1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1670032574
transform -1 0 57776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1670032574
transform -1 0 57776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1670032574
transform -1 0 57592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1670032574
transform -1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1670032574
transform -1 0 57776 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1670032574
transform -1 0 57776 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1670032574
transform -1 0 57224 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1670032574
transform -1 0 56764 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1670032574
transform -1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1670032574
transform -1 0 57592 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1670032574
transform -1 0 57776 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input138_A
timestamp 1670032574
transform -1 0 57776 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input139_A
timestamp 1670032574
transform -1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input140_A
timestamp 1670032574
transform -1 0 57592 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input141_A
timestamp 1670032574
transform -1 0 57776 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input142_A
timestamp 1670032574
transform -1 0 55936 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input143_A
timestamp 1670032574
transform -1 0 57316 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input144_A
timestamp 1670032574
transform -1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input145_A
timestamp 1670032574
transform -1 0 36064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output147_A
timestamp 1670032574
transform -1 0 27416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output148_A
timestamp 1670032574
transform 1 0 28704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output149_A
timestamp 1670032574
transform 1 0 29808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1670032574
transform 1 0 30912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output151_A
timestamp 1670032574
transform -1 0 32476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output152_A
timestamp 1670032574
transform 1 0 33120 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output154_A
timestamp 1670032574
transform 1 0 3496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output155_A
timestamp 1670032574
transform 1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output156_A
timestamp 1670032574
transform 1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output157_A
timestamp 1670032574
transform 1 0 2944 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output158_A
timestamp 1670032574
transform 1 0 3312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output159_A
timestamp 1670032574
transform -1 0 2484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output167_A
timestamp 1670032574
transform 1 0 2300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1670032574
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1670032574
transform 1 0 2300 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1670032574
transform -1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output172_A
timestamp 1670032574
transform -1 0 2484 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output173_A
timestamp 1670032574
transform 1 0 2300 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1670032574
transform 1 0 2300 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1670032574
transform -1 0 2484 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output182_A
timestamp 1670032574
transform 1 0 3956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output183_A
timestamp 1670032574
transform 1 0 3404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output184_A
timestamp 1670032574
transform 1 0 2300 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output186_A
timestamp 1670032574
transform 1 0 2300 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output187_A
timestamp 1670032574
transform -1 0 2484 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output188_A
timestamp 1670032574
transform -1 0 2484 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output189_A
timestamp 1670032574
transform 1 0 2300 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output190_A
timestamp 1670032574
transform 1 0 2300 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output191_A
timestamp 1670032574
transform -1 0 2484 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output196_A
timestamp 1670032574
transform 1 0 2300 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output197_A
timestamp 1670032574
transform 1 0 2300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output198_A
timestamp 1670032574
transform -1 0 2484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output199_A
timestamp 1670032574
transform -1 0 2484 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output200_A
timestamp 1670032574
transform 1 0 2300 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output201_A
timestamp 1670032574
transform -1 0 2484 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output202_A
timestamp 1670032574
transform 1 0 2300 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output203_A
timestamp 1670032574
transform -1 0 2484 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output204_A
timestamp 1670032574
transform -1 0 2484 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output205_A
timestamp 1670032574
transform 1 0 2300 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output206_A
timestamp 1670032574
transform 1 0 2300 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output207_A
timestamp 1670032574
transform -1 0 2484 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output208_A
timestamp 1670032574
transform 1 0 2300 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output209_A
timestamp 1670032574
transform 1 0 2300 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output210_A
timestamp 1670032574
transform -1 0 2484 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1670032574
transform -1 0 2484 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output212_A
timestamp 1670032574
transform 1 0 2300 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output213_A
timestamp 1670032574
transform 1 0 2300 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output214_A
timestamp 1670032574
transform -1 0 2484 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output215_A
timestamp 1670032574
transform -1 0 2484 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output216_A
timestamp 1670032574
transform 1 0 2300 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output217_A
timestamp 1670032574
transform 1 0 37812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output218_A
timestamp 1670032574
transform 1 0 38548 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output219_A
timestamp 1670032574
transform 1 0 39284 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output221_A
timestamp 1670032574
transform 1 0 41768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output223_A
timestamp 1670032574
transform 1 0 43700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output226_A
timestamp 1670032574
transform 1 0 44712 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output227_A
timestamp 1670032574
transform 1 0 45816 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1670032574
transform 1 0 49496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output231_A
timestamp 1670032574
transform 1 0 50692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output232_A
timestamp 1670032574
transform 1 0 51428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10
timestamp 1670032574
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 2668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp 1670032574
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1670032574
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1670032574
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1670032574
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1670032574
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66
timestamp 1670032574
transform 1 0 7176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1670032574
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1670032574
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91
timestamp 1670032574
transform 1 0 9476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97
timestamp 1670032574
transform 1 0 10028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1670032574
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1670032574
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1670032574
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1670032574
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126
timestamp 1670032574
transform 1 0 12696 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1670032574
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1670032574
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1670032574
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_150
timestamp 1670032574
transform 1 0 14904 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1670032574
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1670032574
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_175
timestamp 1670032574
transform 1 0 17204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_181
timestamp 1670032574
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1670032574
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp 1670032574
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1670032574
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_216
timestamp 1670032574
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1670032574
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1670032574
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_229
timestamp 1670032574
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_233
timestamp 1670032574
transform 1 0 22540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_241
timestamp 1670032574
transform 1 0 23276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1670032574
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1670032574
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1670032574
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_261
timestamp 1670032574
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 1670032574
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_272
timestamp 1670032574
transform 1 0 26128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1670032574
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1670032574
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_294
timestamp 1670032574
transform 1 0 28152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1670032574
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1670032574
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_313
timestamp 1670032574
transform 1 0 29900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_318
timestamp 1670032574
transform 1 0 30360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1670032574
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1670032574
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_343
timestamp 1670032574
transform 1 0 32660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_349
timestamp 1670032574
transform 1 0 33212 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_354
timestamp 1670032574
transform 1 0 33672 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1670032574
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1670032574
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_376
timestamp 1670032574
transform 1 0 35696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_386
timestamp 1670032574
transform 1 0 36616 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1670032574
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_399
timestamp 1670032574
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_407
timestamp 1670032574
transform 1 0 38548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1670032574
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1670032574
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1670032574
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_427
timestamp 1670032574
transform 1 0 40388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1670032574
transform 1 0 40940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_438
timestamp 1670032574
transform 1 0 41400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1670032574
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1670032574
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_455
timestamp 1670032574
transform 1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_463
timestamp 1670032574
transform 1 0 43700 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_469
timestamp 1670032574
transform 1 0 44252 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1670032574
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1670032574
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_481
timestamp 1670032574
transform 1 0 45356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_486
timestamp 1670032574
transform 1 0 45816 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1670032574
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1670032574
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_511
timestamp 1670032574
transform 1 0 48116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_517
timestamp 1670032574
transform 1 0 48668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_522
timestamp 1670032574
transform 1 0 49128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_528
timestamp 1670032574
transform 1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1670032574
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1670032574
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_547
timestamp 1670032574
transform 1 0 51428 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_553
timestamp 1670032574
transform 1 0 51980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1670032574
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_561
timestamp 1670032574
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_565
timestamp 1670032574
transform 1 0 53084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_570
timestamp 1670032574
transform 1 0 53544 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_582
timestamp 1670032574
transform 1 0 54648 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1670032574
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_595
timestamp 1670032574
transform 1 0 55844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_601
timestamp 1670032574
transform 1 0 56396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_605
timestamp 1670032574
transform 1 0 56764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1670032574
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1670032574
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1670032574
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1670032574
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_8
timestamp 1670032574
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1670032574
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_28
timestamp 1670032574
transform 1 0 3680 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1670032574
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1670032574
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1670032574
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1670032574
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1670032574
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_101
timestamp 1670032574
transform 1 0 10396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_107
timestamp 1670032574
transform 1 0 10948 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1670032574
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1670032574
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1670032574
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1670032574
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_145
timestamp 1670032574
transform 1 0 14444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_151
timestamp 1670032574
transform 1 0 14996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_154
timestamp 1670032574
transform 1 0 15272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_160
timestamp 1670032574
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1670032574
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1670032574
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_191
timestamp 1670032574
transform 1 0 18676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_205
timestamp 1670032574
transform 1 0 19964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_212
timestamp 1670032574
transform 1 0 20608 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1670032574
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1670032574
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_232
timestamp 1670032574
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1670032574
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_247
timestamp 1670032574
transform 1 0 23828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_255
timestamp 1670032574
transform 1 0 24564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_263
timestamp 1670032574
transform 1 0 25300 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_266 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 25576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1670032574
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp 1670032574
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1670032574
transform 1 0 27416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_294
timestamp 1670032574
transform 1 0 28152 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_302
timestamp 1670032574
transform 1 0 28888 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_310
timestamp 1670032574
transform 1 0 29624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_314
timestamp 1670032574
transform 1 0 29992 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_322
timestamp 1670032574
transform 1 0 30728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_326
timestamp 1670032574
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1670032574
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1670032574
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_341
timestamp 1670032574
transform 1 0 32476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_347
timestamp 1670032574
transform 1 0 33028 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_350
timestamp 1670032574
transform 1 0 33304 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_362
timestamp 1670032574
transform 1 0 34408 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_374
timestamp 1670032574
transform 1 0 35512 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_380
timestamp 1670032574
transform 1 0 36064 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1670032574
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_401
timestamp 1670032574
transform 1 0 37996 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_409
timestamp 1670032574
transform 1 0 38732 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1670032574
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1670032574
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1670032574
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1670032574
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1670032574
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_461
timestamp 1670032574
transform 1 0 43516 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_465
timestamp 1670032574
transform 1 0 43884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_473
timestamp 1670032574
transform 1 0 44620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_476
timestamp 1670032574
transform 1 0 44896 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_484
timestamp 1670032574
transform 1 0 45632 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_488
timestamp 1670032574
transform 1 0 46000 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1670032574
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1670032574
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1670032574
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_529
timestamp 1670032574
transform 1 0 49772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_537
timestamp 1670032574
transform 1 0 50508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_541
timestamp 1670032574
transform 1 0 50876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_549
timestamp 1670032574
transform 1 0 51612 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1670032574
transform 1 0 52348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_561
timestamp 1670032574
transform 1 0 52716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_569
timestamp 1670032574
transform 1 0 53452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_573
timestamp 1670032574
transform 1 0 53820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_579
timestamp 1670032574
transform 1 0 54372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_585
timestamp 1670032574
transform 1 0 54924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_593
timestamp 1670032574
transform 1 0 55660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_600
timestamp 1670032574
transform 1 0 56304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_607
timestamp 1670032574
transform 1 0 56948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1670032574
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_617
timestamp 1670032574
transform 1 0 57868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_622
timestamp 1670032574
transform 1 0 58328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1670032574
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_8
timestamp 1670032574
transform 1 0 1840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1670032574
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1670032574
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1670032574
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_34
timestamp 1670032574
transform 1 0 4232 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1670032574
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1670032574
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_74
timestamp 1670032574
transform 1 0 7912 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1670032574
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1670032574
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1670032574
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_112
timestamp 1670032574
transform 1 0 11408 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_124
timestamp 1670032574
transform 1 0 12512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1670032574
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1670032574
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1670032574
transform 1 0 14812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_155
timestamp 1670032574
transform 1 0 15364 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1670032574
transform 1 0 16100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1670032574
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_190
timestamp 1670032574
transform 1 0 18584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1670032574
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp 1670032574
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_203
timestamp 1670032574
transform 1 0 19780 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_213
timestamp 1670032574
transform 1 0 20700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1670032574
transform 1 0 21252 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_222
timestamp 1670032574
transform 1 0 21528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1670032574
transform 1 0 22172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1670032574
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1670032574
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1670032574
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1670032574
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1670032574
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1670032574
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1670032574
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1670032574
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1670032574
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1670032574
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1670032574
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1670032574
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1670032574
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1670032574
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1670032574
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1670032574
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1670032574
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1670032574
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1670032574
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1670032574
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_421
timestamp 1670032574
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_428
timestamp 1670032574
transform 1 0 40480 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_434
timestamp 1670032574
transform 1 0 41032 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_446
timestamp 1670032574
transform 1 0 42136 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_458
timestamp 1670032574
transform 1 0 43240 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1670032574
transform 1 0 44344 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1670032574
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1670032574
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_501
timestamp 1670032574
transform 1 0 47196 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1670032574
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_518
timestamp 1670032574
transform 1 0 48760 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_530
timestamp 1670032574
transform 1 0 49864 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1670032574
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1670032574
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1670032574
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_569
timestamp 1670032574
transform 1 0 53452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_573
timestamp 1670032574
transform 1 0 53820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_576
timestamp 1670032574
transform 1 0 54096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_583
timestamp 1670032574
transform 1 0 54740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1670032574
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_589
timestamp 1670032574
transform 1 0 55292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_594
timestamp 1670032574
transform 1 0 55752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_601
timestamp 1670032574
transform 1 0 56396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_608
timestamp 1670032574
transform 1 0 57040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_615
timestamp 1670032574
transform 1 0 57684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_622
timestamp 1670032574
transform 1 0 58328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1670032574
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1670032574
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_21
timestamp 1670032574
transform 1 0 3036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp 1670032574
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_34
timestamp 1670032574
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_40
timestamp 1670032574
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1670032574
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1670032574
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_63
timestamp 1670032574
transform 1 0 6900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_75
timestamp 1670032574
transform 1 0 8004 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_87
timestamp 1670032574
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_99
timestamp 1670032574
transform 1 0 10212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1670032574
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1670032574
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1670032574
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1670032574
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1670032574
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1670032574
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1670032574
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1670032574
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_177
timestamp 1670032574
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_180
timestamp 1670032574
transform 1 0 17664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_186
timestamp 1670032574
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_192
timestamp 1670032574
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_198
timestamp 1670032574
transform 1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_211
timestamp 1670032574
transform 1 0 20516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp 1670032574
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1670032574
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_229
timestamp 1670032574
transform 1 0 22172 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_242
timestamp 1670032574
transform 1 0 23368 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_254
timestamp 1670032574
transform 1 0 24472 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_266
timestamp 1670032574
transform 1 0 25576 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1670032574
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1670032574
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1670032574
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1670032574
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1670032574
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1670032574
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1670032574
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1670032574
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1670032574
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1670032574
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1670032574
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1670032574
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1670032574
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1670032574
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1670032574
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1670032574
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1670032574
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1670032574
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1670032574
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1670032574
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1670032574
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1670032574
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1670032574
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1670032574
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1670032574
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1670032574
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1670032574
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1670032574
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1670032574
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1670032574
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1670032574
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1670032574
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1670032574
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_585
timestamp 1670032574
transform 1 0 54924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_590
timestamp 1670032574
transform 1 0 55384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_596
timestamp 1670032574
transform 1 0 55936 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_604
timestamp 1670032574
transform 1 0 56672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_607
timestamp 1670032574
transform 1 0 56948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_614
timestamp 1670032574
transform 1 0 57592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1670032574
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_622
timestamp 1670032574
transform 1 0 58328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1670032574
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1670032574
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1670032574
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1670032574
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1670032574
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1670032574
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1670032574
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1670032574
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1670032574
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1670032574
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1670032574
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1670032574
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1670032574
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1670032574
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1670032574
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1670032574
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1670032574
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1670032574
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1670032574
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1670032574
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1670032574
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1670032574
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1670032574
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_201
timestamp 1670032574
transform 1 0 19596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1670032574
transform 1 0 19872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_210
timestamp 1670032574
transform 1 0 20424 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_218
timestamp 1670032574
transform 1 0 21160 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1670032574
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_236
timestamp 1670032574
transform 1 0 22816 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1670032574
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1670032574
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1670032574
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1670032574
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1670032574
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1670032574
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1670032574
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1670032574
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1670032574
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1670032574
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1670032574
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1670032574
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1670032574
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1670032574
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1670032574
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1670032574
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1670032574
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1670032574
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1670032574
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1670032574
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1670032574
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1670032574
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1670032574
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1670032574
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1670032574
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1670032574
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1670032574
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1670032574
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1670032574
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1670032574
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1670032574
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1670032574
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1670032574
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1670032574
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1670032574
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1670032574
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1670032574
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_589
timestamp 1670032574
transform 1 0 55292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_597
timestamp 1670032574
transform 1 0 56028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_603
timestamp 1670032574
transform 1 0 56580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_609
timestamp 1670032574
transform 1 0 57132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_616
timestamp 1670032574
transform 1 0 57776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1670032574
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1670032574
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1670032574
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1670032574
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1670032574
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1670032574
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1670032574
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1670032574
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1670032574
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1670032574
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1670032574
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1670032574
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1670032574
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1670032574
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1670032574
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1670032574
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1670032574
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1670032574
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1670032574
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1670032574
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1670032574
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1670032574
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1670032574
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1670032574
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1670032574
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_233
timestamp 1670032574
transform 1 0 22540 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_236
timestamp 1670032574
transform 1 0 22816 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_248
timestamp 1670032574
transform 1 0 23920 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_260
timestamp 1670032574
transform 1 0 25024 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_272
timestamp 1670032574
transform 1 0 26128 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1670032574
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1670032574
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1670032574
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1670032574
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1670032574
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1670032574
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1670032574
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1670032574
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1670032574
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1670032574
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1670032574
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1670032574
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1670032574
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1670032574
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1670032574
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1670032574
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1670032574
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1670032574
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1670032574
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1670032574
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1670032574
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1670032574
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1670032574
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1670032574
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1670032574
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1670032574
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1670032574
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1670032574
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1670032574
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1670032574
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1670032574
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1670032574
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1670032574
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_597
timestamp 1670032574
transform 1 0 56028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_602
timestamp 1670032574
transform 1 0 56488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_608
timestamp 1670032574
transform 1 0 57040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_614
timestamp 1670032574
transform 1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_617
timestamp 1670032574
transform 1 0 57868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1670032574
transform 1 0 58420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1670032574
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_9
timestamp 1670032574
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1670032574
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1670032574
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1670032574
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1670032574
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_69
timestamp 1670032574
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1670032574
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1670032574
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1670032574
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_118
timestamp 1670032574
transform 1 0 11960 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp 1670032574
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1670032574
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1670032574
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1670032574
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1670032574
transform 1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1670032574
transform 1 0 16652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_190
timestamp 1670032574
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1670032574
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1670032574
transform 1 0 20608 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_218
timestamp 1670032574
transform 1 0 21160 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1670032574
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_236
timestamp 1670032574
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_242
timestamp 1670032574
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1670032574
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1670032574
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1670032574
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1670032574
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1670032574
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1670032574
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1670032574
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1670032574
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1670032574
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1670032574
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1670032574
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1670032574
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1670032574
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1670032574
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1670032574
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1670032574
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1670032574
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1670032574
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1670032574
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1670032574
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1670032574
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1670032574
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1670032574
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1670032574
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1670032574
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1670032574
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1670032574
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1670032574
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1670032574
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1670032574
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1670032574
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1670032574
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1670032574
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1670032574
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1670032574
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1670032574
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1670032574
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1670032574
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_601
timestamp 1670032574
transform 1 0 56396 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_623
timestamp 1670032574
transform 1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1670032574
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_9
timestamp 1670032574
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1670032574
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_24
timestamp 1670032574
transform 1 0 3312 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_36
timestamp 1670032574
transform 1 0 4416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1670032574
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1670032574
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1670032574
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_96
timestamp 1670032574
transform 1 0 9936 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1670032574
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1670032574
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1670032574
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1670032574
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1670032574
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1670032574
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1670032574
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1670032574
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1670032574
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_200
timestamp 1670032574
transform 1 0 19504 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_207
timestamp 1670032574
transform 1 0 20148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1670032574
transform 1 0 21252 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1670032574
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1670032574
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_234
timestamp 1670032574
transform 1 0 22632 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_247
timestamp 1670032574
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_253
timestamp 1670032574
transform 1 0 24380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_265
timestamp 1670032574
transform 1 0 25484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1670032574
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1670032574
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1670032574
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1670032574
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1670032574
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1670032574
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1670032574
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1670032574
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1670032574
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1670032574
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1670032574
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1670032574
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1670032574
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1670032574
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1670032574
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1670032574
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1670032574
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1670032574
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1670032574
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1670032574
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1670032574
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1670032574
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1670032574
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1670032574
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1670032574
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1670032574
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1670032574
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1670032574
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1670032574
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1670032574
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1670032574
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1670032574
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1670032574
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_585
timestamp 1670032574
transform 1 0 54924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_593
timestamp 1670032574
transform 1 0 55660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_596
timestamp 1670032574
transform 1 0 55936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_602
timestamp 1670032574
transform 1 0 56488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_608
timestamp 1670032574
transform 1 0 57040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_614
timestamp 1670032574
transform 1 0 57592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_617
timestamp 1670032574
transform 1 0 57868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 1670032574
transform 1 0 58420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1670032574
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1670032574
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1670032574
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1670032574
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp 1670032574
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_52
timestamp 1670032574
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_64
timestamp 1670032574
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1670032574
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1670032574
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1670032574
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1670032574
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1670032574
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1670032574
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1670032574
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1670032574
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1670032574
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1670032574
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1670032574
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_189
timestamp 1670032574
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1670032574
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1670032574
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_208
timestamp 1670032574
transform 1 0 20240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_214
timestamp 1670032574
transform 1 0 20792 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_221
timestamp 1670032574
transform 1 0 21436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_234
timestamp 1670032574
transform 1 0 22632 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1670032574
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1670032574
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_257
timestamp 1670032574
transform 1 0 24748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_269
timestamp 1670032574
transform 1 0 25852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_281
timestamp 1670032574
transform 1 0 26956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_293
timestamp 1670032574
transform 1 0 28060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1670032574
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1670032574
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1670032574
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1670032574
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1670032574
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1670032574
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1670032574
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1670032574
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1670032574
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1670032574
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1670032574
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1670032574
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1670032574
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1670032574
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1670032574
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1670032574
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1670032574
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1670032574
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1670032574
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1670032574
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1670032574
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1670032574
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1670032574
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1670032574
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1670032574
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1670032574
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1670032574
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1670032574
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1670032574
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1670032574
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1670032574
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_589
timestamp 1670032574
transform 1 0 55292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_614
timestamp 1670032574
transform 1 0 57592 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_623
timestamp 1670032574
transform 1 0 58420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1670032574
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_20
timestamp 1670032574
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1670032574
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1670032574
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1670032574
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1670032574
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1670032574
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1670032574
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1670032574
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1670032574
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1670032574
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1670032574
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1670032574
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1670032574
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1670032574
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1670032574
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1670032574
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_192
timestamp 1670032574
transform 1 0 18768 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_198
timestamp 1670032574
transform 1 0 19320 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_210
timestamp 1670032574
transform 1 0 20424 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1670032574
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1670032574
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_229
timestamp 1670032574
transform 1 0 22172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1670032574
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_250
timestamp 1670032574
transform 1 0 24104 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_262
timestamp 1670032574
transform 1 0 25208 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_274
timestamp 1670032574
transform 1 0 26312 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1670032574
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1670032574
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1670032574
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1670032574
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1670032574
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1670032574
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1670032574
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1670032574
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1670032574
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1670032574
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1670032574
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1670032574
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1670032574
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1670032574
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1670032574
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1670032574
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1670032574
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1670032574
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1670032574
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1670032574
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1670032574
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1670032574
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1670032574
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1670032574
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1670032574
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1670032574
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1670032574
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1670032574
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1670032574
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1670032574
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1670032574
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1670032574
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1670032574
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_597
timestamp 1670032574
transform 1 0 56028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_602
timestamp 1670032574
transform 1 0 56488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_608
timestamp 1670032574
transform 1 0 57040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1670032574
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_617
timestamp 1670032574
transform 1 0 57868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_623
timestamp 1670032574
transform 1 0 58420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1670032574
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1670032574
transform 1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_17
timestamp 1670032574
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1670032574
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1670032574
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1670032574
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp 1670032574
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_64
timestamp 1670032574
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1670032574
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1670032574
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1670032574
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1670032574
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1670032574
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1670032574
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1670032574
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1670032574
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1670032574
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1670032574
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1670032574
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_189
timestamp 1670032574
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1670032574
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1670032574
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_203
timestamp 1670032574
transform 1 0 19780 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_215
timestamp 1670032574
transform 1 0 20884 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_221
timestamp 1670032574
transform 1 0 21436 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_224
timestamp 1670032574
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_237
timestamp 1670032574
transform 1 0 22908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1670032574
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1670032574
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1670032574
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1670032574
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1670032574
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1670032574
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1670032574
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1670032574
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1670032574
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1670032574
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1670032574
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1670032574
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1670032574
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1670032574
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1670032574
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1670032574
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1670032574
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1670032574
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1670032574
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1670032574
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1670032574
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1670032574
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1670032574
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1670032574
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1670032574
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1670032574
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1670032574
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1670032574
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1670032574
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1670032574
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1670032574
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1670032574
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1670032574
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1670032574
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1670032574
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1670032574
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1670032574
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1670032574
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1670032574
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_601
timestamp 1670032574
transform 1 0 56396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_623
timestamp 1670032574
transform 1 0 58420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1670032574
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_9
timestamp 1670032574
transform 1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1670032574
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_19
timestamp 1670032574
transform 1 0 2852 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_25
timestamp 1670032574
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_37
timestamp 1670032574
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1670032574
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1670032574
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1670032574
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_69
timestamp 1670032574
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_95
timestamp 1670032574
transform 1 0 9844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1670032574
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1670032574
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1670032574
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_135
timestamp 1670032574
transform 1 0 13524 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_147
timestamp 1670032574
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1670032574
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1670032574
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1670032574
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_181
timestamp 1670032574
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_187
timestamp 1670032574
transform 1 0 18308 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_194
timestamp 1670032574
transform 1 0 18952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1670032574
transform 1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1670032574
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1670032574
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp 1670032574
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_234
timestamp 1670032574
transform 1 0 22632 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_246
timestamp 1670032574
transform 1 0 23736 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_258
timestamp 1670032574
transform 1 0 24840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_270
timestamp 1670032574
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1670032574
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1670032574
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1670032574
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1670032574
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1670032574
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1670032574
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1670032574
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1670032574
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1670032574
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1670032574
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1670032574
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1670032574
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1670032574
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1670032574
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1670032574
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1670032574
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1670032574
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1670032574
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1670032574
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1670032574
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1670032574
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1670032574
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1670032574
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1670032574
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1670032574
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1670032574
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1670032574
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1670032574
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1670032574
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1670032574
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1670032574
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1670032574
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1670032574
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1670032574
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_597
timestamp 1670032574
transform 1 0 56028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_605
timestamp 1670032574
transform 1 0 56764 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_608
timestamp 1670032574
transform 1 0 57040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1670032574
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_617
timestamp 1670032574
transform 1 0 57868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_623
timestamp 1670032574
transform 1 0 58420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1670032574
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_11
timestamp 1670032574
transform 1 0 2116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1670032574
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1670032574
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1670032574
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_33
timestamp 1670032574
transform 1 0 4140 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_61
timestamp 1670032574
transform 1 0 6716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_73
timestamp 1670032574
transform 1 0 7820 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1670032574
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1670032574
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_96
timestamp 1670032574
transform 1 0 9936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1670032574
transform 1 0 10488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_106
timestamp 1670032574
transform 1 0 10856 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_130
timestamp 1670032574
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1670032574
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1670032574
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1670032574
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1670032574
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1670032574
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1670032574
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1670032574
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1670032574
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_211
timestamp 1670032574
transform 1 0 20516 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_217
timestamp 1670032574
transform 1 0 21068 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_225
timestamp 1670032574
transform 1 0 21804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1670032574
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_241
timestamp 1670032574
transform 1 0 23276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1670032574
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1670032574
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1670032574
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1670032574
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1670032574
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1670032574
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1670032574
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1670032574
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1670032574
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1670032574
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1670032574
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1670032574
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1670032574
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1670032574
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1670032574
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1670032574
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1670032574
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1670032574
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1670032574
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1670032574
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1670032574
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1670032574
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1670032574
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1670032574
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1670032574
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1670032574
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1670032574
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1670032574
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1670032574
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1670032574
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1670032574
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1670032574
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1670032574
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1670032574
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1670032574
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1670032574
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1670032574
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1670032574
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_601
timestamp 1670032574
transform 1 0 56396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_607
timestamp 1670032574
transform 1 0 56948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_610
timestamp 1670032574
transform 1 0 57224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_616
timestamp 1670032574
transform 1 0 57776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_623
timestamp 1670032574
transform 1 0 58420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1670032574
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_20
timestamp 1670032574
transform 1 0 2944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1670032574
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_33
timestamp 1670032574
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1670032574
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1670032574
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1670032574
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_63
timestamp 1670032574
transform 1 0 6900 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1670032574
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1670032574
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_93
timestamp 1670032574
transform 1 0 9660 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_98
timestamp 1670032574
transform 1 0 10120 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1670032574
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1670032574
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1670032574
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_124
timestamp 1670032574
transform 1 0 12512 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_136
timestamp 1670032574
transform 1 0 13616 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_148
timestamp 1670032574
transform 1 0 14720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1670032574
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1670032574
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1670032574
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_193
timestamp 1670032574
transform 1 0 18860 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_199
timestamp 1670032574
transform 1 0 19412 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_202
timestamp 1670032574
transform 1 0 19688 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1670032574
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1670032574
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1670032574
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_231
timestamp 1670032574
transform 1 0 22356 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_235
timestamp 1670032574
transform 1 0 22724 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_247
timestamp 1670032574
transform 1 0 23828 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_259
timestamp 1670032574
transform 1 0 24932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1670032574
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1670032574
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1670032574
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1670032574
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1670032574
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1670032574
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1670032574
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1670032574
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1670032574
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1670032574
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1670032574
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1670032574
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1670032574
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1670032574
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1670032574
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1670032574
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1670032574
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1670032574
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1670032574
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1670032574
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1670032574
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1670032574
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1670032574
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1670032574
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1670032574
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1670032574
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1670032574
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1670032574
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1670032574
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1670032574
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1670032574
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1670032574
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1670032574
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1670032574
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_585
timestamp 1670032574
transform 1 0 54924 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_591
timestamp 1670032574
transform 1 0 55476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_594
timestamp 1670032574
transform 1 0 55752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_604
timestamp 1670032574
transform 1 0 56672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_614
timestamp 1670032574
transform 1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_617
timestamp 1670032574
transform 1 0 57868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_623
timestamp 1670032574
transform 1 0 58420 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1670032574
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1670032574
transform 1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1670032574
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1670032574
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1670032574
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1670032574
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1670032574
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1670032574
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1670032574
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1670032574
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1670032574
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1670032574
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1670032574
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1670032574
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1670032574
transform 1 0 11868 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_120
timestamp 1670032574
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1670032574
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1670032574
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_153
timestamp 1670032574
transform 1 0 15180 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_161
timestamp 1670032574
transform 1 0 15916 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_185
timestamp 1670032574
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1670032574
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1670032574
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1670032574
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_205
timestamp 1670032574
transform 1 0 19964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_217
timestamp 1670032574
transform 1 0 21068 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_225
timestamp 1670032574
transform 1 0 21804 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_229
timestamp 1670032574
transform 1 0 22172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_242
timestamp 1670032574
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1670032574
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1670032574
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1670032574
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1670032574
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1670032574
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1670032574
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1670032574
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1670032574
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1670032574
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1670032574
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1670032574
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1670032574
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1670032574
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1670032574
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1670032574
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1670032574
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1670032574
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1670032574
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1670032574
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1670032574
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1670032574
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1670032574
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1670032574
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1670032574
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1670032574
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1670032574
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1670032574
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1670032574
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1670032574
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1670032574
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1670032574
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1670032574
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1670032574
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1670032574
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1670032574
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1670032574
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1670032574
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1670032574
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_601
timestamp 1670032574
transform 1 0 56396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_620
timestamp 1670032574
transform 1 0 58144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_624
timestamp 1670032574
transform 1 0 58512 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1670032574
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1670032574
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1670032574
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1670032574
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1670032574
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1670032574
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1670032574
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1670032574
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1670032574
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1670032574
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1670032574
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1670032574
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1670032574
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1670032574
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1670032574
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1670032574
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1670032574
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1670032574
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_194
timestamp 1670032574
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_200
timestamp 1670032574
transform 1 0 19504 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_213
timestamp 1670032574
transform 1 0 20700 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1670032574
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1670032574
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1670032574
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1670032574
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1670032574
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1670032574
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1670032574
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1670032574
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1670032574
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1670032574
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1670032574
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1670032574
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1670032574
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1670032574
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1670032574
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1670032574
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1670032574
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1670032574
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1670032574
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1670032574
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1670032574
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1670032574
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1670032574
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1670032574
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1670032574
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1670032574
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1670032574
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1670032574
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1670032574
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1670032574
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1670032574
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1670032574
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1670032574
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1670032574
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1670032574
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1670032574
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1670032574
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1670032574
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1670032574
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_585
timestamp 1670032574
transform 1 0 54924 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_590
timestamp 1670032574
transform 1 0 55384 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_602
timestamp 1670032574
transform 1 0 56488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_610
timestamp 1670032574
transform 1 0 57224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_614
timestamp 1670032574
transform 1 0 57592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_617
timestamp 1670032574
transform 1 0 57868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_623
timestamp 1670032574
transform 1 0 58420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1670032574
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_9
timestamp 1670032574
transform 1 0 1932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_17
timestamp 1670032574
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1670032574
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1670032574
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1670032574
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1670032574
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1670032574
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1670032574
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1670032574
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1670032574
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1670032574
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1670032574
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1670032574
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1670032574
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1670032574
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1670032574
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1670032574
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1670032574
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1670032574
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1670032574
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1670032574
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1670032574
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1670032574
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1670032574
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_205
timestamp 1670032574
transform 1 0 19964 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_211
timestamp 1670032574
transform 1 0 20516 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_214
timestamp 1670032574
transform 1 0 20792 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_226
timestamp 1670032574
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_230
timestamp 1670032574
transform 1 0 22264 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_234
timestamp 1670032574
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1670032574
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1670032574
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1670032574
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1670032574
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1670032574
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1670032574
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1670032574
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1670032574
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1670032574
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1670032574
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1670032574
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1670032574
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1670032574
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1670032574
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1670032574
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1670032574
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1670032574
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1670032574
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1670032574
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1670032574
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1670032574
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1670032574
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1670032574
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1670032574
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1670032574
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1670032574
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1670032574
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1670032574
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1670032574
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1670032574
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1670032574
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1670032574
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1670032574
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1670032574
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1670032574
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1670032574
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1670032574
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1670032574
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_601
timestamp 1670032574
transform 1 0 56396 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_607
timestamp 1670032574
transform 1 0 56948 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_610
timestamp 1670032574
transform 1 0 57224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_616
timestamp 1670032574
transform 1 0 57776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_623
timestamp 1670032574
transform 1 0 58420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1670032574
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1670032574
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_19
timestamp 1670032574
transform 1 0 2852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_26
timestamp 1670032574
transform 1 0 3496 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_32
timestamp 1670032574
transform 1 0 4048 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1670032574
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1670032574
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1670032574
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1670032574
transform 1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1670032574
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1670032574
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_138
timestamp 1670032574
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_150
timestamp 1670032574
transform 1 0 14904 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1670032574
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1670032574
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1670032574
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1670032574
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_199
timestamp 1670032574
transform 1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_212
timestamp 1670032574
transform 1 0 20608 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1670032574
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1670032574
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_231
timestamp 1670032574
transform 1 0 22356 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_241
timestamp 1670032574
transform 1 0 23276 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_247
timestamp 1670032574
transform 1 0 23828 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_259
timestamp 1670032574
transform 1 0 24932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1670032574
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1670032574
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1670032574
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1670032574
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1670032574
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1670032574
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1670032574
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1670032574
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1670032574
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1670032574
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1670032574
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1670032574
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1670032574
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1670032574
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1670032574
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1670032574
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1670032574
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1670032574
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1670032574
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1670032574
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1670032574
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1670032574
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1670032574
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1670032574
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1670032574
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1670032574
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1670032574
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1670032574
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1670032574
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1670032574
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1670032574
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1670032574
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1670032574
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1670032574
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_585
timestamp 1670032574
transform 1 0 54924 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_614
timestamp 1670032574
transform 1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_617
timestamp 1670032574
transform 1 0 57868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_623
timestamp 1670032574
transform 1 0 58420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1670032574
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_18
timestamp 1670032574
transform 1 0 2760 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1670032574
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1670032574
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_33
timestamp 1670032574
transform 1 0 4140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_45
timestamp 1670032574
transform 1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1670032574
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1670032574
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1670032574
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1670032574
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1670032574
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1670032574
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1670032574
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1670032574
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1670032574
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1670032574
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_149
timestamp 1670032574
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_173
timestamp 1670032574
transform 1 0 17020 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_185
timestamp 1670032574
transform 1 0 18124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1670032574
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1670032574
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_204
timestamp 1670032574
transform 1 0 19872 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_216
timestamp 1670032574
transform 1 0 20976 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_228
timestamp 1670032574
transform 1 0 22080 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_235
timestamp 1670032574
transform 1 0 22724 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1670032574
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1670032574
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1670032574
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1670032574
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1670032574
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1670032574
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1670032574
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1670032574
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1670032574
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1670032574
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1670032574
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1670032574
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1670032574
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1670032574
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1670032574
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1670032574
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1670032574
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1670032574
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1670032574
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1670032574
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1670032574
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1670032574
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1670032574
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1670032574
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1670032574
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1670032574
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1670032574
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1670032574
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1670032574
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1670032574
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1670032574
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1670032574
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1670032574
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1670032574
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1670032574
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1670032574
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1670032574
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1670032574
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1670032574
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_601
timestamp 1670032574
transform 1 0 56396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_607
timestamp 1670032574
transform 1 0 56948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_610
timestamp 1670032574
transform 1 0 57224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_616
timestamp 1670032574
transform 1 0 57776 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_623
timestamp 1670032574
transform 1 0 58420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1670032574
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_9
timestamp 1670032574
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1670032574
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_19
timestamp 1670032574
transform 1 0 2852 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1670032574
transform 1 0 3128 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_28
timestamp 1670032574
transform 1 0 3680 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_40
timestamp 1670032574
transform 1 0 4784 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1670032574
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1670032574
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_69
timestamp 1670032574
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_75
timestamp 1670032574
transform 1 0 8004 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_97
timestamp 1670032574
transform 1 0 10028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_105
timestamp 1670032574
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1670032574
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1670032574
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_135
timestamp 1670032574
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_147
timestamp 1670032574
transform 1 0 14628 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1670032574
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1670032574
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1670032574
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1670032574
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1670032574
transform 1 0 18492 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1670032574
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_199
timestamp 1670032574
transform 1 0 19412 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_212
timestamp 1670032574
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1670032574
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_231
timestamp 1670032574
transform 1 0 22356 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_241
timestamp 1670032574
transform 1 0 23276 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_247
timestamp 1670032574
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_259
timestamp 1670032574
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_271
timestamp 1670032574
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1670032574
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1670032574
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1670032574
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1670032574
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1670032574
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1670032574
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1670032574
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1670032574
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1670032574
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1670032574
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1670032574
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1670032574
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1670032574
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1670032574
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1670032574
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1670032574
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1670032574
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1670032574
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1670032574
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1670032574
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1670032574
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1670032574
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1670032574
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1670032574
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1670032574
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1670032574
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1670032574
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1670032574
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1670032574
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1670032574
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1670032574
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1670032574
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1670032574
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1670032574
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1670032574
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_609
timestamp 1670032574
transform 1 0 57132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_614
timestamp 1670032574
transform 1 0 57592 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_617
timestamp 1670032574
transform 1 0 57868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_623
timestamp 1670032574
transform 1 0 58420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1670032574
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_9
timestamp 1670032574
transform 1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1670032574
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1670032574
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1670032574
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_55
timestamp 1670032574
transform 1 0 6164 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_67
timestamp 1670032574
transform 1 0 7268 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1670032574
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1670032574
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1670032574
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1670032574
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_109
timestamp 1670032574
transform 1 0 11132 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1670032574
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1670032574
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_153
timestamp 1670032574
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_161
timestamp 1670032574
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_184
timestamp 1670032574
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1670032574
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1670032574
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_205
timestamp 1670032574
transform 1 0 19964 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_217
timestamp 1670032574
transform 1 0 21068 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_225
timestamp 1670032574
transform 1 0 21804 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_229
timestamp 1670032574
transform 1 0 22172 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_235
timestamp 1670032574
transform 1 0 22724 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1670032574
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1670032574
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1670032574
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1670032574
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1670032574
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1670032574
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1670032574
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1670032574
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1670032574
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1670032574
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1670032574
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1670032574
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1670032574
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1670032574
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1670032574
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1670032574
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1670032574
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1670032574
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1670032574
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1670032574
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1670032574
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1670032574
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1670032574
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1670032574
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1670032574
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1670032574
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1670032574
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1670032574
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1670032574
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1670032574
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1670032574
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1670032574
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1670032574
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1670032574
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1670032574
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1670032574
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1670032574
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1670032574
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1670032574
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_601
timestamp 1670032574
transform 1 0 56396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_623
timestamp 1670032574
transform 1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1670032574
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1670032574
transform 1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_16
timestamp 1670032574
transform 1 0 2576 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_22
timestamp 1670032574
transform 1 0 3128 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_34
timestamp 1670032574
transform 1 0 4232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1670032574
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1670032574
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1670032574
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1670032574
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1670032574
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1670032574
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_105
timestamp 1670032574
transform 1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1670032574
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1670032574
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_121
timestamp 1670032574
transform 1 0 12236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1670032574
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1670032574
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1670032574
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1670032574
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1670032574
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_193
timestamp 1670032574
transform 1 0 18860 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_201
timestamp 1670032574
transform 1 0 19596 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1670032574
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1670032574
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1670032574
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1670032574
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1670032574
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_244
timestamp 1670032574
transform 1 0 23552 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_256
timestamp 1670032574
transform 1 0 24656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_268
timestamp 1670032574
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1670032574
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1670032574
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1670032574
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1670032574
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1670032574
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1670032574
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1670032574
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1670032574
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1670032574
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1670032574
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1670032574
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1670032574
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1670032574
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1670032574
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1670032574
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1670032574
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1670032574
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1670032574
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1670032574
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1670032574
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1670032574
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1670032574
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1670032574
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1670032574
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1670032574
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1670032574
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1670032574
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1670032574
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1670032574
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1670032574
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1670032574
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1670032574
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_585
timestamp 1670032574
transform 1 0 54924 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_593
timestamp 1670032574
transform 1 0 55660 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_598
timestamp 1670032574
transform 1 0 56120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_608
timestamp 1670032574
transform 1 0 57040 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_617
timestamp 1670032574
transform 1 0 57868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_623
timestamp 1670032574
transform 1 0 58420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1670032574
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_18
timestamp 1670032574
transform 1 0 2760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1670032574
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1670032574
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1670032574
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1670032574
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1670032574
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1670032574
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1670032574
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1670032574
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1670032574
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_101
timestamp 1670032574
transform 1 0 10396 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_125
timestamp 1670032574
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1670032574
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1670032574
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_153
timestamp 1670032574
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_182
timestamp 1670032574
transform 1 0 17848 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1670032574
transform 1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1670032574
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1670032574
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 1670032574
transform 1 0 19780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1670032574
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_219
timestamp 1670032574
transform 1 0 21252 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_227
timestamp 1670032574
transform 1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1670032574
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1670032574
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1670032574
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1670032574
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1670032574
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1670032574
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1670032574
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1670032574
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1670032574
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1670032574
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1670032574
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1670032574
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1670032574
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1670032574
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1670032574
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1670032574
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1670032574
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1670032574
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1670032574
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1670032574
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1670032574
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1670032574
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1670032574
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1670032574
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1670032574
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1670032574
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1670032574
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1670032574
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1670032574
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1670032574
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1670032574
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1670032574
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1670032574
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1670032574
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1670032574
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1670032574
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1670032574
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1670032574
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1670032574
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1670032574
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1670032574
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_613
timestamp 1670032574
transform 1 0 57500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_616
timestamp 1670032574
transform 1 0 57776 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_623
timestamp 1670032574
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1670032574
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_9
timestamp 1670032574
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_16
timestamp 1670032574
transform 1 0 2576 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_22
timestamp 1670032574
transform 1 0 3128 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_34
timestamp 1670032574
transform 1 0 4232 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_46
timestamp 1670032574
transform 1 0 5336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1670032574
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1670032574
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_61
timestamp 1670032574
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_65
timestamp 1670032574
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_86
timestamp 1670032574
transform 1 0 9016 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_98
timestamp 1670032574
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1670032574
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1670032574
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1670032574
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1670032574
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1670032574
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1670032574
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1670032574
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1670032574
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1670032574
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1670032574
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_199
timestamp 1670032574
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_212
timestamp 1670032574
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1670032574
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1670032574
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1670032574
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1670032574
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1670032574
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1670032574
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1670032574
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1670032574
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1670032574
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1670032574
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1670032574
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1670032574
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1670032574
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1670032574
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1670032574
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1670032574
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1670032574
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1670032574
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1670032574
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1670032574
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1670032574
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1670032574
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1670032574
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1670032574
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1670032574
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1670032574
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1670032574
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1670032574
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1670032574
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1670032574
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1670032574
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1670032574
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1670032574
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1670032574
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1670032574
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1670032574
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1670032574
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1670032574
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1670032574
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1670032574
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_609
timestamp 1670032574
transform 1 0 57132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_614
timestamp 1670032574
transform 1 0 57592 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_617
timestamp 1670032574
transform 1 0 57868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_623
timestamp 1670032574
transform 1 0 58420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1670032574
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_18
timestamp 1670032574
transform 1 0 2760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1670032574
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp 1670032574
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_55
timestamp 1670032574
transform 1 0 6164 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_67
timestamp 1670032574
transform 1 0 7268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1670032574
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1670032574
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1670032574
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1670032574
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_122
timestamp 1670032574
transform 1 0 12328 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1670032574
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1670032574
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_153
timestamp 1670032574
transform 1 0 15180 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_176
timestamp 1670032574
transform 1 0 17296 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1670032574
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1670032574
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1670032574
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1670032574
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1670032574
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1670032574
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1670032574
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1670032574
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1670032574
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1670032574
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1670032574
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1670032574
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1670032574
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1670032574
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1670032574
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1670032574
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1670032574
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1670032574
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1670032574
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1670032574
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1670032574
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1670032574
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1670032574
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1670032574
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1670032574
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1670032574
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1670032574
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1670032574
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1670032574
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1670032574
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1670032574
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1670032574
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1670032574
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1670032574
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1670032574
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1670032574
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1670032574
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1670032574
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1670032574
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1670032574
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1670032574
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1670032574
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1670032574
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1670032574
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1670032574
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_613
timestamp 1670032574
transform 1 0 57500 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_623
timestamp 1670032574
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1670032574
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_9
timestamp 1670032574
transform 1 0 1932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_17
timestamp 1670032574
transform 1 0 2668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_20
timestamp 1670032574
transform 1 0 2944 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_26
timestamp 1670032574
transform 1 0 3496 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_38
timestamp 1670032574
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1670032574
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1670032574
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1670032574
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1670032574
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1670032574
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1670032574
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1670032574
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_125
timestamp 1670032574
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1670032574
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1670032574
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1670032574
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1670032574
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1670032574
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1670032574
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1670032574
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1670032574
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1670032574
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1670032574
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1670032574
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1670032574
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1670032574
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1670032574
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1670032574
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1670032574
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1670032574
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1670032574
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1670032574
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1670032574
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1670032574
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1670032574
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1670032574
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1670032574
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1670032574
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1670032574
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1670032574
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1670032574
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1670032574
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1670032574
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1670032574
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1670032574
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1670032574
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1670032574
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1670032574
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1670032574
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1670032574
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1670032574
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1670032574
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1670032574
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1670032574
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1670032574
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1670032574
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1670032574
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1670032574
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1670032574
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1670032574
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1670032574
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1670032574
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1670032574
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1670032574
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_617
timestamp 1670032574
transform 1 0 57868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_623
timestamp 1670032574
transform 1 0 58420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1670032574
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_9
timestamp 1670032574
transform 1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1670032574
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1670032574
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp 1670032574
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_35
timestamp 1670032574
transform 1 0 4324 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_56
timestamp 1670032574
transform 1 0 6256 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_68
timestamp 1670032574
transform 1 0 7360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1670032574
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1670032574
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_107
timestamp 1670032574
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_119
timestamp 1670032574
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp 1670032574
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1670032574
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1670032574
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1670032574
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1670032574
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1670032574
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1670032574
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1670032574
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1670032574
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1670032574
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_212
timestamp 1670032574
transform 1 0 20608 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1670032574
transform 1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1670032574
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1670032574
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1670032574
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1670032574
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1670032574
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1670032574
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1670032574
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1670032574
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1670032574
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1670032574
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1670032574
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1670032574
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1670032574
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1670032574
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1670032574
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1670032574
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1670032574
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1670032574
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1670032574
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1670032574
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1670032574
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1670032574
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1670032574
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1670032574
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1670032574
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1670032574
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1670032574
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1670032574
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1670032574
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1670032574
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1670032574
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1670032574
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1670032574
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1670032574
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1670032574
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1670032574
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1670032574
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1670032574
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1670032574
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1670032574
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1670032574
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_613
timestamp 1670032574
transform 1 0 57500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_616
timestamp 1670032574
transform 1 0 57776 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_623
timestamp 1670032574
transform 1 0 58420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1670032574
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1670032574
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_16
timestamp 1670032574
transform 1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_22
timestamp 1670032574
transform 1 0 3128 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_34
timestamp 1670032574
transform 1 0 4232 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_46
timestamp 1670032574
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1670032574
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1670032574
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1670032574
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1670032574
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1670032574
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1670032574
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1670032574
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1670032574
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1670032574
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1670032574
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1670032574
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1670032574
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1670032574
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1670032574
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_193
timestamp 1670032574
transform 1 0 18860 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_201
timestamp 1670032574
transform 1 0 19596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_213
timestamp 1670032574
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1670032574
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1670032574
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1670032574
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1670032574
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1670032574
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1670032574
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1670032574
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1670032574
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1670032574
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1670032574
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1670032574
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1670032574
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1670032574
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1670032574
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1670032574
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1670032574
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1670032574
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1670032574
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1670032574
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1670032574
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1670032574
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1670032574
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1670032574
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1670032574
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1670032574
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1670032574
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1670032574
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1670032574
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1670032574
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1670032574
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1670032574
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1670032574
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1670032574
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1670032574
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1670032574
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1670032574
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1670032574
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1670032574
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1670032574
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1670032574
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1670032574
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1670032574
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1670032574
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1670032574
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1670032574
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_18
timestamp 1670032574
transform 1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1670032574
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1670032574
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1670032574
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1670032574
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1670032574
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1670032574
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1670032574
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1670032574
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1670032574
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_109
timestamp 1670032574
transform 1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_115
timestamp 1670032574
transform 1 0 11684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1670032574
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1670032574
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1670032574
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_176
timestamp 1670032574
transform 1 0 17296 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1670032574
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1670032574
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1670032574
transform 1 0 20424 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_216
timestamp 1670032574
transform 1 0 20976 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_220
timestamp 1670032574
transform 1 0 21344 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_224
timestamp 1670032574
transform 1 0 21712 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_236
timestamp 1670032574
transform 1 0 22816 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1670032574
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1670032574
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1670032574
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1670032574
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1670032574
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1670032574
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1670032574
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1670032574
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1670032574
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1670032574
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1670032574
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1670032574
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1670032574
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1670032574
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1670032574
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1670032574
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1670032574
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1670032574
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1670032574
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1670032574
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1670032574
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1670032574
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1670032574
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1670032574
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1670032574
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1670032574
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1670032574
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1670032574
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1670032574
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1670032574
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1670032574
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1670032574
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1670032574
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1670032574
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1670032574
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1670032574
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1670032574
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1670032574
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1670032574
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_613
timestamp 1670032574
transform 1 0 57500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_616
timestamp 1670032574
transform 1 0 57776 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_623
timestamp 1670032574
transform 1 0 58420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1670032574
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_18
timestamp 1670032574
transform 1 0 2760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_24
timestamp 1670032574
transform 1 0 3312 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_32
timestamp 1670032574
transform 1 0 4048 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1670032574
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1670032574
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_65
timestamp 1670032574
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_89
timestamp 1670032574
transform 1 0 9292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_101
timestamp 1670032574
transform 1 0 10396 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_107
timestamp 1670032574
transform 1 0 10948 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1670032574
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1670032574
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_123
timestamp 1670032574
transform 1 0 12420 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1670032574
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1670032574
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1670032574
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1670032574
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1670032574
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_193
timestamp 1670032574
transform 1 0 18860 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1670032574
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1670032574
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1670032574
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1670032574
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1670032574
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1670032574
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1670032574
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1670032574
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1670032574
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1670032574
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1670032574
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1670032574
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1670032574
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1670032574
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1670032574
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1670032574
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1670032574
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1670032574
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1670032574
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1670032574
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1670032574
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1670032574
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1670032574
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1670032574
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1670032574
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1670032574
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1670032574
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1670032574
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1670032574
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1670032574
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1670032574
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1670032574
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1670032574
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1670032574
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1670032574
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1670032574
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1670032574
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1670032574
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1670032574
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1670032574
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1670032574
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1670032574
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1670032574
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1670032574
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_609
timestamp 1670032574
transform 1 0 57132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_614
timestamp 1670032574
transform 1 0 57592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_617
timestamp 1670032574
transform 1 0 57868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_623
timestamp 1670032574
transform 1 0 58420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1670032574
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_9
timestamp 1670032574
transform 1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_16
timestamp 1670032574
transform 1 0 2576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1670032574
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1670032574
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1670032574
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1670032574
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1670032574
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1670032574
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1670032574
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1670032574
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_97
timestamp 1670032574
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_105
timestamp 1670032574
transform 1 0 10764 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_126
timestamp 1670032574
transform 1 0 12696 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1670032574
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1670032574
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_149
timestamp 1670032574
transform 1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_175
timestamp 1670032574
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1670032574
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1670032574
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1670032574
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1670032574
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_210
timestamp 1670032574
transform 1 0 20424 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_222
timestamp 1670032574
transform 1 0 21528 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_234
timestamp 1670032574
transform 1 0 22632 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1670032574
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1670032574
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1670032574
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1670032574
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1670032574
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1670032574
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1670032574
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1670032574
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1670032574
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1670032574
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1670032574
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1670032574
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1670032574
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1670032574
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1670032574
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1670032574
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1670032574
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1670032574
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1670032574
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1670032574
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1670032574
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1670032574
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1670032574
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1670032574
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1670032574
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1670032574
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1670032574
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1670032574
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1670032574
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1670032574
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1670032574
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1670032574
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1670032574
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1670032574
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1670032574
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1670032574
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1670032574
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1670032574
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1670032574
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_613
timestamp 1670032574
transform 1 0 57500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_623
timestamp 1670032574
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1670032574
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_9
timestamp 1670032574
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_21
timestamp 1670032574
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_33
timestamp 1670032574
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1670032574
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1670032574
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_69
timestamp 1670032574
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1670032574
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1670032574
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1670032574
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_125
timestamp 1670032574
transform 1 0 12604 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_148
timestamp 1670032574
transform 1 0 14720 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1670032574
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1670032574
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1670032574
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1670032574
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1670032574
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1670032574
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1670032574
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1670032574
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1670032574
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1670032574
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1670032574
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1670032574
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1670032574
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1670032574
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1670032574
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1670032574
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1670032574
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1670032574
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1670032574
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1670032574
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1670032574
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1670032574
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1670032574
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1670032574
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1670032574
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1670032574
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1670032574
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1670032574
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1670032574
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1670032574
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1670032574
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1670032574
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1670032574
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1670032574
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1670032574
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1670032574
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1670032574
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1670032574
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1670032574
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1670032574
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1670032574
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1670032574
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1670032574
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1670032574
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1670032574
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1670032574
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_597
timestamp 1670032574
transform 1 0 56028 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_603
timestamp 1670032574
transform 1 0 56580 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_614
timestamp 1670032574
transform 1 0 57592 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_617
timestamp 1670032574
transform 1 0 57868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_623
timestamp 1670032574
transform 1 0 58420 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1670032574
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_9
timestamp 1670032574
transform 1 0 1932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1670032574
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1670032574
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1670032574
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_41
timestamp 1670032574
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1670032574
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_59
timestamp 1670032574
transform 1 0 6532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_71
timestamp 1670032574
transform 1 0 7636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1670032574
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1670032574
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1670032574
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1670032574
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1670032574
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1670032574
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1670032574
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1670032574
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1670032574
transform 1 0 15180 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_175
timestamp 1670032574
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1670032574
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_191
timestamp 1670032574
transform 1 0 18676 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1670032574
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1670032574
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_201
timestamp 1670032574
transform 1 0 19596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_213
timestamp 1670032574
transform 1 0 20700 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_225
timestamp 1670032574
transform 1 0 21804 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_237
timestamp 1670032574
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1670032574
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1670032574
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1670032574
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1670032574
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1670032574
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1670032574
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1670032574
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1670032574
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1670032574
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1670032574
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1670032574
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1670032574
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1670032574
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1670032574
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1670032574
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1670032574
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1670032574
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1670032574
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1670032574
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1670032574
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1670032574
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1670032574
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1670032574
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1670032574
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1670032574
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1670032574
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1670032574
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1670032574
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1670032574
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1670032574
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1670032574
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1670032574
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1670032574
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1670032574
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1670032574
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1670032574
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1670032574
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1670032574
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1670032574
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_613
timestamp 1670032574
transform 1 0 57500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_616
timestamp 1670032574
transform 1 0 57776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_623
timestamp 1670032574
transform 1 0 58420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1670032574
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_9
timestamp 1670032574
transform 1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_16
timestamp 1670032574
transform 1 0 2576 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_28
timestamp 1670032574
transform 1 0 3680 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1670032574
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1670032574
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1670032574
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_81
timestamp 1670032574
transform 1 0 8556 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1670032574
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1670032574
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1670032574
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1670032574
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1670032574
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1670032574
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1670032574
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1670032574
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1670032574
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1670032574
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1670032574
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_211
timestamp 1670032574
transform 1 0 20516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1670032574
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1670032574
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1670032574
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1670032574
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1670032574
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1670032574
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1670032574
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1670032574
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1670032574
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1670032574
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1670032574
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1670032574
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1670032574
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1670032574
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1670032574
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1670032574
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1670032574
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1670032574
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1670032574
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1670032574
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1670032574
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1670032574
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1670032574
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1670032574
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1670032574
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1670032574
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1670032574
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1670032574
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1670032574
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1670032574
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1670032574
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1670032574
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1670032574
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1670032574
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1670032574
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1670032574
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1670032574
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1670032574
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1670032574
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1670032574
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1670032574
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1670032574
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1670032574
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1670032574
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1670032574
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_18
timestamp 1670032574
transform 1 0 2760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1670032574
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1670032574
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1670032574
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1670032574
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1670032574
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1670032574
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1670032574
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1670032574
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1670032574
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1670032574
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_117
timestamp 1670032574
transform 1 0 11868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1670032574
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1670032574
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_153
timestamp 1670032574
transform 1 0 15180 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_174
timestamp 1670032574
transform 1 0 17112 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_188
timestamp 1670032574
transform 1 0 18400 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1670032574
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1670032574
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1670032574
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_214
timestamp 1670032574
transform 1 0 20792 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_226
timestamp 1670032574
transform 1 0 21896 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_238
timestamp 1670032574
transform 1 0 23000 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1670032574
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1670032574
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1670032574
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1670032574
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1670032574
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1670032574
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1670032574
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1670032574
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1670032574
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1670032574
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1670032574
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1670032574
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1670032574
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1670032574
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1670032574
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1670032574
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1670032574
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1670032574
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1670032574
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1670032574
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1670032574
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1670032574
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1670032574
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1670032574
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1670032574
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1670032574
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1670032574
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1670032574
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1670032574
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1670032574
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1670032574
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1670032574
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1670032574
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1670032574
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1670032574
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1670032574
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1670032574
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1670032574
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1670032574
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_613
timestamp 1670032574
transform 1 0 57500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_616
timestamp 1670032574
transform 1 0 57776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_623
timestamp 1670032574
transform 1 0 58420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1670032574
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_9
timestamp 1670032574
transform 1 0 1932 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_17
timestamp 1670032574
transform 1 0 2668 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_20
timestamp 1670032574
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_32
timestamp 1670032574
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_44
timestamp 1670032574
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1670032574
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1670032574
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1670032574
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1670032574
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1670032574
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1670032574
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1670032574
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1670032574
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_158
timestamp 1670032574
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1670032574
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1670032574
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1670032574
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_193
timestamp 1670032574
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1670032574
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_208
timestamp 1670032574
transform 1 0 20240 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1670032574
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1670032574
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1670032574
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1670032574
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1670032574
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1670032574
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1670032574
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1670032574
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1670032574
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1670032574
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1670032574
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1670032574
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1670032574
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1670032574
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1670032574
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1670032574
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1670032574
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1670032574
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1670032574
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1670032574
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1670032574
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1670032574
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1670032574
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1670032574
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1670032574
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1670032574
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1670032574
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1670032574
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1670032574
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1670032574
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1670032574
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1670032574
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1670032574
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1670032574
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1670032574
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1670032574
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1670032574
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1670032574
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1670032574
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1670032574
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1670032574
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_609
timestamp 1670032574
transform 1 0 57132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_614
timestamp 1670032574
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_617
timestamp 1670032574
transform 1 0 57868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1670032574
transform 1 0 58420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1670032574
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_9
timestamp 1670032574
transform 1 0 1932 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_17
timestamp 1670032574
transform 1 0 2668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1670032574
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1670032574
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_37
timestamp 1670032574
transform 1 0 4508 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_60
timestamp 1670032574
transform 1 0 6624 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_72
timestamp 1670032574
transform 1 0 7728 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1670032574
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1670032574
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1670032574
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1670032574
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1670032574
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1670032574
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1670032574
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1670032574
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_172
timestamp 1670032574
transform 1 0 16928 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_184
timestamp 1670032574
transform 1 0 18032 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1670032574
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1670032574
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1670032574
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1670032574
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1670032574
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1670032574
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1670032574
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1670032574
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1670032574
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1670032574
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1670032574
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1670032574
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1670032574
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1670032574
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1670032574
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1670032574
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1670032574
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1670032574
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1670032574
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1670032574
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1670032574
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1670032574
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1670032574
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1670032574
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1670032574
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1670032574
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1670032574
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1670032574
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1670032574
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1670032574
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1670032574
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1670032574
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1670032574
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1670032574
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1670032574
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1670032574
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1670032574
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1670032574
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1670032574
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1670032574
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1670032574
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1670032574
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1670032574
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1670032574
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1670032574
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_613
timestamp 1670032574
transform 1 0 57500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_616
timestamp 1670032574
transform 1 0 57776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_623
timestamp 1670032574
transform 1 0 58420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1670032574
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_18
timestamp 1670032574
transform 1 0 2760 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_24
timestamp 1670032574
transform 1 0 3312 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_36
timestamp 1670032574
transform 1 0 4416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1670032574
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1670032574
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1670032574
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_77
timestamp 1670032574
transform 1 0 8188 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_99
timestamp 1670032574
transform 1 0 10212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1670032574
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1670032574
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_121
timestamp 1670032574
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_144
timestamp 1670032574
transform 1 0 14352 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_156
timestamp 1670032574
transform 1 0 15456 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1670032574
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1670032574
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_188
timestamp 1670032574
transform 1 0 18400 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_201
timestamp 1670032574
transform 1 0 19596 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_207
timestamp 1670032574
transform 1 0 20148 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1670032574
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1670032574
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1670032574
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1670032574
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1670032574
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1670032574
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1670032574
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1670032574
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1670032574
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1670032574
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1670032574
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1670032574
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1670032574
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1670032574
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1670032574
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1670032574
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1670032574
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1670032574
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1670032574
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1670032574
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1670032574
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1670032574
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1670032574
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1670032574
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1670032574
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1670032574
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1670032574
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1670032574
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1670032574
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1670032574
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1670032574
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1670032574
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1670032574
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1670032574
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1670032574
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1670032574
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1670032574
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1670032574
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1670032574
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1670032574
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1670032574
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1670032574
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_609
timestamp 1670032574
transform 1 0 57132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_614
timestamp 1670032574
transform 1 0 57592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_617
timestamp 1670032574
transform 1 0 57868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1670032574
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1670032574
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_9
timestamp 1670032574
transform 1 0 1932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_16
timestamp 1670032574
transform 1 0 2576 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1670032574
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1670032574
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1670032574
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_33
timestamp 1670032574
transform 1 0 4140 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_61
timestamp 1670032574
transform 1 0 6716 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_73
timestamp 1670032574
transform 1 0 7820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_81
timestamp 1670032574
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1670032574
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_97
timestamp 1670032574
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_124
timestamp 1670032574
transform 1 0 12512 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1670032574
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1670032574
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1670032574
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1670032574
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_177
timestamp 1670032574
transform 1 0 17388 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_185
timestamp 1670032574
transform 1 0 18124 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1670032574
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1670032574
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1670032574
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1670032574
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1670032574
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1670032574
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1670032574
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1670032574
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1670032574
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1670032574
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1670032574
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1670032574
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1670032574
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1670032574
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1670032574
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1670032574
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1670032574
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1670032574
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1670032574
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1670032574
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1670032574
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1670032574
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1670032574
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1670032574
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1670032574
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1670032574
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1670032574
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1670032574
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1670032574
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1670032574
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1670032574
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1670032574
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1670032574
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1670032574
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1670032574
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1670032574
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1670032574
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1670032574
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1670032574
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1670032574
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1670032574
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1670032574
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1670032574
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1670032574
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_601
timestamp 1670032574
transform 1 0 56396 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_609
timestamp 1670032574
transform 1 0 57132 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_620
timestamp 1670032574
transform 1 0 58144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_624
timestamp 1670032574
transform 1 0 58512 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1670032574
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_18
timestamp 1670032574
transform 1 0 2760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_24
timestamp 1670032574
transform 1 0 3312 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1670032574
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1670032574
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1670032574
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1670032574
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_94
timestamp 1670032574
transform 1 0 9752 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_106
timestamp 1670032574
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1670032574
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1670032574
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1670032574
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1670032574
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1670032574
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1670032574
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1670032574
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1670032574
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1670032574
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1670032574
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1670032574
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1670032574
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1670032574
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1670032574
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1670032574
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1670032574
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1670032574
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1670032574
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1670032574
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1670032574
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1670032574
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1670032574
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1670032574
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1670032574
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1670032574
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1670032574
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1670032574
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1670032574
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1670032574
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1670032574
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1670032574
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1670032574
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1670032574
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1670032574
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1670032574
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1670032574
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1670032574
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1670032574
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1670032574
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1670032574
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1670032574
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1670032574
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1670032574
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1670032574
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1670032574
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1670032574
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1670032574
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1670032574
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1670032574
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1670032574
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1670032574
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1670032574
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1670032574
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1670032574
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_617
timestamp 1670032574
transform 1 0 57868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_623
timestamp 1670032574
transform 1 0 58420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1670032574
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_9
timestamp 1670032574
transform 1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_15
timestamp 1670032574
transform 1 0 2484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1670032574
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1670032574
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1670032574
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1670032574
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1670032574
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1670032574
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1670032574
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1670032574
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1670032574
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1670032574
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1670032574
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1670032574
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1670032574
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1670032574
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1670032574
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1670032574
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1670032574
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1670032574
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1670032574
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1670032574
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1670032574
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1670032574
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_211
timestamp 1670032574
transform 1 0 20516 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_223
timestamp 1670032574
transform 1 0 21620 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_235
timestamp 1670032574
transform 1 0 22724 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1670032574
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1670032574
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1670032574
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1670032574
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1670032574
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1670032574
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1670032574
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1670032574
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1670032574
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1670032574
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1670032574
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1670032574
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1670032574
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1670032574
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1670032574
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1670032574
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1670032574
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1670032574
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1670032574
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1670032574
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1670032574
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1670032574
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1670032574
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1670032574
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1670032574
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1670032574
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1670032574
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1670032574
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1670032574
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1670032574
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1670032574
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1670032574
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1670032574
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1670032574
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1670032574
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1670032574
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1670032574
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1670032574
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1670032574
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_601
timestamp 1670032574
transform 1 0 56396 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_607
timestamp 1670032574
transform 1 0 56948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_610
timestamp 1670032574
transform 1 0 57224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_616
timestamp 1670032574
transform 1 0 57776 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_623
timestamp 1670032574
transform 1 0 58420 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1670032574
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_9
timestamp 1670032574
transform 1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp 1670032574
transform 1 0 2484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_21
timestamp 1670032574
transform 1 0 3036 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1670032574
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1670032574
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1670032574
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1670032574
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1670032574
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1670032574
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1670032574
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1670032574
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1670032574
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1670032574
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1670032574
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1670032574
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1670032574
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1670032574
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1670032574
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1670032574
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1670032574
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1670032574
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1670032574
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1670032574
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1670032574
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1670032574
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1670032574
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1670032574
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1670032574
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1670032574
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1670032574
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1670032574
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1670032574
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1670032574
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1670032574
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1670032574
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1670032574
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1670032574
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1670032574
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1670032574
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1670032574
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1670032574
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1670032574
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1670032574
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1670032574
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1670032574
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1670032574
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1670032574
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1670032574
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1670032574
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1670032574
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1670032574
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1670032574
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1670032574
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1670032574
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1670032574
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1670032574
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1670032574
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1670032574
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1670032574
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1670032574
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1670032574
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1670032574
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1670032574
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1670032574
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_597
timestamp 1670032574
transform 1 0 56028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_605
timestamp 1670032574
transform 1 0 56764 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_608
timestamp 1670032574
transform 1 0 57040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_614
timestamp 1670032574
transform 1 0 57592 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_617
timestamp 1670032574
transform 1 0 57868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1670032574
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1670032574
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_9
timestamp 1670032574
transform 1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_13
timestamp 1670032574
transform 1 0 2300 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_17
timestamp 1670032574
transform 1 0 2668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1670032574
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1670032574
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1670032574
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1670032574
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1670032574
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_65
timestamp 1670032574
transform 1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_70
timestamp 1670032574
transform 1 0 7544 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_78
timestamp 1670032574
transform 1 0 8280 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1670032574
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1670032574
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_90
timestamp 1670032574
transform 1 0 9384 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_102
timestamp 1670032574
transform 1 0 10488 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_108
timestamp 1670032574
transform 1 0 11040 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_111
timestamp 1670032574
transform 1 0 11316 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_117
timestamp 1670032574
transform 1 0 11868 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp 1670032574
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1670032574
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1670032574
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_147
timestamp 1670032574
transform 1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1670032574
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_159
timestamp 1670032574
transform 1 0 15732 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_167
timestamp 1670032574
transform 1 0 16468 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_172
timestamp 1670032574
transform 1 0 16928 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_184
timestamp 1670032574
transform 1 0 18032 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1670032574
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1670032574
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1670032574
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1670032574
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1670032574
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1670032574
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1670032574
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1670032574
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1670032574
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1670032574
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1670032574
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1670032574
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1670032574
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1670032574
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1670032574
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1670032574
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1670032574
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1670032574
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1670032574
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1670032574
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1670032574
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1670032574
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1670032574
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1670032574
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1670032574
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1670032574
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1670032574
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1670032574
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1670032574
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1670032574
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1670032574
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1670032574
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1670032574
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1670032574
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1670032574
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1670032574
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1670032574
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1670032574
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1670032574
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1670032574
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1670032574
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1670032574
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1670032574
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_601
timestamp 1670032574
transform 1 0 56396 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_623
timestamp 1670032574
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_3
timestamp 1670032574
transform 1 0 1380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_9
timestamp 1670032574
transform 1 0 1932 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_19
timestamp 1670032574
transform 1 0 2852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_27
timestamp 1670032574
transform 1 0 3588 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_31
timestamp 1670032574
transform 1 0 3956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_39
timestamp 1670032574
transform 1 0 4692 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_42
timestamp 1670032574
transform 1 0 4968 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1670032574
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_57
timestamp 1670032574
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_62
timestamp 1670032574
transform 1 0 6808 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1670032574
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_82
timestamp 1670032574
transform 1 0 8648 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_90
timestamp 1670032574
transform 1 0 9384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_94
timestamp 1670032574
transform 1 0 9752 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 1670032574
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1670032574
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1670032574
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_117
timestamp 1670032574
transform 1 0 11868 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_129
timestamp 1670032574
transform 1 0 12972 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_134
timestamp 1670032574
transform 1 0 13432 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_147
timestamp 1670032574
transform 1 0 14628 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_153
timestamp 1670032574
transform 1 0 15180 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_156
timestamp 1670032574
transform 1 0 15456 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_163
timestamp 1670032574
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1670032574
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1670032574
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_174
timestamp 1670032574
transform 1 0 17112 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_180
timestamp 1670032574
transform 1 0 17664 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_192
timestamp 1670032574
transform 1 0 18768 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_204
timestamp 1670032574
transform 1 0 19872 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1670032574
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1670032574
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1670032574
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1670032574
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1670032574
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1670032574
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1670032574
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1670032574
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1670032574
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1670032574
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1670032574
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1670032574
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1670032574
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1670032574
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1670032574
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1670032574
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1670032574
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1670032574
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1670032574
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1670032574
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1670032574
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1670032574
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1670032574
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1670032574
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1670032574
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1670032574
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1670032574
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1670032574
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1670032574
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1670032574
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1670032574
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1670032574
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1670032574
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1670032574
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1670032574
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1670032574
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1670032574
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1670032574
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1670032574
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1670032574
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_597
timestamp 1670032574
transform 1 0 56028 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_601
timestamp 1670032574
transform 1 0 56396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_607
timestamp 1670032574
transform 1 0 56948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_614
timestamp 1670032574
transform 1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_617
timestamp 1670032574
transform 1 0 57868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1670032574
transform 1 0 58420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1670032574
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_9
timestamp 1670032574
transform 1 0 1932 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1670032574
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1670032574
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_40
timestamp 1670032574
transform 1 0 4784 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_46
timestamp 1670032574
transform 1 0 5336 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_53
timestamp 1670032574
transform 1 0 5980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_66
timestamp 1670032574
transform 1 0 7176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_72
timestamp 1670032574
transform 1 0 7728 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1670032574
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1670032574
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_89
timestamp 1670032574
transform 1 0 9292 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_99
timestamp 1670032574
transform 1 0 10212 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_107
timestamp 1670032574
transform 1 0 10948 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_112
timestamp 1670032574
transform 1 0 11408 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_116
timestamp 1670032574
transform 1 0 11776 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_120
timestamp 1670032574
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1670032574
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_132
timestamp 1670032574
transform 1 0 13248 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1670032574
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1670032574
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_147
timestamp 1670032574
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_157
timestamp 1670032574
transform 1 0 15548 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_170
timestamp 1670032574
transform 1 0 16744 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_183
timestamp 1670032574
transform 1 0 17940 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1670032574
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1670032574
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1670032574
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1670032574
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1670032574
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1670032574
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1670032574
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1670032574
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1670032574
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1670032574
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1670032574
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1670032574
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1670032574
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1670032574
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1670032574
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1670032574
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1670032574
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1670032574
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1670032574
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1670032574
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1670032574
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1670032574
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1670032574
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1670032574
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1670032574
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1670032574
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1670032574
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1670032574
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1670032574
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1670032574
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_469
timestamp 1670032574
transform 1 0 44252 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_473
timestamp 1670032574
transform 1 0 44620 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1670032574
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1670032574
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1670032574
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1670032574
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1670032574
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1670032574
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1670032574
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1670032574
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1670032574
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1670032574
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1670032574
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1670032574
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1670032574
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_601
timestamp 1670032574
transform 1 0 56396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_623
timestamp 1670032574
transform 1 0 58420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1670032574
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_11
timestamp 1670032574
transform 1 0 2116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_23
timestamp 1670032574
transform 1 0 3220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_27
timestamp 1670032574
transform 1 0 3588 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_30
timestamp 1670032574
transform 1 0 3864 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_36
timestamp 1670032574
transform 1 0 4416 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_44
timestamp 1670032574
transform 1 0 5152 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_48
timestamp 1670032574
transform 1 0 5520 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1670032574
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1670032574
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_62
timestamp 1670032574
transform 1 0 6808 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_68
timestamp 1670032574
transform 1 0 7360 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_76
timestamp 1670032574
transform 1 0 8096 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_80
timestamp 1670032574
transform 1 0 8464 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_93
timestamp 1670032574
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1670032574
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1670032574
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_118
timestamp 1670032574
transform 1 0 11960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 1670032574
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_138
timestamp 1670032574
transform 1 0 13800 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_149
timestamp 1670032574
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_155
timestamp 1670032574
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1670032574
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1670032574
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1670032574
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_174
timestamp 1670032574
transform 1 0 17112 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_180
timestamp 1670032574
transform 1 0 17664 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_192
timestamp 1670032574
transform 1 0 18768 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_204
timestamp 1670032574
transform 1 0 19872 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1670032574
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1670032574
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1670032574
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1670032574
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1670032574
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1670032574
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1670032574
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1670032574
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1670032574
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1670032574
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1670032574
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1670032574
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1670032574
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1670032574
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1670032574
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1670032574
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1670032574
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1670032574
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1670032574
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1670032574
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1670032574
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1670032574
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1670032574
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1670032574
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1670032574
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1670032574
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1670032574
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1670032574
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1670032574
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1670032574
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1670032574
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1670032574
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1670032574
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1670032574
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1670032574
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1670032574
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1670032574
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1670032574
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1670032574
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1670032574
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_597
timestamp 1670032574
transform 1 0 56028 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_605
timestamp 1670032574
transform 1 0 56764 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_608
timestamp 1670032574
transform 1 0 57040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_614
timestamp 1670032574
transform 1 0 57592 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_617
timestamp 1670032574
transform 1 0 57868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_623
timestamp 1670032574
transform 1 0 58420 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1670032574
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_9
timestamp 1670032574
transform 1 0 1932 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1670032574
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1670032574
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1670032574
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_41
timestamp 1670032574
transform 1 0 4876 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_51
timestamp 1670032574
transform 1 0 5796 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_64
timestamp 1670032574
transform 1 0 6992 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_71
timestamp 1670032574
transform 1 0 7636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1670032574
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1670032574
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1670032574
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_93
timestamp 1670032574
transform 1 0 9660 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1670032574
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_103
timestamp 1670032574
transform 1 0 10580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_111
timestamp 1670032574
transform 1 0 11316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_116
timestamp 1670032574
transform 1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_122
timestamp 1670032574
transform 1 0 12328 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1670032574
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1670032574
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_145
timestamp 1670032574
transform 1 0 14444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_151
timestamp 1670032574
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_157
timestamp 1670032574
transform 1 0 15548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_169
timestamp 1670032574
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_181
timestamp 1670032574
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1670032574
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1670032574
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1670032574
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1670032574
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1670032574
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1670032574
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1670032574
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1670032574
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1670032574
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1670032574
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1670032574
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1670032574
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1670032574
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1670032574
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1670032574
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1670032574
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1670032574
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1670032574
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1670032574
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1670032574
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1670032574
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1670032574
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1670032574
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1670032574
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1670032574
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1670032574
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1670032574
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1670032574
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1670032574
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1670032574
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1670032574
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1670032574
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1670032574
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1670032574
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1670032574
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1670032574
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1670032574
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1670032574
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1670032574
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1670032574
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1670032574
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1670032574
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1670032574
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1670032574
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_601
timestamp 1670032574
transform 1 0 56396 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_607
timestamp 1670032574
transform 1 0 56948 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_610
timestamp 1670032574
transform 1 0 57224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_616
timestamp 1670032574
transform 1 0 57776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_623
timestamp 1670032574
transform 1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1670032574
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_9
timestamp 1670032574
transform 1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1670032574
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1670032574
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1670032574
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_51
timestamp 1670032574
transform 1 0 5796 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1670032574
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_57
timestamp 1670032574
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_63
timestamp 1670032574
transform 1 0 6900 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_66
timestamp 1670032574
transform 1 0 7176 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_78
timestamp 1670032574
transform 1 0 8280 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_90
timestamp 1670032574
transform 1 0 9384 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_96
timestamp 1670032574
transform 1 0 9936 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_103
timestamp 1670032574
transform 1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1670032574
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1670032574
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1670032574
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_137
timestamp 1670032574
transform 1 0 13708 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1670032574
transform 1 0 13984 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_146
timestamp 1670032574
transform 1 0 14536 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_154
timestamp 1670032574
transform 1 0 15272 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_158
timestamp 1670032574
transform 1 0 15640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1670032574
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1670032574
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1670032574
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1670032574
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1670032574
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1670032574
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1670032574
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1670032574
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1670032574
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1670032574
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1670032574
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1670032574
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1670032574
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1670032574
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1670032574
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1670032574
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1670032574
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1670032574
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1670032574
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1670032574
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1670032574
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1670032574
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1670032574
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1670032574
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1670032574
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1670032574
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1670032574
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1670032574
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1670032574
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1670032574
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1670032574
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1670032574
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1670032574
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1670032574
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1670032574
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1670032574
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1670032574
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1670032574
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1670032574
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1670032574
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1670032574
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1670032574
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1670032574
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1670032574
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1670032574
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1670032574
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1670032574
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_609
timestamp 1670032574
transform 1 0 57132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_614
timestamp 1670032574
transform 1 0 57592 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_617
timestamp 1670032574
transform 1 0 57868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_623
timestamp 1670032574
transform 1 0 58420 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1670032574
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1670032574
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1670032574
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1670032574
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1670032574
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_53
timestamp 1670032574
transform 1 0 5980 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_62
timestamp 1670032574
transform 1 0 6808 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_70
timestamp 1670032574
transform 1 0 7544 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1670032574
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1670032574
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1670032574
transform 1 0 9660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_104
timestamp 1670032574
transform 1 0 10672 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_110
timestamp 1670032574
transform 1 0 11224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_116
timestamp 1670032574
transform 1 0 11776 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_122
timestamp 1670032574
transform 1 0 12328 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_125
timestamp 1670032574
transform 1 0 12604 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1670032574
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1670032574
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_145
timestamp 1670032574
transform 1 0 14444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_157
timestamp 1670032574
transform 1 0 15548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_169
timestamp 1670032574
transform 1 0 16652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_181
timestamp 1670032574
transform 1 0 17756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1670032574
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1670032574
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1670032574
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1670032574
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1670032574
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1670032574
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1670032574
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1670032574
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1670032574
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1670032574
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1670032574
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1670032574
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1670032574
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1670032574
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1670032574
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1670032574
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1670032574
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1670032574
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1670032574
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1670032574
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1670032574
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1670032574
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1670032574
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1670032574
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1670032574
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1670032574
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1670032574
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1670032574
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1670032574
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1670032574
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1670032574
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1670032574
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1670032574
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1670032574
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1670032574
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1670032574
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1670032574
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1670032574
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1670032574
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1670032574
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1670032574
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1670032574
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1670032574
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1670032574
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_601
timestamp 1670032574
transform 1 0 56396 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_607
timestamp 1670032574
transform 1 0 56948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_610
timestamp 1670032574
transform 1 0 57224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_616
timestamp 1670032574
transform 1 0 57776 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_623
timestamp 1670032574
transform 1 0 58420 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1670032574
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_9
timestamp 1670032574
transform 1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1670032574
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1670032574
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1670032574
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1670032574
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1670032574
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1670032574
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_68
timestamp 1670032574
transform 1 0 7360 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_74
timestamp 1670032574
transform 1 0 7912 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_80
timestamp 1670032574
transform 1 0 8464 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_84
timestamp 1670032574
transform 1 0 8832 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_94
timestamp 1670032574
transform 1 0 9752 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_100
timestamp 1670032574
transform 1 0 10304 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_106
timestamp 1670032574
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1670032574
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1670032574
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1670032574
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1670032574
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1670032574
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1670032574
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1670032574
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1670032574
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1670032574
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1670032574
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1670032574
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1670032574
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1670032574
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1670032574
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1670032574
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1670032574
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1670032574
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1670032574
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1670032574
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1670032574
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1670032574
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1670032574
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1670032574
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1670032574
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1670032574
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1670032574
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1670032574
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1670032574
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1670032574
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1670032574
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1670032574
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1670032574
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1670032574
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1670032574
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1670032574
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1670032574
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1670032574
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1670032574
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1670032574
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1670032574
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1670032574
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1670032574
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1670032574
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1670032574
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1670032574
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1670032574
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1670032574
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1670032574
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1670032574
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1670032574
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1670032574
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_597
timestamp 1670032574
transform 1 0 56028 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_605
timestamp 1670032574
transform 1 0 56764 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_608
timestamp 1670032574
transform 1 0 57040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_614
timestamp 1670032574
transform 1 0 57592 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_617
timestamp 1670032574
transform 1 0 57868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_623
timestamp 1670032574
transform 1 0 58420 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1670032574
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_9
timestamp 1670032574
transform 1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1670032574
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1670032574
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1670032574
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1670032574
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1670032574
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1670032574
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1670032574
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1670032574
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1670032574
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_93
timestamp 1670032574
transform 1 0 9660 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_98
timestamp 1670032574
transform 1 0 10120 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_104
timestamp 1670032574
transform 1 0 10672 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_116
timestamp 1670032574
transform 1 0 11776 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_128
timestamp 1670032574
transform 1 0 12880 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1670032574
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1670032574
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1670032574
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1670032574
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1670032574
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1670032574
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1670032574
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1670032574
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1670032574
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1670032574
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1670032574
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1670032574
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1670032574
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1670032574
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1670032574
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1670032574
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1670032574
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1670032574
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1670032574
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1670032574
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1670032574
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1670032574
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1670032574
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1670032574
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1670032574
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1670032574
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1670032574
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1670032574
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1670032574
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1670032574
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1670032574
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1670032574
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1670032574
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1670032574
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1670032574
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1670032574
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1670032574
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1670032574
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1670032574
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1670032574
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1670032574
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1670032574
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1670032574
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1670032574
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1670032574
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1670032574
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1670032574
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1670032574
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1670032574
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_622
timestamp 1670032574
transform 1 0 58328 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1670032574
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1670032574
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1670032574
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1670032574
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1670032574
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1670032574
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1670032574
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1670032574
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1670032574
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1670032574
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1670032574
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1670032574
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1670032574
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1670032574
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1670032574
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1670032574
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1670032574
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1670032574
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1670032574
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1670032574
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1670032574
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1670032574
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1670032574
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1670032574
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1670032574
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1670032574
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1670032574
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1670032574
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1670032574
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1670032574
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1670032574
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1670032574
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1670032574
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1670032574
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1670032574
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1670032574
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1670032574
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1670032574
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1670032574
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1670032574
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1670032574
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1670032574
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1670032574
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1670032574
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1670032574
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1670032574
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1670032574
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1670032574
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1670032574
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1670032574
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1670032574
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1670032574
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1670032574
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1670032574
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1670032574
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1670032574
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1670032574
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1670032574
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1670032574
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1670032574
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1670032574
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1670032574
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1670032574
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_597
timestamp 1670032574
transform 1 0 56028 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_602
timestamp 1670032574
transform 1 0 56488 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_608
timestamp 1670032574
transform 1 0 57040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_614
timestamp 1670032574
transform 1 0 57592 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_617
timestamp 1670032574
transform 1 0 57868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_623
timestamp 1670032574
transform 1 0 58420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1670032574
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1670032574
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1670032574
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1670032574
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1670032574
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1670032574
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1670032574
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1670032574
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1670032574
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1670032574
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1670032574
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1670032574
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1670032574
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1670032574
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1670032574
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1670032574
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1670032574
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1670032574
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1670032574
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1670032574
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1670032574
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1670032574
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1670032574
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1670032574
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1670032574
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1670032574
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1670032574
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1670032574
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1670032574
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1670032574
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1670032574
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1670032574
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1670032574
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1670032574
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1670032574
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1670032574
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1670032574
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1670032574
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1670032574
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1670032574
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1670032574
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1670032574
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1670032574
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1670032574
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1670032574
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1670032574
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1670032574
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1670032574
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1670032574
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1670032574
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1670032574
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1670032574
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1670032574
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1670032574
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1670032574
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1670032574
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1670032574
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1670032574
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1670032574
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1670032574
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1670032574
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1670032574
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1670032574
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1670032574
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1670032574
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_601
timestamp 1670032574
transform 1 0 56396 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_620
timestamp 1670032574
transform 1 0 58144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_624
timestamp 1670032574
transform 1 0 58512 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1670032574
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_9
timestamp 1670032574
transform 1 0 1932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1670032574
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1670032574
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1670032574
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1670032574
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1670032574
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1670032574
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1670032574
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1670032574
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1670032574
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1670032574
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1670032574
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1670032574
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1670032574
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1670032574
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1670032574
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1670032574
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1670032574
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1670032574
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1670032574
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1670032574
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1670032574
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1670032574
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1670032574
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1670032574
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1670032574
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1670032574
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1670032574
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1670032574
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1670032574
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1670032574
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1670032574
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1670032574
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1670032574
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1670032574
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1670032574
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1670032574
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1670032574
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1670032574
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1670032574
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1670032574
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1670032574
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1670032574
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1670032574
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1670032574
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1670032574
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1670032574
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1670032574
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1670032574
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1670032574
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1670032574
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1670032574
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1670032574
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1670032574
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1670032574
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1670032574
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1670032574
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1670032574
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1670032574
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1670032574
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1670032574
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1670032574
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_597
timestamp 1670032574
transform 1 0 56028 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_605
timestamp 1670032574
transform 1 0 56764 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_608
timestamp 1670032574
transform 1 0 57040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_614
timestamp 1670032574
transform 1 0 57592 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_617
timestamp 1670032574
transform 1 0 57868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1670032574
transform 1 0 58420 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1670032574
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1670032574
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1670032574
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1670032574
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1670032574
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1670032574
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1670032574
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1670032574
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1670032574
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1670032574
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1670032574
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1670032574
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1670032574
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1670032574
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1670032574
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1670032574
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1670032574
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1670032574
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1670032574
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1670032574
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1670032574
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1670032574
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1670032574
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1670032574
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1670032574
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1670032574
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1670032574
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1670032574
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1670032574
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1670032574
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1670032574
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1670032574
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1670032574
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1670032574
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1670032574
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1670032574
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1670032574
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1670032574
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1670032574
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1670032574
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1670032574
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1670032574
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1670032574
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1670032574
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1670032574
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1670032574
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1670032574
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1670032574
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1670032574
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1670032574
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1670032574
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1670032574
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1670032574
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1670032574
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1670032574
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1670032574
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1670032574
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1670032574
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1670032574
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1670032574
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1670032574
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1670032574
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1670032574
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_589
timestamp 1670032574
transform 1 0 55292 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_594
timestamp 1670032574
transform 1 0 55752 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_606
timestamp 1670032574
transform 1 0 56856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_616
timestamp 1670032574
transform 1 0 57776 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_620
timestamp 1670032574
transform 1 0 58144 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_623
timestamp 1670032574
transform 1 0 58420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1670032574
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1670032574
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1670032574
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1670032574
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1670032574
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1670032574
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1670032574
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1670032574
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1670032574
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1670032574
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1670032574
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1670032574
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1670032574
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1670032574
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1670032574
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1670032574
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1670032574
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1670032574
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1670032574
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1670032574
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1670032574
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1670032574
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1670032574
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1670032574
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1670032574
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1670032574
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1670032574
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1670032574
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1670032574
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1670032574
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1670032574
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1670032574
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1670032574
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1670032574
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1670032574
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1670032574
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1670032574
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1670032574
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1670032574
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1670032574
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1670032574
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1670032574
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1670032574
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1670032574
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1670032574
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1670032574
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1670032574
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1670032574
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1670032574
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1670032574
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1670032574
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1670032574
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1670032574
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1670032574
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1670032574
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1670032574
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1670032574
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1670032574
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1670032574
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1670032574
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1670032574
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_573
timestamp 1670032574
transform 1 0 53820 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_577
timestamp 1670032574
transform 1 0 54188 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_588
timestamp 1670032574
transform 1 0 55200 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_614
timestamp 1670032574
transform 1 0 57592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_617
timestamp 1670032574
transform 1 0 57868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_623
timestamp 1670032574
transform 1 0 58420 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1670032574
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1670032574
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1670032574
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1670032574
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1670032574
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1670032574
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1670032574
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1670032574
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1670032574
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1670032574
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1670032574
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1670032574
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1670032574
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1670032574
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1670032574
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1670032574
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1670032574
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1670032574
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1670032574
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1670032574
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1670032574
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1670032574
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1670032574
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1670032574
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1670032574
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1670032574
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1670032574
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1670032574
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1670032574
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1670032574
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1670032574
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1670032574
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1670032574
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1670032574
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1670032574
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1670032574
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1670032574
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1670032574
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1670032574
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1670032574
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1670032574
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1670032574
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1670032574
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1670032574
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1670032574
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1670032574
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1670032574
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1670032574
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1670032574
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1670032574
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1670032574
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1670032574
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1670032574
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1670032574
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1670032574
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1670032574
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1670032574
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1670032574
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1670032574
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1670032574
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1670032574
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1670032574
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1670032574
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1670032574
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_589
timestamp 1670032574
transform 1 0 55292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_593
timestamp 1670032574
transform 1 0 55660 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_596
timestamp 1670032574
transform 1 0 55936 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_623
timestamp 1670032574
transform 1 0 58420 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1670032574
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1670032574
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1670032574
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1670032574
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1670032574
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1670032574
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1670032574
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1670032574
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1670032574
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1670032574
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1670032574
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1670032574
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1670032574
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1670032574
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1670032574
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1670032574
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1670032574
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1670032574
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1670032574
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1670032574
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1670032574
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1670032574
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1670032574
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1670032574
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1670032574
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1670032574
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1670032574
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1670032574
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1670032574
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1670032574
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1670032574
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1670032574
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1670032574
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1670032574
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1670032574
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1670032574
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1670032574
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1670032574
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1670032574
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1670032574
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1670032574
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1670032574
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1670032574
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1670032574
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1670032574
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1670032574
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1670032574
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1670032574
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1670032574
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1670032574
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1670032574
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1670032574
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1670032574
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1670032574
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1670032574
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1670032574
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1670032574
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1670032574
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1670032574
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1670032574
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1670032574
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1670032574
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1670032574
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_597
timestamp 1670032574
transform 1 0 56028 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_600
timestamp 1670032574
transform 1 0 56304 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_606
timestamp 1670032574
transform 1 0 56856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_614
timestamp 1670032574
transform 1 0 57592 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_617
timestamp 1670032574
transform 1 0 57868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_623
timestamp 1670032574
transform 1 0 58420 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1670032574
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_9
timestamp 1670032574
transform 1 0 1932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1670032574
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1670032574
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1670032574
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1670032574
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1670032574
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1670032574
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1670032574
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1670032574
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1670032574
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1670032574
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1670032574
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1670032574
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1670032574
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1670032574
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1670032574
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1670032574
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1670032574
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1670032574
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1670032574
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1670032574
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1670032574
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1670032574
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1670032574
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1670032574
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1670032574
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1670032574
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1670032574
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1670032574
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1670032574
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1670032574
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1670032574
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1670032574
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1670032574
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1670032574
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1670032574
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1670032574
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1670032574
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1670032574
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1670032574
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1670032574
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1670032574
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1670032574
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1670032574
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1670032574
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1670032574
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1670032574
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1670032574
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1670032574
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1670032574
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1670032574
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1670032574
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1670032574
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1670032574
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1670032574
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1670032574
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1670032574
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1670032574
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1670032574
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1670032574
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_569
timestamp 1670032574
transform 1 0 53452 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_579
timestamp 1670032574
transform 1 0 54372 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1670032574
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1670032574
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_601
timestamp 1670032574
transform 1 0 56396 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_607
timestamp 1670032574
transform 1 0 56948 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_610
timestamp 1670032574
transform 1 0 57224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_616
timestamp 1670032574
transform 1 0 57776 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_623
timestamp 1670032574
transform 1 0 58420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1670032574
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1670032574
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1670032574
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1670032574
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1670032574
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1670032574
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1670032574
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1670032574
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1670032574
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1670032574
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1670032574
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1670032574
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1670032574
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1670032574
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1670032574
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1670032574
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1670032574
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1670032574
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1670032574
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1670032574
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1670032574
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1670032574
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1670032574
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1670032574
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1670032574
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1670032574
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1670032574
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1670032574
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1670032574
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1670032574
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1670032574
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1670032574
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1670032574
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1670032574
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1670032574
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1670032574
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1670032574
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1670032574
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1670032574
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1670032574
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1670032574
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1670032574
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1670032574
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1670032574
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1670032574
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1670032574
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1670032574
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1670032574
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1670032574
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1670032574
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1670032574
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1670032574
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1670032574
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1670032574
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1670032574
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1670032574
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1670032574
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1670032574
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_541
timestamp 1670032574
transform 1 0 50876 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_547
timestamp 1670032574
transform 1 0 51428 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_558
timestamp 1670032574
transform 1 0 52440 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1670032574
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_575
timestamp 1670032574
transform 1 0 54004 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_600
timestamp 1670032574
transform 1 0 56304 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_606
timestamp 1670032574
transform 1 0 56856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_614
timestamp 1670032574
transform 1 0 57592 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_617
timestamp 1670032574
transform 1 0 57868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1670032574
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1670032574
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1670032574
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1670032574
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1670032574
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1670032574
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1670032574
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1670032574
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1670032574
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1670032574
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1670032574
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1670032574
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1670032574
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1670032574
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1670032574
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1670032574
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1670032574
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1670032574
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1670032574
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1670032574
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1670032574
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1670032574
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1670032574
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1670032574
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1670032574
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1670032574
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1670032574
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1670032574
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1670032574
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1670032574
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1670032574
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1670032574
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1670032574
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1670032574
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1670032574
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1670032574
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1670032574
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1670032574
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1670032574
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1670032574
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1670032574
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1670032574
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1670032574
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1670032574
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1670032574
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1670032574
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1670032574
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1670032574
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1670032574
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1670032574
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1670032574
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1670032574
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1670032574
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1670032574
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1670032574
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1670032574
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1670032574
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1670032574
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1670032574
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1670032574
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1670032574
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_569
timestamp 1670032574
transform 1 0 53452 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_585
timestamp 1670032574
transform 1 0 54924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_589
timestamp 1670032574
transform 1 0 55292 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_593
timestamp 1670032574
transform 1 0 55660 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_596
timestamp 1670032574
transform 1 0 55936 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1670032574
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1670032574
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1670032574
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1670032574
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1670032574
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1670032574
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1670032574
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1670032574
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1670032574
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1670032574
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1670032574
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1670032574
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1670032574
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1670032574
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1670032574
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1670032574
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1670032574
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1670032574
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1670032574
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1670032574
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1670032574
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1670032574
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1670032574
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1670032574
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1670032574
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1670032574
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1670032574
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1670032574
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1670032574
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1670032574
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1670032574
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1670032574
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1670032574
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1670032574
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1670032574
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1670032574
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1670032574
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1670032574
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1670032574
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1670032574
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1670032574
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1670032574
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1670032574
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1670032574
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1670032574
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1670032574
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1670032574
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1670032574
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1670032574
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1670032574
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1670032574
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1670032574
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1670032574
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1670032574
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1670032574
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1670032574
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1670032574
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1670032574
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1670032574
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1670032574
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1670032574
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1670032574
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1670032574
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1670032574
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1670032574
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_597
timestamp 1670032574
transform 1 0 56028 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_600
timestamp 1670032574
transform 1 0 56304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_614
timestamp 1670032574
transform 1 0 57592 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_617
timestamp 1670032574
transform 1 0 57868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_623
timestamp 1670032574
transform 1 0 58420 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1670032574
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1670032574
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1670032574
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1670032574
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1670032574
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1670032574
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1670032574
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1670032574
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1670032574
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1670032574
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1670032574
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1670032574
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1670032574
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1670032574
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1670032574
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1670032574
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1670032574
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1670032574
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1670032574
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1670032574
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1670032574
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1670032574
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1670032574
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1670032574
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1670032574
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1670032574
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1670032574
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1670032574
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1670032574
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1670032574
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1670032574
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1670032574
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1670032574
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1670032574
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1670032574
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1670032574
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1670032574
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1670032574
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1670032574
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1670032574
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1670032574
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1670032574
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1670032574
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1670032574
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1670032574
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1670032574
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1670032574
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1670032574
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1670032574
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1670032574
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1670032574
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1670032574
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1670032574
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1670032574
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1670032574
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1670032574
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1670032574
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1670032574
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1670032574
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1670032574
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1670032574
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1670032574
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1670032574
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1670032574
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1670032574
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_601
timestamp 1670032574
transform 1 0 56396 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_607
timestamp 1670032574
transform 1 0 56948 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_610
timestamp 1670032574
transform 1 0 57224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_616
timestamp 1670032574
transform 1 0 57776 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_623
timestamp 1670032574
transform 1 0 58420 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1670032574
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1670032574
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1670032574
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1670032574
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1670032574
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1670032574
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1670032574
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1670032574
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1670032574
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1670032574
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1670032574
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1670032574
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1670032574
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1670032574
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1670032574
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1670032574
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1670032574
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1670032574
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1670032574
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1670032574
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1670032574
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1670032574
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1670032574
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1670032574
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1670032574
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1670032574
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1670032574
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1670032574
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1670032574
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1670032574
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1670032574
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1670032574
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1670032574
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1670032574
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1670032574
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1670032574
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1670032574
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1670032574
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1670032574
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1670032574
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1670032574
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1670032574
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1670032574
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1670032574
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1670032574
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1670032574
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1670032574
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1670032574
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1670032574
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1670032574
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1670032574
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1670032574
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1670032574
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1670032574
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1670032574
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1670032574
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1670032574
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1670032574
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1670032574
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1670032574
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1670032574
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1670032574
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1670032574
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_597
timestamp 1670032574
transform 1 0 56028 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_605
timestamp 1670032574
transform 1 0 56764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_611
timestamp 1670032574
transform 1 0 57316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_614
timestamp 1670032574
transform 1 0 57592 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_617
timestamp 1670032574
transform 1 0 57868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_623
timestamp 1670032574
transform 1 0 58420 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1670032574
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1670032574
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1670032574
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1670032574
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1670032574
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1670032574
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1670032574
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1670032574
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1670032574
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1670032574
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1670032574
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1670032574
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1670032574
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1670032574
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1670032574
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1670032574
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1670032574
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1670032574
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1670032574
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1670032574
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1670032574
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1670032574
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1670032574
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1670032574
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1670032574
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1670032574
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1670032574
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1670032574
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1670032574
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1670032574
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1670032574
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1670032574
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1670032574
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1670032574
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1670032574
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1670032574
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1670032574
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1670032574
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1670032574
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1670032574
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1670032574
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1670032574
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1670032574
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1670032574
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1670032574
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1670032574
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1670032574
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1670032574
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1670032574
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1670032574
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1670032574
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1670032574
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1670032574
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1670032574
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1670032574
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1670032574
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1670032574
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1670032574
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1670032574
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1670032574
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1670032574
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_569
timestamp 1670032574
transform 1 0 53452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_577
timestamp 1670032574
transform 1 0 54188 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_580
timestamp 1670032574
transform 1 0 54464 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_589
timestamp 1670032574
transform 1 0 55292 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_597
timestamp 1670032574
transform 1 0 56028 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_601
timestamp 1670032574
transform 1 0 56396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_623
timestamp 1670032574
transform 1 0 58420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1670032574
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_9
timestamp 1670032574
transform 1 0 1932 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1670032574
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1670032574
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1670032574
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1670032574
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1670032574
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1670032574
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1670032574
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1670032574
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1670032574
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1670032574
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1670032574
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1670032574
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1670032574
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1670032574
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1670032574
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1670032574
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1670032574
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1670032574
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1670032574
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1670032574
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1670032574
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1670032574
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1670032574
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1670032574
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1670032574
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1670032574
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1670032574
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1670032574
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1670032574
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1670032574
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1670032574
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1670032574
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1670032574
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1670032574
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1670032574
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1670032574
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1670032574
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1670032574
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1670032574
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1670032574
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1670032574
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1670032574
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1670032574
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1670032574
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1670032574
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1670032574
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1670032574
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1670032574
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1670032574
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1670032574
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1670032574
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1670032574
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1670032574
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1670032574
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1670032574
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1670032574
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1670032574
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1670032574
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1670032574
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1670032574
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_573
timestamp 1670032574
transform 1 0 53820 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_576
timestamp 1670032574
transform 1 0 54096 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_598
timestamp 1670032574
transform 1 0 56120 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_604
timestamp 1670032574
transform 1 0 56672 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_614
timestamp 1670032574
transform 1 0 57592 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_617
timestamp 1670032574
transform 1 0 57868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_623
timestamp 1670032574
transform 1 0 58420 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1670032574
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1670032574
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1670032574
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1670032574
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1670032574
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1670032574
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1670032574
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1670032574
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1670032574
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1670032574
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1670032574
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1670032574
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1670032574
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1670032574
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1670032574
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1670032574
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1670032574
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1670032574
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1670032574
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1670032574
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1670032574
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1670032574
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1670032574
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1670032574
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1670032574
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1670032574
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1670032574
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1670032574
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1670032574
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1670032574
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1670032574
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1670032574
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1670032574
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1670032574
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1670032574
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1670032574
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1670032574
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1670032574
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1670032574
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1670032574
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1670032574
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1670032574
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1670032574
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1670032574
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1670032574
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1670032574
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1670032574
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1670032574
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1670032574
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1670032574
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1670032574
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1670032574
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1670032574
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1670032574
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1670032574
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1670032574
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1670032574
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1670032574
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1670032574
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1670032574
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1670032574
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1670032574
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1670032574
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_589
timestamp 1670032574
transform 1 0 55292 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_595
timestamp 1670032574
transform 1 0 55844 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_601
timestamp 1670032574
transform 1 0 56396 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_623
timestamp 1670032574
transform 1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1670032574
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_9
timestamp 1670032574
transform 1 0 1932 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1670032574
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1670032574
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1670032574
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1670032574
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1670032574
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1670032574
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1670032574
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1670032574
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1670032574
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1670032574
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1670032574
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1670032574
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1670032574
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1670032574
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1670032574
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1670032574
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1670032574
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1670032574
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1670032574
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1670032574
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1670032574
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1670032574
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1670032574
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1670032574
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1670032574
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1670032574
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1670032574
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1670032574
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1670032574
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1670032574
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1670032574
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1670032574
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1670032574
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1670032574
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1670032574
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1670032574
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1670032574
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1670032574
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1670032574
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1670032574
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1670032574
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1670032574
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1670032574
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1670032574
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1670032574
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1670032574
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1670032574
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1670032574
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1670032574
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1670032574
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1670032574
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1670032574
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1670032574
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1670032574
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1670032574
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1670032574
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1670032574
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1670032574
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1670032574
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1670032574
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1670032574
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_585
timestamp 1670032574
transform 1 0 54924 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_591
timestamp 1670032574
transform 1 0 55476 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_605
timestamp 1670032574
transform 1 0 56764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_611
timestamp 1670032574
transform 1 0 57316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_614
timestamp 1670032574
transform 1 0 57592 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_617
timestamp 1670032574
transform 1 0 57868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_623
timestamp 1670032574
transform 1 0 58420 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1670032574
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_9
timestamp 1670032574
transform 1 0 1932 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1670032574
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1670032574
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1670032574
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1670032574
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1670032574
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1670032574
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1670032574
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1670032574
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1670032574
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1670032574
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1670032574
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1670032574
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1670032574
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1670032574
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1670032574
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1670032574
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1670032574
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1670032574
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1670032574
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1670032574
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1670032574
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1670032574
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1670032574
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1670032574
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1670032574
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1670032574
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1670032574
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1670032574
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1670032574
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1670032574
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1670032574
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1670032574
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1670032574
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1670032574
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1670032574
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1670032574
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1670032574
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1670032574
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1670032574
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1670032574
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1670032574
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1670032574
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1670032574
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1670032574
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1670032574
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1670032574
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1670032574
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1670032574
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1670032574
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1670032574
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1670032574
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1670032574
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1670032574
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1670032574
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1670032574
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1670032574
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1670032574
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1670032574
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1670032574
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1670032574
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_581
timestamp 1670032574
transform 1 0 54556 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_586
timestamp 1670032574
transform 1 0 55016 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_589
timestamp 1670032574
transform 1 0 55292 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_609
timestamp 1670032574
transform 1 0 57132 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_615
timestamp 1670032574
transform 1 0 57684 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_619
timestamp 1670032574
transform 1 0 58052 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_623
timestamp 1670032574
transform 1 0 58420 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1670032574
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1670032574
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1670032574
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1670032574
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1670032574
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1670032574
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1670032574
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1670032574
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1670032574
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1670032574
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1670032574
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1670032574
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1670032574
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1670032574
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1670032574
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1670032574
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1670032574
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1670032574
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1670032574
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1670032574
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1670032574
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1670032574
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1670032574
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1670032574
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1670032574
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1670032574
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1670032574
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1670032574
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1670032574
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1670032574
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1670032574
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1670032574
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1670032574
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1670032574
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1670032574
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1670032574
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1670032574
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1670032574
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1670032574
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1670032574
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1670032574
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1670032574
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1670032574
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1670032574
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1670032574
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1670032574
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1670032574
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1670032574
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1670032574
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1670032574
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1670032574
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1670032574
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1670032574
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1670032574
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1670032574
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1670032574
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1670032574
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1670032574
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1670032574
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1670032574
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1670032574
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1670032574
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1670032574
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1670032574
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_609
timestamp 1670032574
transform 1 0 57132 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_614
timestamp 1670032574
transform 1 0 57592 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_617
timestamp 1670032574
transform 1 0 57868 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_623
timestamp 1670032574
transform 1 0 58420 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1670032574
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_9
timestamp 1670032574
transform 1 0 1932 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1670032574
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1670032574
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1670032574
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1670032574
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1670032574
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1670032574
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1670032574
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1670032574
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1670032574
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1670032574
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1670032574
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1670032574
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1670032574
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1670032574
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1670032574
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1670032574
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1670032574
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1670032574
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1670032574
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1670032574
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1670032574
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1670032574
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1670032574
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1670032574
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1670032574
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1670032574
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1670032574
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1670032574
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1670032574
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1670032574
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1670032574
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1670032574
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1670032574
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1670032574
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1670032574
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1670032574
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1670032574
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1670032574
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1670032574
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1670032574
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1670032574
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1670032574
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1670032574
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1670032574
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1670032574
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1670032574
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1670032574
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1670032574
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1670032574
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1670032574
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1670032574
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1670032574
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1670032574
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1670032574
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1670032574
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1670032574
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1670032574
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1670032574
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1670032574
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1670032574
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1670032574
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1670032574
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1670032574
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1670032574
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_613
timestamp 1670032574
transform 1 0 57500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_616
timestamp 1670032574
transform 1 0 57776 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_623
timestamp 1670032574
transform 1 0 58420 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1670032574
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_9
timestamp 1670032574
transform 1 0 1932 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1670032574
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1670032574
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1670032574
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1670032574
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1670032574
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1670032574
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1670032574
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1670032574
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1670032574
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1670032574
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1670032574
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1670032574
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1670032574
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1670032574
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1670032574
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1670032574
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1670032574
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1670032574
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1670032574
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1670032574
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1670032574
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1670032574
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1670032574
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1670032574
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1670032574
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1670032574
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1670032574
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1670032574
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1670032574
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1670032574
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1670032574
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1670032574
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1670032574
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1670032574
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1670032574
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1670032574
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1670032574
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1670032574
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1670032574
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1670032574
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1670032574
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1670032574
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1670032574
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1670032574
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1670032574
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1670032574
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1670032574
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1670032574
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1670032574
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1670032574
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1670032574
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1670032574
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1670032574
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1670032574
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1670032574
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1670032574
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1670032574
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1670032574
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1670032574
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1670032574
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1670032574
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1670032574
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1670032574
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1670032574
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1670032574
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_617
timestamp 1670032574
transform 1 0 57868 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_623
timestamp 1670032574
transform 1 0 58420 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1670032574
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1670032574
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1670032574
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1670032574
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1670032574
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1670032574
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1670032574
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1670032574
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1670032574
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1670032574
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1670032574
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1670032574
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1670032574
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1670032574
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1670032574
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1670032574
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1670032574
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1670032574
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1670032574
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1670032574
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1670032574
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1670032574
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1670032574
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1670032574
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1670032574
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1670032574
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1670032574
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1670032574
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1670032574
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1670032574
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1670032574
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1670032574
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1670032574
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1670032574
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1670032574
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1670032574
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1670032574
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1670032574
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1670032574
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1670032574
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1670032574
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1670032574
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1670032574
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1670032574
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1670032574
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1670032574
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1670032574
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1670032574
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1670032574
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1670032574
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1670032574
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1670032574
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1670032574
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1670032574
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1670032574
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1670032574
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1670032574
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1670032574
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1670032574
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1670032574
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1670032574
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1670032574
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1670032574
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1670032574
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1670032574
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_613
timestamp 1670032574
transform 1 0 57500 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_623
timestamp 1670032574
transform 1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1670032574
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_9
timestamp 1670032574
transform 1 0 1932 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1670032574
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1670032574
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1670032574
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1670032574
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1670032574
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1670032574
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1670032574
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1670032574
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1670032574
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1670032574
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1670032574
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1670032574
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1670032574
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1670032574
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1670032574
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1670032574
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1670032574
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1670032574
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1670032574
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1670032574
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1670032574
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1670032574
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1670032574
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1670032574
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1670032574
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1670032574
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1670032574
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1670032574
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1670032574
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1670032574
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1670032574
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1670032574
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1670032574
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1670032574
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1670032574
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1670032574
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1670032574
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1670032574
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1670032574
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1670032574
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1670032574
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1670032574
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1670032574
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1670032574
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1670032574
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1670032574
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1670032574
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1670032574
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1670032574
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1670032574
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1670032574
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1670032574
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1670032574
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1670032574
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1670032574
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1670032574
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1670032574
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1670032574
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1670032574
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1670032574
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1670032574
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1670032574
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1670032574
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_609
timestamp 1670032574
transform 1 0 57132 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_614
timestamp 1670032574
transform 1 0 57592 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_617
timestamp 1670032574
transform 1 0 57868 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_623
timestamp 1670032574
transform 1 0 58420 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1670032574
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_9
timestamp 1670032574
transform 1 0 1932 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1670032574
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1670032574
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1670032574
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1670032574
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1670032574
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1670032574
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1670032574
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1670032574
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1670032574
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1670032574
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1670032574
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1670032574
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1670032574
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1670032574
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1670032574
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1670032574
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1670032574
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1670032574
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1670032574
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1670032574
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1670032574
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1670032574
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1670032574
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1670032574
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1670032574
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1670032574
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1670032574
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1670032574
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1670032574
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1670032574
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1670032574
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1670032574
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1670032574
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1670032574
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1670032574
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1670032574
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1670032574
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1670032574
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1670032574
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1670032574
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1670032574
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1670032574
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1670032574
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1670032574
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1670032574
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1670032574
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1670032574
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1670032574
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1670032574
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1670032574
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1670032574
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1670032574
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1670032574
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1670032574
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1670032574
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1670032574
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1670032574
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1670032574
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1670032574
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1670032574
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1670032574
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1670032574
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1670032574
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1670032574
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_613
timestamp 1670032574
transform 1 0 57500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_616
timestamp 1670032574
transform 1 0 57776 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_623
timestamp 1670032574
transform 1 0 58420 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1670032574
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1670032574
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1670032574
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1670032574
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1670032574
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1670032574
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1670032574
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1670032574
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1670032574
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1670032574
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1670032574
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1670032574
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1670032574
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1670032574
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1670032574
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1670032574
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1670032574
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1670032574
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1670032574
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1670032574
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1670032574
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1670032574
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1670032574
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1670032574
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1670032574
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1670032574
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1670032574
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1670032574
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1670032574
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1670032574
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1670032574
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1670032574
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1670032574
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1670032574
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1670032574
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1670032574
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1670032574
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1670032574
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1670032574
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1670032574
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1670032574
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1670032574
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1670032574
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1670032574
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1670032574
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1670032574
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1670032574
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1670032574
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1670032574
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1670032574
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1670032574
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1670032574
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1670032574
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1670032574
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1670032574
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1670032574
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1670032574
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1670032574
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1670032574
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1670032574
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1670032574
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1670032574
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1670032574
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1670032574
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1670032574
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1670032574
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1670032574
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1670032574
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_9
timestamp 1670032574
transform 1 0 1932 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1670032574
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1670032574
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1670032574
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1670032574
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1670032574
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1670032574
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1670032574
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1670032574
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1670032574
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1670032574
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1670032574
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1670032574
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1670032574
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1670032574
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1670032574
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1670032574
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1670032574
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1670032574
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1670032574
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1670032574
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1670032574
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1670032574
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1670032574
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1670032574
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1670032574
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1670032574
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1670032574
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1670032574
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1670032574
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1670032574
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1670032574
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1670032574
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1670032574
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1670032574
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1670032574
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1670032574
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1670032574
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1670032574
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1670032574
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1670032574
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1670032574
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1670032574
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1670032574
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1670032574
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1670032574
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1670032574
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1670032574
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1670032574
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1670032574
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1670032574
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1670032574
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1670032574
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1670032574
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1670032574
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1670032574
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1670032574
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1670032574
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1670032574
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1670032574
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1670032574
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1670032574
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1670032574
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1670032574
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1670032574
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_613
timestamp 1670032574
transform 1 0 57500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_616
timestamp 1670032574
transform 1 0 57776 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_623
timestamp 1670032574
transform 1 0 58420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1670032574
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_9
timestamp 1670032574
transform 1 0 1932 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1670032574
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1670032574
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1670032574
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1670032574
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1670032574
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1670032574
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1670032574
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1670032574
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1670032574
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1670032574
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1670032574
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1670032574
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1670032574
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1670032574
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1670032574
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1670032574
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1670032574
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1670032574
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1670032574
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1670032574
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1670032574
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1670032574
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1670032574
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1670032574
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1670032574
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1670032574
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1670032574
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1670032574
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1670032574
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1670032574
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1670032574
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1670032574
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1670032574
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1670032574
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1670032574
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1670032574
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1670032574
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1670032574
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1670032574
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1670032574
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1670032574
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1670032574
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1670032574
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1670032574
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1670032574
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1670032574
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1670032574
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1670032574
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1670032574
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1670032574
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1670032574
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1670032574
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1670032574
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1670032574
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1670032574
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1670032574
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1670032574
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1670032574
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1670032574
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1670032574
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1670032574
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1670032574
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1670032574
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1670032574
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1670032574
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_617
timestamp 1670032574
transform 1 0 57868 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_623
timestamp 1670032574
transform 1 0 58420 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1670032574
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1670032574
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1670032574
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1670032574
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1670032574
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1670032574
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1670032574
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1670032574
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1670032574
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1670032574
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1670032574
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1670032574
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1670032574
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1670032574
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1670032574
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1670032574
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1670032574
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1670032574
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1670032574
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1670032574
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1670032574
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1670032574
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1670032574
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1670032574
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1670032574
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1670032574
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1670032574
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1670032574
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1670032574
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1670032574
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1670032574
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1670032574
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1670032574
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1670032574
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1670032574
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1670032574
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1670032574
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1670032574
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1670032574
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1670032574
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1670032574
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1670032574
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1670032574
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1670032574
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1670032574
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1670032574
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1670032574
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1670032574
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1670032574
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1670032574
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1670032574
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1670032574
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1670032574
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1670032574
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1670032574
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1670032574
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1670032574
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1670032574
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1670032574
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1670032574
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1670032574
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1670032574
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1670032574
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1670032574
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1670032574
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_613
timestamp 1670032574
transform 1 0 57500 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_623
timestamp 1670032574
transform 1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1670032574
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_9
timestamp 1670032574
transform 1 0 1932 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1670032574
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1670032574
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1670032574
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1670032574
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1670032574
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1670032574
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1670032574
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1670032574
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1670032574
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1670032574
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1670032574
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1670032574
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1670032574
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1670032574
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1670032574
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1670032574
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1670032574
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1670032574
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1670032574
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1670032574
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1670032574
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1670032574
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1670032574
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1670032574
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1670032574
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1670032574
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1670032574
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1670032574
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1670032574
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1670032574
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1670032574
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1670032574
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1670032574
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1670032574
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1670032574
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1670032574
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1670032574
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1670032574
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1670032574
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1670032574
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1670032574
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1670032574
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1670032574
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1670032574
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1670032574
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1670032574
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1670032574
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1670032574
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1670032574
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1670032574
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1670032574
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1670032574
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1670032574
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1670032574
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1670032574
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1670032574
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1670032574
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1670032574
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1670032574
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1670032574
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1670032574
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1670032574
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1670032574
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_609
timestamp 1670032574
transform 1 0 57132 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_614
timestamp 1670032574
transform 1 0 57592 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_617
timestamp 1670032574
transform 1 0 57868 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_623
timestamp 1670032574
transform 1 0 58420 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1670032574
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_9
timestamp 1670032574
transform 1 0 1932 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1670032574
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1670032574
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1670032574
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1670032574
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1670032574
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1670032574
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1670032574
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1670032574
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1670032574
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1670032574
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1670032574
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1670032574
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1670032574
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1670032574
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1670032574
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1670032574
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1670032574
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1670032574
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1670032574
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1670032574
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1670032574
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1670032574
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1670032574
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1670032574
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1670032574
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1670032574
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1670032574
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1670032574
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1670032574
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1670032574
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1670032574
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1670032574
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1670032574
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1670032574
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1670032574
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1670032574
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1670032574
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1670032574
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1670032574
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1670032574
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1670032574
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1670032574
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1670032574
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1670032574
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1670032574
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1670032574
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1670032574
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1670032574
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1670032574
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1670032574
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1670032574
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1670032574
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1670032574
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1670032574
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1670032574
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1670032574
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1670032574
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1670032574
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1670032574
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1670032574
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1670032574
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1670032574
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1670032574
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1670032574
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_613
timestamp 1670032574
transform 1 0 57500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_616
timestamp 1670032574
transform 1 0 57776 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_623
timestamp 1670032574
transform 1 0 58420 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1670032574
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1670032574
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1670032574
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1670032574
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1670032574
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1670032574
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1670032574
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1670032574
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1670032574
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1670032574
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1670032574
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1670032574
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1670032574
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1670032574
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1670032574
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1670032574
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1670032574
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1670032574
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1670032574
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1670032574
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1670032574
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1670032574
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1670032574
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1670032574
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1670032574
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1670032574
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1670032574
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1670032574
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1670032574
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1670032574
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1670032574
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1670032574
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1670032574
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1670032574
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1670032574
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1670032574
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1670032574
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1670032574
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1670032574
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1670032574
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1670032574
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1670032574
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1670032574
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1670032574
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1670032574
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1670032574
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1670032574
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1670032574
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1670032574
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1670032574
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1670032574
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1670032574
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1670032574
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1670032574
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1670032574
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1670032574
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1670032574
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1670032574
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1670032574
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1670032574
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1670032574
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1670032574
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1670032574
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1670032574
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1670032574
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1670032574
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1670032574
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1670032574
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_9
timestamp 1670032574
transform 1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1670032574
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1670032574
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1670032574
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1670032574
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1670032574
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1670032574
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1670032574
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1670032574
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1670032574
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1670032574
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1670032574
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1670032574
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1670032574
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1670032574
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1670032574
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1670032574
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1670032574
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1670032574
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1670032574
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1670032574
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1670032574
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1670032574
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1670032574
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1670032574
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1670032574
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1670032574
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1670032574
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1670032574
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1670032574
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1670032574
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1670032574
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1670032574
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1670032574
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1670032574
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1670032574
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1670032574
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1670032574
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1670032574
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1670032574
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1670032574
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1670032574
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1670032574
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1670032574
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1670032574
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1670032574
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1670032574
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1670032574
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1670032574
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1670032574
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1670032574
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1670032574
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1670032574
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1670032574
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1670032574
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1670032574
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1670032574
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1670032574
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1670032574
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1670032574
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1670032574
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1670032574
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1670032574
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1670032574
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1670032574
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_613
timestamp 1670032574
transform 1 0 57500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_616
timestamp 1670032574
transform 1 0 57776 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_623
timestamp 1670032574
transform 1 0 58420 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1670032574
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_9
timestamp 1670032574
transform 1 0 1932 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1670032574
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1670032574
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1670032574
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1670032574
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1670032574
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1670032574
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1670032574
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1670032574
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1670032574
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1670032574
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1670032574
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1670032574
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1670032574
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1670032574
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1670032574
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1670032574
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1670032574
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1670032574
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1670032574
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1670032574
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1670032574
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1670032574
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1670032574
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1670032574
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1670032574
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1670032574
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1670032574
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1670032574
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1670032574
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1670032574
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1670032574
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1670032574
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1670032574
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1670032574
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1670032574
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1670032574
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1670032574
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1670032574
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1670032574
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1670032574
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1670032574
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1670032574
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1670032574
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1670032574
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1670032574
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1670032574
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1670032574
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1670032574
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1670032574
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1670032574
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1670032574
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1670032574
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1670032574
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1670032574
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1670032574
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1670032574
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1670032574
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1670032574
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1670032574
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1670032574
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1670032574
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1670032574
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1670032574
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1670032574
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1670032574
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_617
timestamp 1670032574
transform 1 0 57868 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_623
timestamp 1670032574
transform 1 0 58420 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1670032574
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1670032574
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1670032574
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1670032574
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1670032574
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1670032574
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1670032574
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1670032574
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1670032574
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1670032574
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1670032574
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1670032574
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1670032574
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1670032574
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1670032574
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1670032574
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1670032574
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1670032574
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1670032574
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1670032574
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1670032574
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1670032574
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1670032574
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1670032574
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1670032574
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1670032574
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1670032574
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1670032574
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1670032574
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1670032574
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1670032574
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1670032574
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1670032574
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1670032574
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1670032574
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1670032574
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1670032574
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1670032574
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1670032574
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1670032574
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1670032574
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1670032574
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1670032574
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1670032574
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1670032574
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1670032574
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1670032574
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1670032574
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1670032574
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1670032574
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1670032574
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1670032574
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1670032574
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1670032574
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1670032574
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1670032574
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1670032574
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1670032574
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1670032574
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1670032574
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1670032574
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1670032574
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1670032574
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1670032574
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1670032574
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_613
timestamp 1670032574
transform 1 0 57500 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_623
timestamp 1670032574
transform 1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1670032574
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_9
timestamp 1670032574
transform 1 0 1932 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1670032574
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1670032574
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1670032574
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1670032574
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1670032574
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1670032574
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1670032574
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1670032574
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1670032574
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1670032574
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1670032574
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1670032574
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1670032574
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1670032574
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1670032574
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1670032574
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1670032574
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1670032574
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1670032574
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1670032574
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1670032574
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1670032574
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1670032574
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1670032574
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1670032574
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1670032574
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1670032574
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1670032574
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1670032574
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1670032574
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1670032574
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1670032574
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1670032574
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1670032574
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1670032574
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1670032574
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1670032574
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1670032574
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1670032574
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1670032574
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1670032574
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1670032574
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1670032574
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1670032574
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1670032574
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1670032574
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1670032574
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1670032574
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1670032574
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1670032574
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1670032574
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1670032574
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1670032574
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1670032574
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1670032574
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1670032574
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1670032574
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1670032574
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1670032574
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1670032574
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1670032574
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1670032574
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1670032574
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_609
timestamp 1670032574
transform 1 0 57132 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_614
timestamp 1670032574
transform 1 0 57592 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_85_617
timestamp 1670032574
transform 1 0 57868 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_623
timestamp 1670032574
transform 1 0 58420 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1670032574
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_9
timestamp 1670032574
transform 1 0 1932 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1670032574
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1670032574
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1670032574
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1670032574
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1670032574
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1670032574
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1670032574
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1670032574
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1670032574
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1670032574
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1670032574
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1670032574
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1670032574
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1670032574
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1670032574
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1670032574
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1670032574
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1670032574
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1670032574
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1670032574
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1670032574
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1670032574
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1670032574
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1670032574
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1670032574
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1670032574
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1670032574
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1670032574
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1670032574
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1670032574
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1670032574
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1670032574
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1670032574
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1670032574
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1670032574
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1670032574
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1670032574
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1670032574
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1670032574
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1670032574
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1670032574
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1670032574
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1670032574
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1670032574
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1670032574
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1670032574
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1670032574
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1670032574
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1670032574
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1670032574
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1670032574
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1670032574
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1670032574
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1670032574
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1670032574
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1670032574
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1670032574
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1670032574
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1670032574
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1670032574
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1670032574
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1670032574
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1670032574
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1670032574
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_613
timestamp 1670032574
transform 1 0 57500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_616
timestamp 1670032574
transform 1 0 57776 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_623
timestamp 1670032574
transform 1 0 58420 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1670032574
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1670032574
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1670032574
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1670032574
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1670032574
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1670032574
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1670032574
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1670032574
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1670032574
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1670032574
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1670032574
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1670032574
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1670032574
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1670032574
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1670032574
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1670032574
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1670032574
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1670032574
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1670032574
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1670032574
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1670032574
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1670032574
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1670032574
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1670032574
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1670032574
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1670032574
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1670032574
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1670032574
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1670032574
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1670032574
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1670032574
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1670032574
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1670032574
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1670032574
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1670032574
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1670032574
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1670032574
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1670032574
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1670032574
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1670032574
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1670032574
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1670032574
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1670032574
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1670032574
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1670032574
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1670032574
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1670032574
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1670032574
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1670032574
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1670032574
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1670032574
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1670032574
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1670032574
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1670032574
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1670032574
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1670032574
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1670032574
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1670032574
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1670032574
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1670032574
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1670032574
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1670032574
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1670032574
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1670032574
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1670032574
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1670032574
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1670032574
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1670032574
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_9
timestamp 1670032574
transform 1 0 1932 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1670032574
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1670032574
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1670032574
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1670032574
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1670032574
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1670032574
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1670032574
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1670032574
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1670032574
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1670032574
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1670032574
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1670032574
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1670032574
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1670032574
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1670032574
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1670032574
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1670032574
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1670032574
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1670032574
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1670032574
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1670032574
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1670032574
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1670032574
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1670032574
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1670032574
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1670032574
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1670032574
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1670032574
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1670032574
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1670032574
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1670032574
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1670032574
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1670032574
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1670032574
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1670032574
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1670032574
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1670032574
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1670032574
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1670032574
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1670032574
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1670032574
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1670032574
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1670032574
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1670032574
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1670032574
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1670032574
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1670032574
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1670032574
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1670032574
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1670032574
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1670032574
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1670032574
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1670032574
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1670032574
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1670032574
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1670032574
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1670032574
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1670032574
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1670032574
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1670032574
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1670032574
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1670032574
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1670032574
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1670032574
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_613
timestamp 1670032574
transform 1 0 57500 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_616
timestamp 1670032574
transform 1 0 57776 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_623
timestamp 1670032574
transform 1 0 58420 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1670032574
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_9
timestamp 1670032574
transform 1 0 1932 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1670032574
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1670032574
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1670032574
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1670032574
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1670032574
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1670032574
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1670032574
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1670032574
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1670032574
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1670032574
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1670032574
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1670032574
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1670032574
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1670032574
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1670032574
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1670032574
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1670032574
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1670032574
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1670032574
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1670032574
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1670032574
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1670032574
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1670032574
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1670032574
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1670032574
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1670032574
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1670032574
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1670032574
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1670032574
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1670032574
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1670032574
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1670032574
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1670032574
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1670032574
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1670032574
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1670032574
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1670032574
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1670032574
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1670032574
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1670032574
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1670032574
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1670032574
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1670032574
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1670032574
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1670032574
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1670032574
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1670032574
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1670032574
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1670032574
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1670032574
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1670032574
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1670032574
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1670032574
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1670032574
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1670032574
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1670032574
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1670032574
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1670032574
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1670032574
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1670032574
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1670032574
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1670032574
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1670032574
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1670032574
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1670032574
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_89_617
timestamp 1670032574
transform 1 0 57868 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_623
timestamp 1670032574
transform 1 0 58420 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1670032574
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1670032574
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1670032574
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1670032574
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1670032574
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1670032574
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1670032574
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1670032574
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1670032574
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1670032574
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1670032574
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1670032574
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1670032574
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1670032574
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1670032574
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1670032574
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1670032574
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1670032574
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1670032574
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1670032574
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1670032574
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1670032574
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1670032574
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1670032574
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1670032574
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1670032574
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1670032574
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1670032574
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1670032574
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1670032574
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1670032574
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1670032574
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1670032574
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1670032574
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1670032574
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1670032574
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1670032574
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1670032574
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1670032574
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1670032574
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1670032574
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1670032574
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1670032574
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1670032574
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1670032574
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1670032574
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1670032574
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1670032574
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1670032574
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1670032574
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1670032574
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1670032574
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1670032574
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1670032574
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1670032574
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1670032574
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1670032574
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1670032574
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1670032574
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1670032574
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1670032574
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1670032574
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1670032574
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1670032574
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1670032574
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_613
timestamp 1670032574
transform 1 0 57500 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_623
timestamp 1670032574
transform 1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1670032574
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_9
timestamp 1670032574
transform 1 0 1932 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1670032574
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1670032574
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1670032574
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1670032574
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1670032574
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1670032574
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1670032574
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1670032574
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1670032574
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1670032574
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1670032574
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1670032574
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1670032574
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1670032574
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1670032574
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1670032574
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1670032574
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1670032574
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1670032574
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1670032574
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1670032574
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1670032574
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1670032574
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1670032574
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1670032574
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1670032574
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1670032574
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1670032574
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1670032574
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1670032574
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1670032574
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1670032574
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1670032574
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1670032574
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1670032574
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1670032574
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1670032574
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1670032574
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1670032574
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1670032574
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1670032574
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1670032574
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1670032574
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1670032574
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1670032574
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1670032574
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1670032574
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1670032574
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1670032574
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1670032574
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1670032574
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1670032574
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1670032574
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1670032574
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1670032574
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1670032574
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1670032574
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1670032574
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1670032574
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1670032574
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1670032574
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1670032574
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1670032574
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_609
timestamp 1670032574
transform 1 0 57132 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_614
timestamp 1670032574
transform 1 0 57592 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_91_617
timestamp 1670032574
transform 1 0 57868 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_623
timestamp 1670032574
transform 1 0 58420 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1670032574
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_9
timestamp 1670032574
transform 1 0 1932 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1670032574
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1670032574
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1670032574
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1670032574
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1670032574
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1670032574
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1670032574
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1670032574
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1670032574
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1670032574
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1670032574
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1670032574
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1670032574
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1670032574
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1670032574
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1670032574
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1670032574
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1670032574
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1670032574
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1670032574
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1670032574
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1670032574
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1670032574
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1670032574
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1670032574
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1670032574
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1670032574
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1670032574
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1670032574
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1670032574
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1670032574
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1670032574
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1670032574
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1670032574
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1670032574
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1670032574
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1670032574
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1670032574
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1670032574
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1670032574
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1670032574
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1670032574
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1670032574
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1670032574
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1670032574
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1670032574
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1670032574
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1670032574
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1670032574
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1670032574
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1670032574
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1670032574
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1670032574
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1670032574
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1670032574
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1670032574
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1670032574
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1670032574
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1670032574
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1670032574
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1670032574
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1670032574
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1670032574
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1670032574
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_613
timestamp 1670032574
transform 1 0 57500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_616
timestamp 1670032574
transform 1 0 57776 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_623
timestamp 1670032574
transform 1 0 58420 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1670032574
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1670032574
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1670032574
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1670032574
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1670032574
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1670032574
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1670032574
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1670032574
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1670032574
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1670032574
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1670032574
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1670032574
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1670032574
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1670032574
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1670032574
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1670032574
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1670032574
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1670032574
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1670032574
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1670032574
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1670032574
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1670032574
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1670032574
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1670032574
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1670032574
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1670032574
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1670032574
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1670032574
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1670032574
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1670032574
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1670032574
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_293
timestamp 1670032574
transform 1 0 28060 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_297
timestamp 1670032574
transform 1 0 28428 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_305
timestamp 1670032574
transform 1 0 29164 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_315
timestamp 1670032574
transform 1 0 30084 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_327
timestamp 1670032574
transform 1 0 31188 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1670032574
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1670032574
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1670032574
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1670032574
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1670032574
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1670032574
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1670032574
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_393
timestamp 1670032574
transform 1 0 37260 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_401
timestamp 1670032574
transform 1 0 37996 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_404
timestamp 1670032574
transform 1 0 38272 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_416
timestamp 1670032574
transform 1 0 39376 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_428
timestamp 1670032574
transform 1 0 40480 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_440
timestamp 1670032574
transform 1 0 41584 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1670032574
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1670032574
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1670032574
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1670032574
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1670032574
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1670032574
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1670032574
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1670032574
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1670032574
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1670032574
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1670032574
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1670032574
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1670032574
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1670032574
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1670032574
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1670032574
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1670032574
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1670032574
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1670032574
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1670032574
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_9
timestamp 1670032574
transform 1 0 1932 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1670032574
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1670032574
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1670032574
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1670032574
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1670032574
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1670032574
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1670032574
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1670032574
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1670032574
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1670032574
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1670032574
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1670032574
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1670032574
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1670032574
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1670032574
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1670032574
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1670032574
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1670032574
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1670032574
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1670032574
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1670032574
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1670032574
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1670032574
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1670032574
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1670032574
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1670032574
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1670032574
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_265
timestamp 1670032574
transform 1 0 25484 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_273
timestamp 1670032574
transform 1 0 26220 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_276
timestamp 1670032574
transform 1 0 26496 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_288
timestamp 1670032574
transform 1 0 27600 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_292
timestamp 1670032574
transform 1 0 27968 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_295
timestamp 1670032574
transform 1 0 28244 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_306
timestamp 1670032574
transform 1 0 29256 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_309
timestamp 1670032574
transform 1 0 29532 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_324
timestamp 1670032574
transform 1 0 30912 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_328
timestamp 1670032574
transform 1 0 31280 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_331
timestamp 1670032574
transform 1 0 31556 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_348
timestamp 1670032574
transform 1 0 33120 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_360
timestamp 1670032574
transform 1 0 34224 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1670032574
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_377
timestamp 1670032574
transform 1 0 35788 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_385
timestamp 1670032574
transform 1 0 36524 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_388
timestamp 1670032574
transform 1 0 36800 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_396
timestamp 1670032574
transform 1 0 37536 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_94_410
timestamp 1670032574
transform 1 0 38824 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_418
timestamp 1670032574
transform 1 0 39560 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_421
timestamp 1670032574
transform 1 0 39836 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_425
timestamp 1670032574
transform 1 0 40204 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_431
timestamp 1670032574
transform 1 0 40756 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_443
timestamp 1670032574
transform 1 0 41860 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_455
timestamp 1670032574
transform 1 0 42964 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_467
timestamp 1670032574
transform 1 0 44068 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1670032574
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1670032574
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1670032574
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1670032574
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1670032574
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1670032574
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1670032574
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1670032574
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1670032574
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1670032574
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1670032574
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1670032574
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1670032574
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1670032574
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1670032574
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_613
timestamp 1670032574
transform 1 0 57500 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_616
timestamp 1670032574
transform 1 0 57776 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_623
timestamp 1670032574
transform 1 0 58420 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1670032574
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_9
timestamp 1670032574
transform 1 0 1932 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1670032574
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1670032574
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1670032574
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1670032574
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1670032574
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1670032574
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1670032574
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1670032574
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1670032574
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1670032574
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1670032574
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1670032574
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1670032574
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1670032574
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1670032574
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1670032574
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1670032574
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1670032574
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1670032574
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1670032574
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1670032574
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_222
timestamp 1670032574
transform 1 0 21528 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1670032574
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_237
timestamp 1670032574
transform 1 0 22908 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_240
timestamp 1670032574
transform 1 0 23184 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_252
timestamp 1670032574
transform 1 0 24288 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_264
timestamp 1670032574
transform 1 0 25392 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_278
timestamp 1670032574
transform 1 0 26680 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_281
timestamp 1670032574
transform 1 0 26956 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_291
timestamp 1670032574
transform 1 0 27876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_303
timestamp 1670032574
transform 1 0 28980 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_311
timestamp 1670032574
transform 1 0 29716 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_323
timestamp 1670032574
transform 1 0 30820 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_327
timestamp 1670032574
transform 1 0 31188 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_334
timestamp 1670032574
transform 1 0 31832 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_337
timestamp 1670032574
transform 1 0 32108 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_347
timestamp 1670032574
transform 1 0 33028 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_353
timestamp 1670032574
transform 1 0 33580 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_359
timestamp 1670032574
transform 1 0 34132 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_368
timestamp 1670032574
transform 1 0 34960 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_380
timestamp 1670032574
transform 1 0 36064 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_393
timestamp 1670032574
transform 1 0 37260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_402
timestamp 1670032574
transform 1 0 38088 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_412
timestamp 1670032574
transform 1 0 39008 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_418
timestamp 1670032574
transform 1 0 39560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_421
timestamp 1670032574
transform 1 0 39836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_432
timestamp 1670032574
transform 1 0 40848 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_438
timestamp 1670032574
transform 1 0 41400 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_446
timestamp 1670032574
transform 1 0 42136 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1670032574
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1670032574
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1670032574
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1670032574
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1670032574
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1670032574
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1670032574
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1670032574
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1670032574
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1670032574
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1670032574
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1670032574
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1670032574
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1670032574
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1670032574
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1670032574
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1670032574
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1670032574
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_95_617
timestamp 1670032574
transform 1 0 57868 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_623
timestamp 1670032574
transform 1 0 58420 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1670032574
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1670032574
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1670032574
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1670032574
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1670032574
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1670032574
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1670032574
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1670032574
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1670032574
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1670032574
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1670032574
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1670032574
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1670032574
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1670032574
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1670032574
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1670032574
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1670032574
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1670032574
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1670032574
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1670032574
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1670032574
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1670032574
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_209
timestamp 1670032574
transform 1 0 20332 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_217
timestamp 1670032574
transform 1 0 21068 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_96_225
timestamp 1670032574
transform 1 0 21804 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_237
timestamp 1670032574
transform 1 0 22908 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_249
timestamp 1670032574
transform 1 0 24012 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_253
timestamp 1670032574
transform 1 0 24380 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_261
timestamp 1670032574
transform 1 0 25116 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_273
timestamp 1670032574
transform 1 0 26220 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_285
timestamp 1670032574
transform 1 0 27324 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_297
timestamp 1670032574
transform 1 0 28428 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_305
timestamp 1670032574
transform 1 0 29164 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1670032574
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1670032574
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_333
timestamp 1670032574
transform 1 0 31740 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_337
timestamp 1670032574
transform 1 0 32108 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_341
timestamp 1670032574
transform 1 0 32476 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_347
timestamp 1670032574
transform 1 0 33028 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_359
timestamp 1670032574
transform 1 0 34132 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1670032574
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_365
timestamp 1670032574
transform 1 0 34684 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_369
timestamp 1670032574
transform 1 0 35052 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_378
timestamp 1670032574
transform 1 0 35880 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_390
timestamp 1670032574
transform 1 0 36984 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_402
timestamp 1670032574
transform 1 0 38088 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_96_406
timestamp 1670032574
transform 1 0 38456 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_414
timestamp 1670032574
transform 1 0 39192 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_418
timestamp 1670032574
transform 1 0 39560 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_96_421
timestamp 1670032574
transform 1 0 39836 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_431
timestamp 1670032574
transform 1 0 40756 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_440
timestamp 1670032574
transform 1 0 41584 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_452
timestamp 1670032574
transform 1 0 42688 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_464
timestamp 1670032574
transform 1 0 43792 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1670032574
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1670032574
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1670032574
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1670032574
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1670032574
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1670032574
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1670032574
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1670032574
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1670032574
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1670032574
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1670032574
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1670032574
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1670032574
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1670032574
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_613
timestamp 1670032574
transform 1 0 57500 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_623
timestamp 1670032574
transform 1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_3
timestamp 1670032574
transform 1 0 1380 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_9
timestamp 1670032574
transform 1 0 1932 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1670032574
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1670032574
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1670032574
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1670032574
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1670032574
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1670032574
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1670032574
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1670032574
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1670032574
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1670032574
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1670032574
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1670032574
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1670032574
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1670032574
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1670032574
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1670032574
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1670032574
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1670032574
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1670032574
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1670032574
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1670032574
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1670032574
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1670032574
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1670032574
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1670032574
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1670032574
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1670032574
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1670032574
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1670032574
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1670032574
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1670032574
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1670032574
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1670032574
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_329
timestamp 1670032574
transform 1 0 31372 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_334
timestamp 1670032574
transform 1 0 31832 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_337
timestamp 1670032574
transform 1 0 32108 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_346
timestamp 1670032574
transform 1 0 32936 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_358
timestamp 1670032574
transform 1 0 34040 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_370
timestamp 1670032574
transform 1 0 35144 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_382
timestamp 1670032574
transform 1 0 36248 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_390
timestamp 1670032574
transform 1 0 36984 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1670032574
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1670032574
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_417
timestamp 1670032574
transform 1 0 39468 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_422
timestamp 1670032574
transform 1 0 39928 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_428
timestamp 1670032574
transform 1 0 40480 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_434
timestamp 1670032574
transform 1 0 41032 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_440
timestamp 1670032574
transform 1 0 41584 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_97_449
timestamp 1670032574
transform 1 0 42412 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_457
timestamp 1670032574
transform 1 0 43148 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_467
timestamp 1670032574
transform 1 0 44068 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_479
timestamp 1670032574
transform 1 0 45172 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_491
timestamp 1670032574
transform 1 0 46276 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1670032574
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1670032574
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1670032574
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1670032574
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1670032574
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1670032574
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1670032574
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1670032574
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1670032574
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1670032574
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1670032574
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_609
timestamp 1670032574
transform 1 0 57132 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_614
timestamp 1670032574
transform 1 0 57592 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_97_617
timestamp 1670032574
transform 1 0 57868 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_623
timestamp 1670032574
transform 1 0 58420 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_3
timestamp 1670032574
transform 1 0 1380 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_9
timestamp 1670032574
transform 1 0 1932 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1670032574
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1670032574
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1670032574
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1670032574
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1670032574
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1670032574
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1670032574
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1670032574
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1670032574
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1670032574
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1670032574
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1670032574
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1670032574
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1670032574
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1670032574
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1670032574
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1670032574
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1670032574
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1670032574
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1670032574
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1670032574
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_209
timestamp 1670032574
transform 1 0 20332 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_217
timestamp 1670032574
transform 1 0 21068 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_98_224
timestamp 1670032574
transform 1 0 21712 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_232
timestamp 1670032574
transform 1 0 22448 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_235
timestamp 1670032574
transform 1 0 22724 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_247
timestamp 1670032574
transform 1 0 23828 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1670032574
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_253
timestamp 1670032574
transform 1 0 24380 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_261
timestamp 1670032574
transform 1 0 25116 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_265
timestamp 1670032574
transform 1 0 25484 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_274
timestamp 1670032574
transform 1 0 26312 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_286
timestamp 1670032574
transform 1 0 27416 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_292
timestamp 1670032574
transform 1 0 27968 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_299
timestamp 1670032574
transform 1 0 28612 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_303
timestamp 1670032574
transform 1 0 28980 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_306
timestamp 1670032574
transform 1 0 29256 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_309
timestamp 1670032574
transform 1 0 29532 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_319
timestamp 1670032574
transform 1 0 30452 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_325
timestamp 1670032574
transform 1 0 31004 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_337
timestamp 1670032574
transform 1 0 32108 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_98_353
timestamp 1670032574
transform 1 0 33580 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_361
timestamp 1670032574
transform 1 0 34316 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_98_365
timestamp 1670032574
transform 1 0 34684 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_375
timestamp 1670032574
transform 1 0 35604 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_381
timestamp 1670032574
transform 1 0 36156 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_389
timestamp 1670032574
transform 1 0 36892 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_397
timestamp 1670032574
transform 1 0 37628 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_402
timestamp 1670032574
transform 1 0 38088 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1670032574
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1670032574
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1670032574
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_433
timestamp 1670032574
transform 1 0 40940 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_98_447
timestamp 1670032574
transform 1 0 42228 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_455
timestamp 1670032574
transform 1 0 42964 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_98_466
timestamp 1670032574
transform 1 0 43976 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_474
timestamp 1670032574
transform 1 0 44712 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1670032574
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1670032574
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1670032574
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1670032574
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1670032574
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1670032574
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1670032574
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1670032574
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1670032574
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1670032574
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1670032574
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1670032574
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1670032574
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_601
timestamp 1670032574
transform 1 0 56396 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_607
timestamp 1670032574
transform 1 0 56948 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_610
timestamp 1670032574
transform 1 0 57224 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_616
timestamp 1670032574
transform 1 0 57776 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_623
timestamp 1670032574
transform 1 0 58420 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1670032574
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1670032574
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1670032574
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1670032574
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1670032574
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1670032574
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1670032574
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1670032574
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1670032574
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1670032574
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1670032574
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1670032574
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1670032574
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1670032574
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1670032574
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1670032574
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1670032574
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1670032574
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1670032574
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1670032574
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1670032574
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1670032574
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_222
timestamp 1670032574
transform 1 0 21528 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_225
timestamp 1670032574
transform 1 0 21804 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_232
timestamp 1670032574
transform 1 0 22448 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_240
timestamp 1670032574
transform 1 0 23184 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_249
timestamp 1670032574
transform 1 0 24012 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_257
timestamp 1670032574
transform 1 0 24748 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_266
timestamp 1670032574
transform 1 0 25576 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_278
timestamp 1670032574
transform 1 0 26680 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1670032574
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_293
timestamp 1670032574
transform 1 0 28060 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_303
timestamp 1670032574
transform 1 0 28980 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_311
timestamp 1670032574
transform 1 0 29716 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_321
timestamp 1670032574
transform 1 0 30636 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_99_333
timestamp 1670032574
transform 1 0 31740 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_99_337
timestamp 1670032574
transform 1 0 32108 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_343
timestamp 1670032574
transform 1 0 32660 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_352
timestamp 1670032574
transform 1 0 33488 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_364
timestamp 1670032574
transform 1 0 34592 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_378
timestamp 1670032574
transform 1 0 35880 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_390
timestamp 1670032574
transform 1 0 36984 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_393
timestamp 1670032574
transform 1 0 37260 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_401
timestamp 1670032574
transform 1 0 37996 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_411
timestamp 1670032574
transform 1 0 38916 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_422
timestamp 1670032574
transform 1 0 39928 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_434
timestamp 1670032574
transform 1 0 41032 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_444
timestamp 1670032574
transform 1 0 41952 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_449
timestamp 1670032574
transform 1 0 42412 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_457
timestamp 1670032574
transform 1 0 43148 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_466
timestamp 1670032574
transform 1 0 43976 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_478
timestamp 1670032574
transform 1 0 45080 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_490
timestamp 1670032574
transform 1 0 46184 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_502
timestamp 1670032574
transform 1 0 47288 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1670032574
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1670032574
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1670032574
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1670032574
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1670032574
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1670032574
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1670032574
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1670032574
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1670032574
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_599
timestamp 1670032574
transform 1 0 56212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_605
timestamp 1670032574
transform 1 0 56764 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_611
timestamp 1670032574
transform 1 0 57316 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1670032574
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_617
timestamp 1670032574
transform 1 0 57868 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1670032574
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_3
timestamp 1670032574
transform 1 0 1380 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_9
timestamp 1670032574
transform 1 0 1932 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_23
timestamp 1670032574
transform 1 0 3220 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1670032574
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_29
timestamp 1670032574
transform 1 0 3772 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_35
timestamp 1670032574
transform 1 0 4324 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_47
timestamp 1670032574
transform 1 0 5428 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_55
timestamp 1670032574
transform 1 0 6164 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_61
timestamp 1670032574
transform 1 0 6716 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_73
timestamp 1670032574
transform 1 0 7820 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_79
timestamp 1670032574
transform 1 0 8372 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_82
timestamp 1670032574
transform 1 0 8648 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_85
timestamp 1670032574
transform 1 0 8924 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_89
timestamp 1670032574
transform 1 0 9292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_101
timestamp 1670032574
transform 1 0 10396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_113
timestamp 1670032574
transform 1 0 11500 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_121
timestamp 1670032574
transform 1 0 12236 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_126
timestamp 1670032574
transform 1 0 12696 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_138
timestamp 1670032574
transform 1 0 13800 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_141
timestamp 1670032574
transform 1 0 14076 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_149
timestamp 1670032574
transform 1 0 14812 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_152
timestamp 1670032574
transform 1 0 15088 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_164
timestamp 1670032574
transform 1 0 16192 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_178
timestamp 1670032574
transform 1 0 17480 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_190
timestamp 1670032574
transform 1 0 18584 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_197
timestamp 1670032574
transform 1 0 19228 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_201
timestamp 1670032574
transform 1 0 19596 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_204
timestamp 1670032574
transform 1 0 19872 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_216
timestamp 1670032574
transform 1 0 20976 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_224
timestamp 1670032574
transform 1 0 21712 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_230
timestamp 1670032574
transform 1 0 22264 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_242
timestamp 1670032574
transform 1 0 23368 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_250
timestamp 1670032574
transform 1 0 24104 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_253
timestamp 1670032574
transform 1 0 24380 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_257
timestamp 1670032574
transform 1 0 24748 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_265
timestamp 1670032574
transform 1 0 25484 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_270
timestamp 1670032574
transform 1 0 25944 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_282
timestamp 1670032574
transform 1 0 27048 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_290
timestamp 1670032574
transform 1 0 27784 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_295
timestamp 1670032574
transform 1 0 28244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1670032574
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_309
timestamp 1670032574
transform 1 0 29532 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_317
timestamp 1670032574
transform 1 0 30268 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_329
timestamp 1670032574
transform 1 0 31372 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_339
timestamp 1670032574
transform 1 0 32292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_351
timestamp 1670032574
transform 1 0 33396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1670032574
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_365
timestamp 1670032574
transform 1 0 34684 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_371
timestamp 1670032574
transform 1 0 35236 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_374
timestamp 1670032574
transform 1 0 35512 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_382
timestamp 1670032574
transform 1 0 36248 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_386
timestamp 1670032574
transform 1 0 36616 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_398
timestamp 1670032574
transform 1 0 37720 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_402
timestamp 1670032574
transform 1 0 38088 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_405
timestamp 1670032574
transform 1 0 38364 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_416
timestamp 1670032574
transform 1 0 39376 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1670032574
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_433
timestamp 1670032574
transform 1 0 40940 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_438
timestamp 1670032574
transform 1 0 41400 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_450
timestamp 1670032574
transform 1 0 42504 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_458
timestamp 1670032574
transform 1 0 43240 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_468
timestamp 1670032574
transform 1 0 44160 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_477
timestamp 1670032574
transform 1 0 44988 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_481
timestamp 1670032574
transform 1 0 45356 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_493
timestamp 1670032574
transform 1 0 46460 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_507
timestamp 1670032574
transform 1 0 47748 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_519
timestamp 1670032574
transform 1 0 48852 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1670032574
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_533
timestamp 1670032574
transform 1 0 50140 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_537
timestamp 1670032574
transform 1 0 50508 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_549
timestamp 1670032574
transform 1 0 51612 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_555
timestamp 1670032574
transform 1 0 52164 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_567
timestamp 1670032574
transform 1 0 53268 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1670032574
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1670032574
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_589
timestamp 1670032574
transform 1 0 55292 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_593
timestamp 1670032574
transform 1 0 55660 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_596
timestamp 1670032574
transform 1 0 55936 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_602
timestamp 1670032574
transform 1 0 56488 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_609
timestamp 1670032574
transform 1 0 57132 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_616
timestamp 1670032574
transform 1 0 57776 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_623
timestamp 1670032574
transform 1 0 58420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_3
timestamp 1670032574
transform 1 0 1380 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_19
timestamp 1670032574
transform 1 0 2852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_26
timestamp 1670032574
transform 1 0 3496 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_29
timestamp 1670032574
transform 1 0 3772 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_38
timestamp 1670032574
transform 1 0 4600 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1670032574
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_57
timestamp 1670032574
transform 1 0 6348 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_64
timestamp 1670032574
transform 1 0 6992 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_82
timestamp 1670032574
transform 1 0 8648 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_85
timestamp 1670032574
transform 1 0 8924 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_90
timestamp 1670032574
transform 1 0 9384 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_96
timestamp 1670032574
transform 1 0 9936 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_103
timestamp 1670032574
transform 1 0 10580 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_107
timestamp 1670032574
transform 1 0 10948 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_110
timestamp 1670032574
transform 1 0 11224 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_113
timestamp 1670032574
transform 1 0 11500 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_118
timestamp 1670032574
transform 1 0 11960 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_101_129
timestamp 1670032574
transform 1 0 12972 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_135
timestamp 1670032574
transform 1 0 13524 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_138
timestamp 1670032574
transform 1 0 13800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_141
timestamp 1670032574
transform 1 0 14076 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_146
timestamp 1670032574
transform 1 0 14536 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_155
timestamp 1670032574
transform 1 0 15364 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_163
timestamp 1670032574
transform 1 0 16100 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_166
timestamp 1670032574
transform 1 0 16376 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_169
timestamp 1670032574
transform 1 0 16652 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_174
timestamp 1670032574
transform 1 0 17112 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_181
timestamp 1670032574
transform 1 0 17756 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_187
timestamp 1670032574
transform 1 0 18308 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_194
timestamp 1670032574
transform 1 0 18952 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_197
timestamp 1670032574
transform 1 0 19228 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_203
timestamp 1670032574
transform 1 0 19780 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_207
timestamp 1670032574
transform 1 0 20148 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_213
timestamp 1670032574
transform 1 0 20700 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_220
timestamp 1670032574
transform 1 0 21344 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_225
timestamp 1670032574
transform 1 0 21804 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_229
timestamp 1670032574
transform 1 0 22172 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_233
timestamp 1670032574
transform 1 0 22540 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_239
timestamp 1670032574
transform 1 0 23092 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_246
timestamp 1670032574
transform 1 0 23736 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_101_253
timestamp 1670032574
transform 1 0 24380 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_259
timestamp 1670032574
transform 1 0 24932 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_265
timestamp 1670032574
transform 1 0 25484 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_272
timestamp 1670032574
transform 1 0 26128 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_278
timestamp 1670032574
transform 1 0 26680 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_281
timestamp 1670032574
transform 1 0 26956 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_286
timestamp 1670032574
transform 1 0 27416 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_294
timestamp 1670032574
transform 1 0 28152 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_298
timestamp 1670032574
transform 1 0 28520 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_306
timestamp 1670032574
transform 1 0 29256 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_309
timestamp 1670032574
transform 1 0 29532 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_314
timestamp 1670032574
transform 1 0 29992 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_320
timestamp 1670032574
transform 1 0 30544 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_324
timestamp 1670032574
transform 1 0 30912 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_330
timestamp 1670032574
transform 1 0 31464 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_101_337
timestamp 1670032574
transform 1 0 32108 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_342
timestamp 1670032574
transform 1 0 32568 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_346
timestamp 1670032574
transform 1 0 32936 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_350
timestamp 1670032574
transform 1 0 33304 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_356
timestamp 1670032574
transform 1 0 33856 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_362
timestamp 1670032574
transform 1 0 34408 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_365
timestamp 1670032574
transform 1 0 34684 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_370
timestamp 1670032574
transform 1 0 35144 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_377
timestamp 1670032574
transform 1 0 35788 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_385
timestamp 1670032574
transform 1 0 36524 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1670032574
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_393
timestamp 1670032574
transform 1 0 37260 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_402
timestamp 1670032574
transform 1 0 38088 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_408
timestamp 1670032574
transform 1 0 38640 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_415
timestamp 1670032574
transform 1 0 39284 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_419
timestamp 1670032574
transform 1 0 39652 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_421
timestamp 1670032574
transform 1 0 39836 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_428
timestamp 1670032574
transform 1 0 40480 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_434
timestamp 1670032574
transform 1 0 41032 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1670032574
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1670032574
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_449
timestamp 1670032574
transform 1 0 42412 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_454
timestamp 1670032574
transform 1 0 42872 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_460
timestamp 1670032574
transform 1 0 43424 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_467
timestamp 1670032574
transform 1 0 44068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_473
timestamp 1670032574
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_477
timestamp 1670032574
transform 1 0 44988 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_482
timestamp 1670032574
transform 1 0 45448 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_493
timestamp 1670032574
transform 1 0 46460 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_499
timestamp 1670032574
transform 1 0 47012 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1670032574
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_505
timestamp 1670032574
transform 1 0 47564 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_510
timestamp 1670032574
transform 1 0 48024 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_519
timestamp 1670032574
transform 1 0 48852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_525
timestamp 1670032574
transform 1 0 49404 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_531
timestamp 1670032574
transform 1 0 49956 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1670032574
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_538
timestamp 1670032574
transform 1 0 50600 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_545
timestamp 1670032574
transform 1 0 51244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_551
timestamp 1670032574
transform 1 0 51796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_558
timestamp 1670032574
transform 1 0 52440 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_561
timestamp 1670032574
transform 1 0 52716 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_567
timestamp 1670032574
transform 1 0 53268 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_571
timestamp 1670032574
transform 1 0 53636 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_577
timestamp 1670032574
transform 1 0 54188 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_584
timestamp 1670032574
transform 1 0 54832 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_589
timestamp 1670032574
transform 1 0 55292 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_593
timestamp 1670032574
transform 1 0 55660 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_597
timestamp 1670032574
transform 1 0 56028 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_603
timestamp 1670032574
transform 1 0 56580 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_610
timestamp 1670032574
transform 1 0 57224 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_101_617
timestamp 1670032574
transform 1 0 57868 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_623
timestamp 1670032574
transform 1 0 58420 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1670032574
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1670032574
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1670032574
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1670032574
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1670032574
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1670032574
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1670032574
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1670032574
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1670032574
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1670032574
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1670032574
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1670032574
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1670032574
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1670032574
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1670032574
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1670032574
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1670032574
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1670032574
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1670032574
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1670032574
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1670032574
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1670032574
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1670032574
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1670032574
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1670032574
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1670032574
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1670032574
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1670032574
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1670032574
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1670032574
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1670032574
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1670032574
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1670032574
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1670032574
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1670032574
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1670032574
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1670032574
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1670032574
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1670032574
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1670032574
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1670032574
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1670032574
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1670032574
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1670032574
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1670032574
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1670032574
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1670032574
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1670032574
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1670032574
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1670032574
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1670032574
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1670032574
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1670032574
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1670032574
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1670032574
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1670032574
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1670032574
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1670032574
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1670032574
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1670032574
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1670032574
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1670032574
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1670032574
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1670032574
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1670032574
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1670032574
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1670032574
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1670032574
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1670032574
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1670032574
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1670032574
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1670032574
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1670032574
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1670032574
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1670032574
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1670032574
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1670032574
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1670032574
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1670032574
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1670032574
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1670032574
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1670032574
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1670032574
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1670032574
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1670032574
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1670032574
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1670032574
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1670032574
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1670032574
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1670032574
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1670032574
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1670032574
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1670032574
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1670032574
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1670032574
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1670032574
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1670032574
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1670032574
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1670032574
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1670032574
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1670032574
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1670032574
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1670032574
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1670032574
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1670032574
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1670032574
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1670032574
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1670032574
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1670032574
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1670032574
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1670032574
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1670032574
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1670032574
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1670032574
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1670032574
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1670032574
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1670032574
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1670032574
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1670032574
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1670032574
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1670032574
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1670032574
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1670032574
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1670032574
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1670032574
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1670032574
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1670032574
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1670032574
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1670032574
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1670032574
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1670032574
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1670032574
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1670032574
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1670032574
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1670032574
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1670032574
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1670032574
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1670032574
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1670032574
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1670032574
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1670032574
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1670032574
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1670032574
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1670032574
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1670032574
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1670032574
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1670032574
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1670032574
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1670032574
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1670032574
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1670032574
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1670032574
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1670032574
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1670032574
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1670032574
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1670032574
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1670032574
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1670032574
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1670032574
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1670032574
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1670032574
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1670032574
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1670032574
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1670032574
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1670032574
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1670032574
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1670032574
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1670032574
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1670032574
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1670032574
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1670032574
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1670032574
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1670032574
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1670032574
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1670032574
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1670032574
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1670032574
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1670032574
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1670032574
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1670032574
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1670032574
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1670032574
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1670032574
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1670032574
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1670032574
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1670032574
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1670032574
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1670032574
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1670032574
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1670032574
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1670032574
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1670032574
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1670032574
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1670032574
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1670032574
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1670032574
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1670032574
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1670032574
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1670032574
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1670032574
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1670032574
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1670032574
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1670032574
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1670032574
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1670032574
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1670032574
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1670032574
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1670032574
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1670032574
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1670032574
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1670032574
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1670032574
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1670032574
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1670032574
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1670032574
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1670032574
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1670032574
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1670032574
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1670032574
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1670032574
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1670032574
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1670032574
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1670032574
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1670032574
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1670032574
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1670032574
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1670032574
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1670032574
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1670032574
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1670032574
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1670032574
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1670032574
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1670032574
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1670032574
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1670032574
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1670032574
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1670032574
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1670032574
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1670032574
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1670032574
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1670032574
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1670032574
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1670032574
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1670032574
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1670032574
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1670032574
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1670032574
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1670032574
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1670032574
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1670032574
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1670032574
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1670032574
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1670032574
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1670032574
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1670032574
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1670032574
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1670032574
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1670032574
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1670032574
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1670032574
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1670032574
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1670032574
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1670032574
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1670032574
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1670032574
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1670032574
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1670032574
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1670032574
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1670032574
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1670032574
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1670032574
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1670032574
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1670032574
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1670032574
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1670032574
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1670032574
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1670032574
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1670032574
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1670032574
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1670032574
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1670032574
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1670032574
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1670032574
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1670032574
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1670032574
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1670032574
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1670032574
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1670032574
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1670032574
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1670032574
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1670032574
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1670032574
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1670032574
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1670032574
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1670032574
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1670032574
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1670032574
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1670032574
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1670032574
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1670032574
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1670032574
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1670032574
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1670032574
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1670032574
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1670032574
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1670032574
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1670032574
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1670032574
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1670032574
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1670032574
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1670032574
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1670032574
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1670032574
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1670032574
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1670032574
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1670032574
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1670032574
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1670032574
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1670032574
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1670032574
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1670032574
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1670032574
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1670032574
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1670032574
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1670032574
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1670032574
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1670032574
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1670032574
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1670032574
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1670032574
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1670032574
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1670032574
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1670032574
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1670032574
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1670032574
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1670032574
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1670032574
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1670032574
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1670032574
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1670032574
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1670032574
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1670032574
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1670032574
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1670032574
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1670032574
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1670032574
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1670032574
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1670032574
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1670032574
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1670032574
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1670032574
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1670032574
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1670032574
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1670032574
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1670032574
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1670032574
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1670032574
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1670032574
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1670032574
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1670032574
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1670032574
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1670032574
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1670032574
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1670032574
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1670032574
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1670032574
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1670032574
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1670032574
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1670032574
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1670032574
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1670032574
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1670032574
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1670032574
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1670032574
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1670032574
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1670032574
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1670032574
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1670032574
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1670032574
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1670032574
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1670032574
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1670032574
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1670032574
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1670032574
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1670032574
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1670032574
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1670032574
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1670032574
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1670032574
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1670032574
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1670032574
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1670032574
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1670032574
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1670032574
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1670032574
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1670032574
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1670032574
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1670032574
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1670032574
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1670032574
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1670032574
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1670032574
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1670032574
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1670032574
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1670032574
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1670032574
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1670032574
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1670032574
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1670032574
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1670032574
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1670032574
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1670032574
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1670032574
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1670032574
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1670032574
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1670032574
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1670032574
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1670032574
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1670032574
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1670032574
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1670032574
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1670032574
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1670032574
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1670032574
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1670032574
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1670032574
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1670032574
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1670032574
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1670032574
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1670032574
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1670032574
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1670032574
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1670032574
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1670032574
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1670032574
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1670032574
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1670032574
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1670032574
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1670032574
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1670032574
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1670032574
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1670032574
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1670032574
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1670032574
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1670032574
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1670032574
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1670032574
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1670032574
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1670032574
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1670032574
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1670032574
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1670032574
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1670032574
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1670032574
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1670032574
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1670032574
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1670032574
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1670032574
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1670032574
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1670032574
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1670032574
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1670032574
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1670032574
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1670032574
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1670032574
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1670032574
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1670032574
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1670032574
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1670032574
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1670032574
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1670032574
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1670032574
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1670032574
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1670032574
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1670032574
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1670032574
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1670032574
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1670032574
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1670032574
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1670032574
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1670032574
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1670032574
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1670032574
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1670032574
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1670032574
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1670032574
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1670032574
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1670032574
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1670032574
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1670032574
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1670032574
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1670032574
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1670032574
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1670032574
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1670032574
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1670032574
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1670032574
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1670032574
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1670032574
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1670032574
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1670032574
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1670032574
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1670032574
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1670032574
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1670032574
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1670032574
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1670032574
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1670032574
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1670032574
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1670032574
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1670032574
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1670032574
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1670032574
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1670032574
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1670032574
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1670032574
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1670032574
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1670032574
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1670032574
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1670032574
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1670032574
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1670032574
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1670032574
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1670032574
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1670032574
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1670032574
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1670032574
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1670032574
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1670032574
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1670032574
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1670032574
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1670032574
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1670032574
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1670032574
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1670032574
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1670032574
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1670032574
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1670032574
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1670032574
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1670032574
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1670032574
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1670032574
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1670032574
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1670032574
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1670032574
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1670032574
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1670032574
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1670032574
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1670032574
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1670032574
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1670032574
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1670032574
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1670032574
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1670032574
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1670032574
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1670032574
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1670032574
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1670032574
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1670032574
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1670032574
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1670032574
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1670032574
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1670032574
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1670032574
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1670032574
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1670032574
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1670032574
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1670032574
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1670032574
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1670032574
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1670032574
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1670032574
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1670032574
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1670032574
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1670032574
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1670032574
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1670032574
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1670032574
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1670032574
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1670032574
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1670032574
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1670032574
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1670032574
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1670032574
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1670032574
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1670032574
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1670032574
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1670032574
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1670032574
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1670032574
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1670032574
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1670032574
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1670032574
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1670032574
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1670032574
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1670032574
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1670032574
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1670032574
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1670032574
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1670032574
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1670032574
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1670032574
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1670032574
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1670032574
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1670032574
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1670032574
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1670032574
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1670032574
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1670032574
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1670032574
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1670032574
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1670032574
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1670032574
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1670032574
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1670032574
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1670032574
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1670032574
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1670032574
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1670032574
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1670032574
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1670032574
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1670032574
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1670032574
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1670032574
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1670032574
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1670032574
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1670032574
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1670032574
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1670032574
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1670032574
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1670032574
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1670032574
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1670032574
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1670032574
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1670032574
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1670032574
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1670032574
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1670032574
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1670032574
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1670032574
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1670032574
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1670032574
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1670032574
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1670032574
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1670032574
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1670032574
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1670032574
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1670032574
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1670032574
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1670032574
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1670032574
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1670032574
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1670032574
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1670032574
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1670032574
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1670032574
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1670032574
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1670032574
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1670032574
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1670032574
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1670032574
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1670032574
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1670032574
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1670032574
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1670032574
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1670032574
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1670032574
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1670032574
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1670032574
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1670032574
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1670032574
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1670032574
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1670032574
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1670032574
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1670032574
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1670032574
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1670032574
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1670032574
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1670032574
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1670032574
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1670032574
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1670032574
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1670032574
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1670032574
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1670032574
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1670032574
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1670032574
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1670032574
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1670032574
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1670032574
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1670032574
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1670032574
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1670032574
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1670032574
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1670032574
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1670032574
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1670032574
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1670032574
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1670032574
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1670032574
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1670032574
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1670032574
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1670032574
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1670032574
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1670032574
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1670032574
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1670032574
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1670032574
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1670032574
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1670032574
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1670032574
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1670032574
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1670032574
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1670032574
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1670032574
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1670032574
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1670032574
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1670032574
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1670032574
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1670032574
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1670032574
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1670032574
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1670032574
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1670032574
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1670032574
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1670032574
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1670032574
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1670032574
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1670032574
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1670032574
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1670032574
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1670032574
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1670032574
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1670032574
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1670032574
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1670032574
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1670032574
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1670032574
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1670032574
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1670032574
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1670032574
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1670032574
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1670032574
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1670032574
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1670032574
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1670032574
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1670032574
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1670032574
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1670032574
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1670032574
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1670032574
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1670032574
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1670032574
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1670032574
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1670032574
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1670032574
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1670032574
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1670032574
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1670032574
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1670032574
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1670032574
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1670032574
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1670032574
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1670032574
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1670032574
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1670032574
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1670032574
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1670032574
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1670032574
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1670032574
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1670032574
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1670032574
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1670032574
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1670032574
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1670032574
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1670032574
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1670032574
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1670032574
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1670032574
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1670032574
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1670032574
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1670032574
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1670032574
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1670032574
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1670032574
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1670032574
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1670032574
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1670032574
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1670032574
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1670032574
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1670032574
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1670032574
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1670032574
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1670032574
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1670032574
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1670032574
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1670032574
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1670032574
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1670032574
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1670032574
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1670032574
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1670032574
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1670032574
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1670032574
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1670032574
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1670032574
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1670032574
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1670032574
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1670032574
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1670032574
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1670032574
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1670032574
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1670032574
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1670032574
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1670032574
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1670032574
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1670032574
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1670032574
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1670032574
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1670032574
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1670032574
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1670032574
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1670032574
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1670032574
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1670032574
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1670032574
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1670032574
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1670032574
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1670032574
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1670032574
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1670032574
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1670032574
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1670032574
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1670032574
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1670032574
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1670032574
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1670032574
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1670032574
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1670032574
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1670032574
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1670032574
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1670032574
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1670032574
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1670032574
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1670032574
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1670032574
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1670032574
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1670032574
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1670032574
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1670032574
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1670032574
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1670032574
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1670032574
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1670032574
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1670032574
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1670032574
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1670032574
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1670032574
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1670032574
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1670032574
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1670032574
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1670032574
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1670032574
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1670032574
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1670032574
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1670032574
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1670032574
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1670032574
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1670032574
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1670032574
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1670032574
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1670032574
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1670032574
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1670032574
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1670032574
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1670032574
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1670032574
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1670032574
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1670032574
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1670032574
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1670032574
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1670032574
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1670032574
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1670032574
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1670032574
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1670032574
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1670032574
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1670032574
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1670032574
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1670032574
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1670032574
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1670032574
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1670032574
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1670032574
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1670032574
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1670032574
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1670032574
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1670032574
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1670032574
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1670032574
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1670032574
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1670032574
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1670032574
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1670032574
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1670032574
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1670032574
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1670032574
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1670032574
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1670032574
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1670032574
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1670032574
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1670032574
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1670032574
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1670032574
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1670032574
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1670032574
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1670032574
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1670032574
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1670032574
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1670032574
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1670032574
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1670032574
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1670032574
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1670032574
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1670032574
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1670032574
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1670032574
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1670032574
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1670032574
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1670032574
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1670032574
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1670032574
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1670032574
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1670032574
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1670032574
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1670032574
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1670032574
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1670032574
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1670032574
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1670032574
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1670032574
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1670032574
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1670032574
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1670032574
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1670032574
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1670032574
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1670032574
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1670032574
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1670032574
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1670032574
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1670032574
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1670032574
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1670032574
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1670032574
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1670032574
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1670032574
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1670032574
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1670032574
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1670032574
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1670032574
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1670032574
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1670032574
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1670032574
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1670032574
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1670032574
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1670032574
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1670032574
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1670032574
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1670032574
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1670032574
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1670032574
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1670032574
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1670032574
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1670032574
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1670032574
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1670032574
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1670032574
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1670032574
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1670032574
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1670032574
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1670032574
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1670032574
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1670032574
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1670032574
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1670032574
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1670032574
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1670032574
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1670032574
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1670032574
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1670032574
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1670032574
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1670032574
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1670032574
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1670032574
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1670032574
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1670032574
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1670032574
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1670032574
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1670032574
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1670032574
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1670032574
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1670032574
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1670032574
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1670032574
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1670032574
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1670032574
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1670032574
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1670032574
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1670032574
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1670032574
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1670032574
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1670032574
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1670032574
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1670032574
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1670032574
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1670032574
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1670032574
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1670032574
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1670032574
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1670032574
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1670032574
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1670032574
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1670032574
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1670032574
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1670032574
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1670032574
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1670032574
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1670032574
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1670032574
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1670032574
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1670032574
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1670032574
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1670032574
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1670032574
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1670032574
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1670032574
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1670032574
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1670032574
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1670032574
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1670032574
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1670032574
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1670032574
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1670032574
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1670032574
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1670032574
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1670032574
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1670032574
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1670032574
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1670032574
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1670032574
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1670032574
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1670032574
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1670032574
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1670032574
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1670032574
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1670032574
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1670032574
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1670032574
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1670032574
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1670032574
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1670032574
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1670032574
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1670032574
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1670032574
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1670032574
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1670032574
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1670032574
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1670032574
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1670032574
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1670032574
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1670032574
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1670032574
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1670032574
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1670032574
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1670032574
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1670032574
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1670032574
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1670032574
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1670032574
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1670032574
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1670032574
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1670032574
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1670032574
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1670032574
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1670032574
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1670032574
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1670032574
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1670032574
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1670032574
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1670032574
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1670032574
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1670032574
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1670032574
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1670032574
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1670032574
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1670032574
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1670032574
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1670032574
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1670032574
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1670032574
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1670032574
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1670032574
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1670032574
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1670032574
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1670032574
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1670032574
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1670032574
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1670032574
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1670032574
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1670032574
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1670032574
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1670032574
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1670032574
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1670032574
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1670032574
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1670032574
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1670032574
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1670032574
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1670032574
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1670032574
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1670032574
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1670032574
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1670032574
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1670032574
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1670032574
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1670032574
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1670032574
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1670032574
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1670032574
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1670032574
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1670032574
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1670032574
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1670032574
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1670032574
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1670032574
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1670032574
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1670032574
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1670032574
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1670032574
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1670032574
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1670032574
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1670032574
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1670032574
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1670032574
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1670032574
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1670032574
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1670032574
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1670032574
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1670032574
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1670032574
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1670032574
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1670032574
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1670032574
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1670032574
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1670032574
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1670032574
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1670032574
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1670032574
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1670032574
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1670032574
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1670032574
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1670032574
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1670032574
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1670032574
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1670032574
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1670032574
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1670032574
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1670032574
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1670032574
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1670032574
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1670032574
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1670032574
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1670032574
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1670032574
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1670032574
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1670032574
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1670032574
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1670032574
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1670032574
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1670032574
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1670032574
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1670032574
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1670032574
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1670032574
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1670032574
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1670032574
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1670032574
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1670032574
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1670032574
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1670032574
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1670032574
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1670032574
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1670032574
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1670032574
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1670032574
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1670032574
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1670032574
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1670032574
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1670032574
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1670032574
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1670032574
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1670032574
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1670032574
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1670032574
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1670032574
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1670032574
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1670032574
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1670032574
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1670032574
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1670032574
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1670032574
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1670032574
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1670032574
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1670032574
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1670032574
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1670032574
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1670032574
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1670032574
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1670032574
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1670032574
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1670032574
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1670032574
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1670032574
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1670032574
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1670032574
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1670032574
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1670032574
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1670032574
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1670032574
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1670032574
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1670032574
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1670032574
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1670032574
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1670032574
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1670032574
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1670032574
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1670032574
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1670032574
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1670032574
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1670032574
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1670032574
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1670032574
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1670032574
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1670032574
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1670032574
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1670032574
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1670032574
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1670032574
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1670032574
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1670032574
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1670032574
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1670032574
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1670032574
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1670032574
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1670032574
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1670032574
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1670032574
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1670032574
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1670032574
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1670032574
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1670032574
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1670032574
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1670032574
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1670032574
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1670032574
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1670032574
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1670032574
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1670032574
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1670032574
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1670032574
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1670032574
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1670032574
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1670032574
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1670032574
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1670032574
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1670032574
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1670032574
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1670032574
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1670032574
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1670032574
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1670032574
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1670032574
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1670032574
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1670032574
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1670032574
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1670032574
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1670032574
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1670032574
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1670032574
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1670032574
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1670032574
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1670032574
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1670032574
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1670032574
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1670032574
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1670032574
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1670032574
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1670032574
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1670032574
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1670032574
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1670032574
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1670032574
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1670032574
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1670032574
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1670032574
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1670032574
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1670032574
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1670032574
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1670032574
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1670032574
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1670032574
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1670032574
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1670032574
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1670032574
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1670032574
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1670032574
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1670032574
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1670032574
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1670032574
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1670032574
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1670032574
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1670032574
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1670032574
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1670032574
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1670032574
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1670032574
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1670032574
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1670032574
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1670032574
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1670032574
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1670032574
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1670032574
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1670032574
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1670032574
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1670032574
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1670032574
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1670032574
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1670032574
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1670032574
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1670032574
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1670032574
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1670032574
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1670032574
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1670032574
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1670032574
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1670032574
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1670032574
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _208_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 2760 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _209_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 3220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 1670032574
transform -1 0 13800 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1670032574
transform -1 0 15640 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 1670032574
transform 1 0 6532 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1670032574
transform -1 0 6808 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 1670032574
transform -1 0 11224 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1670032574
transform -1 0 11960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1670032574
transform 1 0 14720 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1670032574
transform 1 0 14536 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1670032574
transform 1 0 15916 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1670032574
transform 1 0 15824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1670032574
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1670032574
transform 1 0 18492 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1670032574
transform 1 0 19596 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1670032574
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1670032574
transform 1 0 22172 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1670032574
transform 1 0 22264 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _226_
timestamp 1670032574
transform 1 0 19688 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1670032574
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1670032574
transform 1 0 22080 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1670032574
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1670032574
transform 1 0 22448 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1670032574
transform 1 0 22448 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _232_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 38272 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _233_
timestamp 1670032574
transform 1 0 38456 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _234_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 33120 0 1 53312
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _235_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 32476 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _236_
timestamp 1670032574
transform -1 0 30912 0 1 53312
box -38 -48 1234 592
use sky130_fd_sc_hd__or3b_2  _237_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 28612 0 1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _238_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 30084 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _239_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 25576 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _240_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 32292 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _241_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 37536 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _242_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 36248 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _243_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 41124 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _244_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 40204 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _245_
timestamp 1670032574
transform 1 0 40112 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _246_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 41952 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _247_
timestamp 1670032574
transform -1 0 34960 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _248_
timestamp 1670032574
transform -1 0 33580 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _249_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 31832 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _250_
timestamp 1670032574
transform 1 0 25576 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _251_
timestamp 1670032574
transform 1 0 32292 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _252_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 21068 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _253_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 25944 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _254_
timestamp 1670032574
transform -1 0 44160 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _255_
timestamp 1670032574
transform 1 0 38272 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _256_
timestamp 1670032574
transform -1 0 33488 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _257_
timestamp 1670032574
transform 1 0 24564 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _258_
timestamp 1670032574
transform -1 0 24012 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _259_
timestamp 1670032574
transform 1 0 21988 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _260_
timestamp 1670032574
transform 1 0 23092 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _261_
timestamp 1670032574
transform -1 0 43976 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _262_
timestamp 1670032574
transform 1 0 37444 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _263_
timestamp 1670032574
transform -1 0 35880 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _264_
timestamp 1670032574
transform 1 0 24564 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _265_
timestamp 1670032574
transform -1 0 25392 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _266_
timestamp 1670032574
transform 1 0 21344 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _267_
timestamp 1670032574
transform 1 0 23552 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _268_
timestamp 1670032574
transform -1 0 44068 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _269_
timestamp 1670032574
transform 1 0 38732 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _270_
timestamp 1670032574
transform -1 0 35604 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _271_
timestamp 1670032574
transform 1 0 26128 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _272_
timestamp 1670032574
transform -1 0 27876 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _273_
timestamp 1670032574
transform 1 0 21068 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _274_
timestamp 1670032574
transform 1 0 26864 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _275_
timestamp 1670032574
transform -1 0 42228 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _276_
timestamp 1670032574
transform -1 0 39928 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _277_
timestamp 1670032574
transform -1 0 35880 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _278_
timestamp 1670032574
transform 1 0 28060 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _279_
timestamp 1670032574
transform 1 0 28244 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _280_
timestamp 1670032574
transform 1 0 21252 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _281_
timestamp 1670032574
transform 1 0 29716 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _282_
timestamp 1670032574
transform -1 0 43976 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _283_
timestamp 1670032574
transform 1 0 38456 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _284_
timestamp 1670032574
transform -1 0 36984 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _285_
timestamp 1670032574
transform -1 0 30268 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _286_
timestamp 1670032574
transform 1 0 29900 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _287_
timestamp 1670032574
transform 1 0 21252 0 1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _288_
timestamp 1670032574
transform 1 0 31004 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _289_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 56488 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _290_
timestamp 1670032574
transform 1 0 56120 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _291_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 56488 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1670032574
transform 1 0 58052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _293_
timestamp 1670032574
transform -1 0 57592 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1670032574
transform 1 0 56120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _295_
timestamp 1670032574
transform 1 0 56488 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1670032574
transform 1 0 58052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _297_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 58144 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1670032574
transform 1 0 40204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _299_
timestamp 1670032574
transform -1 0 57592 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1670032574
transform 1 0 55108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _301_
timestamp 1670032574
transform -1 0 58420 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1670032574
transform 1 0 58052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _303_
timestamp 1670032574
transform -1 0 58420 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1670032574
transform 1 0 44344 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _305_
timestamp 1670032574
transform -1 0 58420 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _306_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 58144 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _307_
timestamp 1670032574
transform -1 0 58328 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _308_
timestamp 1670032574
transform -1 0 57592 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_2  _309_
timestamp 1670032574
transform -1 0 58144 0 1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp 1670032574
transform 1 0 57316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _311_
timestamp 1670032574
transform -1 0 57592 0 -1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1670032574
transform 1 0 47932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _313_
timestamp 1670032574
transform -1 0 58420 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _314_
timestamp 1670032574
transform -1 0 55200 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _315_
timestamp 1670032574
transform -1 0 56304 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _316_
timestamp 1670032574
transform -1 0 54924 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _317_
timestamp 1670032574
transform -1 0 58236 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _318_
timestamp 1670032574
transform -1 0 52440 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_2  _319_
timestamp 1670032574
transform -1 0 58420 0 1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1670032574
transform 1 0 57316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _321_
timestamp 1670032574
transform -1 0 56120 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1670032574
transform 1 0 54464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _323_
timestamp 1670032574
transform -1 0 57132 0 1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1670032574
transform 1 0 55476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _325_
timestamp 1670032574
transform -1 0 58420 0 1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1670032574
transform 1 0 56764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _327_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 23000 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _328_
timestamp 1670032574
transform -1 0 19964 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1670032574
transform -1 0 5796 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1670032574
transform -1 0 6808 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1670032574
transform -1 0 6992 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1670032574
transform -1 0 7636 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1670032574
transform 1 0 8832 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp 1670032574
transform -1 0 8464 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1670032574
transform -1 0 8648 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1670032574
transform -1 0 9384 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1670032574
transform -1 0 7176 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1670032574
transform -1 0 7452 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1670032574
transform -1 0 9752 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1670032574
transform -1 0 10580 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1670032574
transform 1 0 9844 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1670032574
transform 1 0 9660 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1670032574
transform 1 0 12880 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1670032574
transform -1 0 12604 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1670032574
transform 1 0 12972 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1670032574
transform -1 0 12144 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1670032574
transform 1 0 17112 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1670032574
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1670032574
transform -1 0 19964 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp 1670032574
transform 1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1670032574
transform -1 0 20332 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1670032574
transform 1 0 20148 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1670032574
transform 1 0 19872 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1670032574
transform 1 0 19688 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1670032574
transform 1 0 19780 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1670032574
transform 1 0 19688 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1670032574
transform -1 0 22632 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1670032574
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1670032574
transform 1 0 22448 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _360_
timestamp 1670032574
transform 1 0 22356 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _361_
timestamp 1670032574
transform 1 0 22816 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _362_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 24104 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _363_
timestamp 1670032574
transform -1 0 21436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1670032574
transform -1 0 3036 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _365_
timestamp 1670032574
transform -1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _366_
timestamp 1670032574
transform -1 0 3036 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp 1670032574
transform -1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1670032574
transform -1 0 3036 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _369_
timestamp 1670032574
transform -1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1670032574
transform -1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _371_
timestamp 1670032574
transform -1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1670032574
transform -1 0 2944 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1670032574
transform -1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1670032574
transform -1 0 3036 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1670032574
transform -1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1670032574
transform -1 0 2944 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1670032574
transform -1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1670032574
transform 1 0 9108 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1670032574
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1670032574
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1670032574
transform 1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1670032574
transform 1 0 19320 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _383_
timestamp 1670032574
transform 1 0 18676 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1670032574
transform 1 0 19688 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1670032574
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1670032574
transform 1 0 19780 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _387_
timestamp 1670032574
transform 1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1670032574
transform 1 0 19872 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _389_
timestamp 1670032574
transform 1 0 19228 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1670032574
transform -1 0 20700 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _391_
timestamp 1670032574
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1670032574
transform 1 0 22540 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _393_
timestamp 1670032574
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1670032574
transform 1 0 22540 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _395_
timestamp 1670032574
transform 1 0 22172 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _396_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 23092 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  _397_
timestamp 1670032574
transform -1 0 20608 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1670032574
transform -1 0 2760 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1670032574
transform -1 0 2576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1670032574
transform -1 0 2760 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _401_
timestamp 1670032574
transform -1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1670032574
transform -1 0 2760 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1670032574
transform -1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1670032574
transform -1 0 2760 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp 1670032574
transform -1 0 2576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1670032574
transform -1 0 2760 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1670032574
transform -1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1670032574
transform -1 0 2852 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1670032574
transform -1 0 3496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1670032574
transform -1 0 2760 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1670032574
transform -1 0 2576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1670032574
transform 1 0 10120 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1670032574
transform 1 0 9476 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1670032574
transform 1 0 13800 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 1670032574
transform 1 0 13156 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _416_
timestamp 1670032574
transform 1 0 18768 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _417_
timestamp 1670032574
transform 1 0 18124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp 1670032574
transform 1 0 19780 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _419_
timestamp 1670032574
transform 1 0 19596 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp 1670032574
transform 1 0 19780 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _421_
timestamp 1670032574
transform 1 0 19688 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp 1670032574
transform 1 0 21712 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _423_
timestamp 1670032574
transform 1 0 21436 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _424_
timestamp 1670032574
transform 1 0 19872 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _425_
timestamp 1670032574
transform 1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _426_
timestamp 1670032574
transform 1 0 22448 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _427_
timestamp 1670032574
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _428_
timestamp 1670032574
transform 1 0 22540 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 1670032574
transform 1 0 22448 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _430_
timestamp 1670032574
transform -1 0 24012 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  _431_
timestamp 1670032574
transform -1 0 19688 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _432_
timestamp 1670032574
transform -1 0 2852 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _433_
timestamp 1670032574
transform -1 0 2668 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _434_
timestamp 1670032574
transform -1 0 4784 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1670032574
transform -1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1670032574
transform -1 0 3496 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _437_
timestamp 1670032574
transform -1 0 3956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _438_
timestamp 1670032574
transform -1 0 2760 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _439_
timestamp 1670032574
transform -1 0 2576 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _440_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 9292 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _441_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 7728 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _442_
timestamp 1670032574
transform 1 0 8096 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _443_
timestamp 1670032574
transform -1 0 15640 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _444_
timestamp 1670032574
transform -1 0 9752 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _445_
timestamp 1670032574
transform -1 0 12512 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _446_
timestamp 1670032574
transform 1 0 9108 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _447_
timestamp 1670032574
transform 1 0 12420 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _448_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform -1 0 12604 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _449_
timestamp 1670032574
transform 1 0 14996 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _450_
timestamp 1670032574
transform 1 0 15732 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _451_
timestamp 1670032574
transform 1 0 15088 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _452_
timestamp 1670032574
transform -1 0 17020 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _453_
timestamp 1670032574
transform 1 0 8740 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _454_
timestamp 1670032574
transform -1 0 9936 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _455_
timestamp 1670032574
transform 1 0 16836 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _456_
timestamp 1670032574
transform -1 0 6808 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _457_
timestamp 1670032574
transform -1 0 6072 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _458_
timestamp 1670032574
transform -1 0 9844 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _459_
timestamp 1670032574
transform -1 0 7452 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _460_
timestamp 1670032574
transform -1 0 5888 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _461_
timestamp 1670032574
transform -1 0 6992 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _462_
timestamp 1670032574
transform -1 0 6716 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _463_
timestamp 1670032574
transform 1 0 8004 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _464_
timestamp 1670032574
transform -1 0 11960 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1670032574
transform -1 0 13524 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 1670032574
transform -1 0 18676 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _467_
timestamp 1670032574
transform -1 0 13708 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _468_
timestamp 1670032574
transform -1 0 18584 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 1670032574
transform 1 0 9568 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _470_
timestamp 1670032574
transform -1 0 18216 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _471_
timestamp 1670032574
transform -1 0 14444 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1670032574
transform -1 0 6164 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _473_
timestamp 1670032574
transform -1 0 7912 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _474_
timestamp 1670032574
transform -1 0 6072 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _475_
timestamp 1670032574
transform -1 0 6164 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1670032574
transform -1 0 6256 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1670032574
transform -1 0 5980 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 1670032574
transform -1 0 6072 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _479_
timestamp 1670032574
transform 1 0 9108 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _480_
timestamp 1670032574
transform 1 0 12880 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _481_
timestamp 1670032574
transform 1 0 15364 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _482_
timestamp 1670032574
transform -1 0 13800 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _483_
timestamp 1670032574
transform -1 0 18032 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1670032574
transform -1 0 12696 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _485_
timestamp 1670032574
transform -1 0 18124 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _486_
timestamp 1670032574
transform 1 0 16836 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _487_
timestamp 1670032574
transform -1 0 16284 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1670032574
transform -1 0 5888 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1670032574
transform -1 0 10212 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1670032574
transform -1 0 6072 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 1670032574
transform -1 0 6716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 1670032574
transform -1 0 6624 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 1670032574
transform 1 0 15272 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1670032574
transform 1 0 7176 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1670032574
transform -1 0 13800 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _496_
timestamp 1670032574
transform -1 0 12328 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _497_
timestamp 1670032574
transform -1 0 13708 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _498_
timestamp 1670032574
transform 1 0 15364 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _499_
timestamp 1670032574
transform 1 0 15364 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _500_
timestamp 1670032574
transform -1 0 15640 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _501_
timestamp 1670032574
transform -1 0 13064 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _502_
timestamp 1670032574
transform -1 0 15916 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _503_
timestamp 1670032574
transform -1 0 13800 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1670032574
transform -1 0 57684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_reg_wr_i pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 11684 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_reg_wr_i
timestamp 1670032574
transform -1 0 9660 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_reg_wr_i
timestamp 1670032574
transform -1 0 9660 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_reg_wr_i
timestamp 1670032574
transform 1 0 12972 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_reg_wr_i
timestamp 1670032574
transform 1 0 12972 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_reg_wr_i
timestamp 1670032574
transform -1 0 9660 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_reg_wr_i
timestamp 1670032574
transform -1 0 9660 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_reg_wr_i
timestamp 1670032574
transform 1 0 12972 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_reg_wr_i
timestamp 1670032574
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout235
timestamp 1670032574
transform -1 0 7084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout236
timestamp 1670032574
transform 1 0 6532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout237
timestamp 1670032574
transform 1 0 14260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout238 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 12144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout239
timestamp 1670032574
transform -1 0 5980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout240
timestamp 1670032574
transform 1 0 5612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout241
timestamp 1670032574
transform -1 0 12236 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout242
timestamp 1670032574
transform -1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout243
timestamp 1670032574
transform 1 0 6532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1670032574
transform -1 0 56764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1670032574
transform 1 0 1932 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1670032574
transform -1 0 3496 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1670032574
transform -1 0 4600 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1670032574
transform -1 0 6072 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1670032574
transform -1 0 6992 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1670032574
transform -1 0 8648 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1670032574
transform -1 0 9384 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1670032574
transform -1 0 10580 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1670032574
transform -1 0 11960 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1670032574
transform -1 0 12972 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1670032574
transform -1 0 14536 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1670032574
transform -1 0 15364 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1670032574
transform -1 0 17112 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1670032574
transform -1 0 17756 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1670032574
transform -1 0 18952 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1670032574
transform -1 0 20148 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1670032574
transform -1 0 21344 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1670032574
transform -1 0 22540 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1670032574
transform -1 0 23736 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1670032574
transform -1 0 24932 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1670032574
transform 1 0 25852 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1670032574
transform 1 0 27140 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1670032574
transform -1 0 28520 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1670032574
transform 1 0 29716 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1670032574
transform -1 0 30912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1670032574
transform -1 0 32568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1670032574
transform -1 0 33304 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1670032574
transform -1 0 35144 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1670032574
transform 1 0 35512 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1670032574
transform 1 0 36616 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1670032574
transform 1 0 37812 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1670032574
transform 1 0 39008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1670032574
transform 1 0 40204 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1670032574
transform 1 0 41400 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1670032574
transform 1 0 42596 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1670032574
transform 1 0 43792 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1670032574
transform 1 0 45172 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1670032574
transform 1 0 46184 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1670032574
transform 1 0 47748 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1670032574
transform 1 0 48576 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1670032574
transform 1 0 50324 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1670032574
transform 1 0 50968 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1670032574
transform 1 0 52164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1670032574
transform 1 0 53360 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1670032574
transform 1 0 54556 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1670032574
transform 1 0 55752 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1670032574
transform 1 0 56948 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1670032574
transform 1 0 58144 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input50
timestamp 1670032574
transform 1 0 24564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input51
timestamp 1670032574
transform 1 0 25576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input52 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 27140 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  input53
timestamp 1670032574
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1670032574
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1670032574
transform -1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1670032574
transform 1 0 17848 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1670032574
transform 1 0 19044 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1670032574
transform 1 0 20056 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1670032574
transform 1 0 21160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1670032574
transform -1 0 22540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1670032574
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1670032574
transform -1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1670032574
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1670032574
transform -1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1670032574
transform -1 0 11224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input66
timestamp 1670032574
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1670032574
transform -1 0 13800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1670032574
transform -1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1670032574
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1670032574
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1670032574
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1670032574
transform 1 0 56672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1670032574
transform -1 0 56304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1670032574
transform 1 0 57316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1670032574
transform 1 0 57500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1670032574
transform 1 0 58144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1670032574
transform 1 0 58144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1670032574
transform 1 0 58144 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1670032574
transform 1 0 58144 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1670032574
transform 1 0 58144 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1670032574
transform 1 0 58144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1670032574
transform 1 0 58144 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1670032574
transform 1 0 58144 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1670032574
transform 1 0 58144 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1670032574
transform 1 0 58144 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1670032574
transform 1 0 57316 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1670032574
transform 1 0 58144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1670032574
transform 1 0 58144 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1670032574
transform 1 0 58144 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1670032574
transform 1 0 58144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1670032574
transform 1 0 58144 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1670032574
transform 1 0 58144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1670032574
transform 1 0 58144 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1670032574
transform 1 0 58144 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1670032574
transform -1 0 58420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1670032574
transform -1 0 58420 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1670032574
transform 1 0 58144 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1670032574
transform 1 0 58144 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1670032574
transform -1 0 58420 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1670032574
transform 1 0 58144 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1670032574
transform 1 0 58144 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1670032574
transform 1 0 58144 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1670032574
transform -1 0 58420 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1670032574
transform 1 0 58144 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1670032574
transform 1 0 58144 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1670032574
transform 1 0 58144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1670032574
transform 1 0 58144 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1670032574
transform 1 0 58144 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1670032574
transform 1 0 58144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1670032574
transform 1 0 58144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1670032574
transform 1 0 58144 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1670032574
transform 1 0 58144 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1670032574
transform 1 0 58144 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1670032574
transform 1 0 58144 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1670032574
transform 1 0 58144 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1670032574
transform 1 0 58144 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1670032574
transform 1 0 58144 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1670032574
transform 1 0 58144 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1670032574
transform 1 0 58144 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1670032574
transform 1 0 58144 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1670032574
transform 1 0 58144 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1670032574
transform 1 0 58144 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1670032574
transform 1 0 58144 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1670032574
transform 1 0 58144 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1670032574
transform 1 0 58144 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1670032574
transform 1 0 58144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1670032574
transform 1 0 58144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1670032574
transform 1 0 58144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1670032574
transform 1 0 58144 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1670032574
transform 1 0 58144 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1670032574
transform 1 0 58144 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1670032574
transform 1 0 58144 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1670032574
transform 1 0 58144 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1670032574
transform -1 0 57776 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1670032574
transform 1 0 58144 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1670032574
transform 1 0 58144 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1670032574
transform 1 0 58144 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input138
timestamp 1670032574
transform 1 0 58144 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1670032574
transform 1 0 58144 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1670032574
transform 1 0 58144 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1670032574
transform 1 0 58144 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1670032574
transform 1 0 58144 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1670032574
transform 1 0 56856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input144 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1670032574
transform 1 0 34868 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input145
timestamp 1670032574
transform 1 0 36064 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1670032574
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1670032574
transform 1 0 27784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1670032574
transform 1 0 28888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1670032574
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1670032574
transform 1 0 31096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1670032574
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1670032574
transform 1 0 33304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1670032574
transform -1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1670032574
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1670032574
transform -1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1670032574
transform -1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1670032574
transform -1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1670032574
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1670032574
transform -1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1670032574
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1670032574
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1670032574
transform -1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1670032574
transform -1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1670032574
transform -1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1670032574
transform -1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1670032574
transform -1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1670032574
transform -1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1670032574
transform -1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1670032574
transform -1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1670032574
transform -1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1670032574
transform -1 0 1932 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1670032574
transform -1 0 1932 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1670032574
transform -1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1670032574
transform -1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1670032574
transform -1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1670032574
transform -1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1670032574
transform -1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1670032574
transform -1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1670032574
transform -1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1670032574
transform -1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1670032574
transform -1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1670032574
transform -1 0 1932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1670032574
transform -1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1670032574
transform -1 0 1932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1670032574
transform -1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1670032574
transform -1 0 1932 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1670032574
transform -1 0 1932 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1670032574
transform -1 0 1932 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1670032574
transform -1 0 1932 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1670032574
transform -1 0 1932 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1670032574
transform -1 0 1932 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1670032574
transform -1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1670032574
transform -1 0 1932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1670032574
transform -1 0 1932 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1670032574
transform -1 0 1932 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1670032574
transform -1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1670032574
transform -1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1670032574
transform -1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1670032574
transform -1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1670032574
transform -1 0 1932 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1670032574
transform -1 0 1932 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1670032574
transform -1 0 1932 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1670032574
transform -1 0 1932 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1670032574
transform -1 0 1932 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1670032574
transform -1 0 1932 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1670032574
transform -1 0 1932 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1670032574
transform -1 0 1932 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1670032574
transform -1 0 1932 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1670032574
transform -1 0 1932 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1670032574
transform -1 0 1932 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1670032574
transform -1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1670032574
transform -1 0 1932 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1670032574
transform -1 0 1932 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1670032574
transform -1 0 1932 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1670032574
transform -1 0 1932 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1670032574
transform -1 0 1932 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1670032574
transform -1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1670032574
transform -1 0 38548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1670032574
transform -1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1670032574
transform -1 0 40388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1670032574
transform -1 0 41400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1670032574
transform -1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1670032574
transform -1 0 43700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1670032574
transform -1 0 54648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1670032574
transform -1 0 55844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1670032574
transform -1 0 44712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1670032574
transform -1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1670032574
transform -1 0 46920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1670032574
transform -1 0 48116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1670032574
transform -1 0 49128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1670032574
transform -1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1670032574
transform -1 0 51428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1670032574
transform -1 0 52440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1670032574
transform -1 0 53544 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 56414 0 56470 800 0 FreeSans 224 90 0 0 loopback_i
port 0 nsew signal input
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 loopback_o
port 1 nsew signal tristate
flabel metal2 s 1858 59200 1914 60000 0 FreeSans 224 90 0 0 mux0_i[0]
port 2 nsew signal input
flabel metal2 s 3054 59200 3110 60000 0 FreeSans 224 90 0 0 mux0_i[1]
port 3 nsew signal input
flabel metal2 s 4250 59200 4306 60000 0 FreeSans 224 90 0 0 mux0_i[2]
port 4 nsew signal input
flabel metal2 s 5446 59200 5502 60000 0 FreeSans 224 90 0 0 mux0_i[3]
port 5 nsew signal input
flabel metal2 s 6642 59200 6698 60000 0 FreeSans 224 90 0 0 mux0_i[4]
port 6 nsew signal input
flabel metal2 s 7838 59200 7894 60000 0 FreeSans 224 90 0 0 mux0_i[5]
port 7 nsew signal input
flabel metal2 s 9034 59200 9090 60000 0 FreeSans 224 90 0 0 mux1_i[0]
port 8 nsew signal input
flabel metal2 s 10230 59200 10286 60000 0 FreeSans 224 90 0 0 mux1_i[1]
port 9 nsew signal input
flabel metal2 s 11426 59200 11482 60000 0 FreeSans 224 90 0 0 mux1_i[2]
port 10 nsew signal input
flabel metal2 s 12622 59200 12678 60000 0 FreeSans 224 90 0 0 mux1_i[3]
port 11 nsew signal input
flabel metal2 s 13818 59200 13874 60000 0 FreeSans 224 90 0 0 mux1_i[4]
port 12 nsew signal input
flabel metal2 s 15014 59200 15070 60000 0 FreeSans 224 90 0 0 mux1_i[5]
port 13 nsew signal input
flabel metal2 s 16210 59200 16266 60000 0 FreeSans 224 90 0 0 mux2_i[0]
port 14 nsew signal input
flabel metal2 s 17406 59200 17462 60000 0 FreeSans 224 90 0 0 mux2_i[1]
port 15 nsew signal input
flabel metal2 s 18602 59200 18658 60000 0 FreeSans 224 90 0 0 mux2_i[2]
port 16 nsew signal input
flabel metal2 s 19798 59200 19854 60000 0 FreeSans 224 90 0 0 mux2_i[3]
port 17 nsew signal input
flabel metal2 s 20994 59200 21050 60000 0 FreeSans 224 90 0 0 mux2_i[4]
port 18 nsew signal input
flabel metal2 s 22190 59200 22246 60000 0 FreeSans 224 90 0 0 mux2_i[5]
port 19 nsew signal input
flabel metal2 s 23386 59200 23442 60000 0 FreeSans 224 90 0 0 mux3_i[0]
port 20 nsew signal input
flabel metal2 s 24582 59200 24638 60000 0 FreeSans 224 90 0 0 mux3_i[1]
port 21 nsew signal input
flabel metal2 s 25778 59200 25834 60000 0 FreeSans 224 90 0 0 mux3_i[2]
port 22 nsew signal input
flabel metal2 s 26974 59200 27030 60000 0 FreeSans 224 90 0 0 mux3_i[3]
port 23 nsew signal input
flabel metal2 s 28170 59200 28226 60000 0 FreeSans 224 90 0 0 mux3_i[4]
port 24 nsew signal input
flabel metal2 s 29366 59200 29422 60000 0 FreeSans 224 90 0 0 mux3_i[5]
port 25 nsew signal input
flabel metal2 s 30562 59200 30618 60000 0 FreeSans 224 90 0 0 mux4_i[0]
port 26 nsew signal input
flabel metal2 s 31758 59200 31814 60000 0 FreeSans 224 90 0 0 mux4_i[1]
port 27 nsew signal input
flabel metal2 s 32954 59200 33010 60000 0 FreeSans 224 90 0 0 mux4_i[2]
port 28 nsew signal input
flabel metal2 s 34150 59200 34206 60000 0 FreeSans 224 90 0 0 mux4_i[3]
port 29 nsew signal input
flabel metal2 s 35346 59200 35402 60000 0 FreeSans 224 90 0 0 mux4_i[4]
port 30 nsew signal input
flabel metal2 s 36542 59200 36598 60000 0 FreeSans 224 90 0 0 mux4_i[5]
port 31 nsew signal input
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 mux5_i[0]
port 32 nsew signal input
flabel metal2 s 38934 59200 38990 60000 0 FreeSans 224 90 0 0 mux5_i[1]
port 33 nsew signal input
flabel metal2 s 40130 59200 40186 60000 0 FreeSans 224 90 0 0 mux5_i[2]
port 34 nsew signal input
flabel metal2 s 41326 59200 41382 60000 0 FreeSans 224 90 0 0 mux5_i[3]
port 35 nsew signal input
flabel metal2 s 42522 59200 42578 60000 0 FreeSans 224 90 0 0 mux5_i[4]
port 36 nsew signal input
flabel metal2 s 43718 59200 43774 60000 0 FreeSans 224 90 0 0 mux5_i[5]
port 37 nsew signal input
flabel metal2 s 44914 59200 44970 60000 0 FreeSans 224 90 0 0 mux6_i[0]
port 38 nsew signal input
flabel metal2 s 46110 59200 46166 60000 0 FreeSans 224 90 0 0 mux6_i[1]
port 39 nsew signal input
flabel metal2 s 47306 59200 47362 60000 0 FreeSans 224 90 0 0 mux6_i[2]
port 40 nsew signal input
flabel metal2 s 48502 59200 48558 60000 0 FreeSans 224 90 0 0 mux6_i[3]
port 41 nsew signal input
flabel metal2 s 49698 59200 49754 60000 0 FreeSans 224 90 0 0 mux6_i[4]
port 42 nsew signal input
flabel metal2 s 50894 59200 50950 60000 0 FreeSans 224 90 0 0 mux6_i[5]
port 43 nsew signal input
flabel metal2 s 52090 59200 52146 60000 0 FreeSans 224 90 0 0 mux7_i[0]
port 44 nsew signal input
flabel metal2 s 53286 59200 53342 60000 0 FreeSans 224 90 0 0 mux7_i[1]
port 45 nsew signal input
flabel metal2 s 54482 59200 54538 60000 0 FreeSans 224 90 0 0 mux7_i[2]
port 46 nsew signal input
flabel metal2 s 55678 59200 55734 60000 0 FreeSans 224 90 0 0 mux7_i[3]
port 47 nsew signal input
flabel metal2 s 56874 59200 56930 60000 0 FreeSans 224 90 0 0 mux7_i[4]
port 48 nsew signal input
flabel metal2 s 58070 59200 58126 60000 0 FreeSans 224 90 0 0 mux7_i[5]
port 49 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 mux_adr_i[0]
port 50 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 mux_adr_i[1]
port 51 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 mux_adr_i[2]
port 52 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 mux_o[0]
port 53 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 mux_o[1]
port 54 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 mux_o[2]
port 55 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 mux_o[3]
port 56 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 mux_o[4]
port 57 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 mux_o[5]
port 58 nsew signal tristate
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 reg0_o[0]
port 59 nsew signal tristate
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 reg0_o[10]
port 60 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 reg0_o[11]
port 61 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 reg0_o[12]
port 62 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 reg0_o[13]
port 63 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 reg0_o[14]
port 64 nsew signal tristate
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 reg0_o[15]
port 65 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 reg0_o[1]
port 66 nsew signal tristate
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 reg0_o[2]
port 67 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 reg0_o[3]
port 68 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 reg0_o[4]
port 69 nsew signal tristate
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 reg0_o[5]
port 70 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 reg0_o[6]
port 71 nsew signal tristate
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 reg0_o[7]
port 72 nsew signal tristate
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 reg0_o[8]
port 73 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 reg0_o[9]
port 74 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 reg1_o[0]
port 75 nsew signal tristate
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 reg1_o[10]
port 76 nsew signal tristate
flabel metal3 s 0 26256 800 26376 0 FreeSans 480 0 0 0 reg1_o[11]
port 77 nsew signal tristate
flabel metal3 s 0 27072 800 27192 0 FreeSans 480 0 0 0 reg1_o[12]
port 78 nsew signal tristate
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 reg1_o[13]
port 79 nsew signal tristate
flabel metal3 s 0 28704 800 28824 0 FreeSans 480 0 0 0 reg1_o[14]
port 80 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 reg1_o[15]
port 81 nsew signal tristate
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 reg1_o[1]
port 82 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 reg1_o[2]
port 83 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 reg1_o[3]
port 84 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 reg1_o[4]
port 85 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 reg1_o[5]
port 86 nsew signal tristate
flabel metal3 s 0 22176 800 22296 0 FreeSans 480 0 0 0 reg1_o[6]
port 87 nsew signal tristate
flabel metal3 s 0 22992 800 23112 0 FreeSans 480 0 0 0 reg1_o[7]
port 88 nsew signal tristate
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 reg1_o[8]
port 89 nsew signal tristate
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 reg1_o[9]
port 90 nsew signal tristate
flabel metal3 s 0 30336 800 30456 0 FreeSans 480 0 0 0 reg2_o[0]
port 91 nsew signal tristate
flabel metal3 s 0 38496 800 38616 0 FreeSans 480 0 0 0 reg2_o[10]
port 92 nsew signal tristate
flabel metal3 s 0 39312 800 39432 0 FreeSans 480 0 0 0 reg2_o[11]
port 93 nsew signal tristate
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 reg2_o[12]
port 94 nsew signal tristate
flabel metal3 s 0 40944 800 41064 0 FreeSans 480 0 0 0 reg2_o[13]
port 95 nsew signal tristate
flabel metal3 s 0 41760 800 41880 0 FreeSans 480 0 0 0 reg2_o[14]
port 96 nsew signal tristate
flabel metal3 s 0 42576 800 42696 0 FreeSans 480 0 0 0 reg2_o[15]
port 97 nsew signal tristate
flabel metal3 s 0 31152 800 31272 0 FreeSans 480 0 0 0 reg2_o[1]
port 98 nsew signal tristate
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 reg2_o[2]
port 99 nsew signal tristate
flabel metal3 s 0 32784 800 32904 0 FreeSans 480 0 0 0 reg2_o[3]
port 100 nsew signal tristate
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 reg2_o[4]
port 101 nsew signal tristate
flabel metal3 s 0 34416 800 34536 0 FreeSans 480 0 0 0 reg2_o[5]
port 102 nsew signal tristate
flabel metal3 s 0 35232 800 35352 0 FreeSans 480 0 0 0 reg2_o[6]
port 103 nsew signal tristate
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 reg2_o[7]
port 104 nsew signal tristate
flabel metal3 s 0 36864 800 36984 0 FreeSans 480 0 0 0 reg2_o[8]
port 105 nsew signal tristate
flabel metal3 s 0 37680 800 37800 0 FreeSans 480 0 0 0 reg2_o[9]
port 106 nsew signal tristate
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 reg3_o[0]
port 107 nsew signal tristate
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 reg3_o[10]
port 108 nsew signal tristate
flabel metal3 s 0 52368 800 52488 0 FreeSans 480 0 0 0 reg3_o[11]
port 109 nsew signal tristate
flabel metal3 s 0 53184 800 53304 0 FreeSans 480 0 0 0 reg3_o[12]
port 110 nsew signal tristate
flabel metal3 s 0 54000 800 54120 0 FreeSans 480 0 0 0 reg3_o[13]
port 111 nsew signal tristate
flabel metal3 s 0 54816 800 54936 0 FreeSans 480 0 0 0 reg3_o[14]
port 112 nsew signal tristate
flabel metal3 s 0 55632 800 55752 0 FreeSans 480 0 0 0 reg3_o[15]
port 113 nsew signal tristate
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 reg3_o[1]
port 114 nsew signal tristate
flabel metal3 s 0 45024 800 45144 0 FreeSans 480 0 0 0 reg3_o[2]
port 115 nsew signal tristate
flabel metal3 s 0 45840 800 45960 0 FreeSans 480 0 0 0 reg3_o[3]
port 116 nsew signal tristate
flabel metal3 s 0 46656 800 46776 0 FreeSans 480 0 0 0 reg3_o[4]
port 117 nsew signal tristate
flabel metal3 s 0 47472 800 47592 0 FreeSans 480 0 0 0 reg3_o[5]
port 118 nsew signal tristate
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 reg3_o[6]
port 119 nsew signal tristate
flabel metal3 s 0 49104 800 49224 0 FreeSans 480 0 0 0 reg3_o[7]
port 120 nsew signal tristate
flabel metal3 s 0 49920 800 50040 0 FreeSans 480 0 0 0 reg3_o[8]
port 121 nsew signal tristate
flabel metal3 s 0 50736 800 50856 0 FreeSans 480 0 0 0 reg3_o[9]
port 122 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 reg_adr_i[0]
port 123 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 reg_adr_i[1]
port 124 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 reg_dat_i[0]
port 125 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 reg_dat_i[10]
port 126 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 reg_dat_i[11]
port 127 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 reg_dat_i[12]
port 128 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 reg_dat_i[13]
port 129 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 reg_dat_i[14]
port 130 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 reg_dat_i[15]
port 131 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 reg_dat_i[1]
port 132 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 reg_dat_i[2]
port 133 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 reg_dat_i[3]
port 134 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 reg_dat_i[4]
port 135 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 reg_dat_i[5]
port 136 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 reg_dat_i[6]
port 137 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 reg_dat_i[7]
port 138 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 reg_dat_i[8]
port 139 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 reg_dat_i[9]
port 140 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 reg_wr_i
port 141 nsew signal input
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 rst_n_i
port 142 nsew signal input
flabel metal3 s 59200 960 60000 1080 0 FreeSans 480 0 0 0 temp0_dac_i[0]
port 143 nsew signal input
flabel metal3 s 59200 1776 60000 1896 0 FreeSans 480 0 0 0 temp0_dac_i[1]
port 144 nsew signal input
flabel metal3 s 59200 2592 60000 2712 0 FreeSans 480 0 0 0 temp0_dac_i[2]
port 145 nsew signal input
flabel metal3 s 59200 3408 60000 3528 0 FreeSans 480 0 0 0 temp0_dac_i[3]
port 146 nsew signal input
flabel metal3 s 59200 4224 60000 4344 0 FreeSans 480 0 0 0 temp0_dac_i[4]
port 147 nsew signal input
flabel metal3 s 59200 5040 60000 5160 0 FreeSans 480 0 0 0 temp0_dac_i[5]
port 148 nsew signal input
flabel metal3 s 59200 20544 60000 20664 0 FreeSans 480 0 0 0 temp0_ticks_i[0]
port 149 nsew signal input
flabel metal3 s 59200 28704 60000 28824 0 FreeSans 480 0 0 0 temp0_ticks_i[10]
port 150 nsew signal input
flabel metal3 s 59200 29520 60000 29640 0 FreeSans 480 0 0 0 temp0_ticks_i[11]
port 151 nsew signal input
flabel metal3 s 59200 21360 60000 21480 0 FreeSans 480 0 0 0 temp0_ticks_i[1]
port 152 nsew signal input
flabel metal3 s 59200 22176 60000 22296 0 FreeSans 480 0 0 0 temp0_ticks_i[2]
port 153 nsew signal input
flabel metal3 s 59200 22992 60000 23112 0 FreeSans 480 0 0 0 temp0_ticks_i[3]
port 154 nsew signal input
flabel metal3 s 59200 23808 60000 23928 0 FreeSans 480 0 0 0 temp0_ticks_i[4]
port 155 nsew signal input
flabel metal3 s 59200 24624 60000 24744 0 FreeSans 480 0 0 0 temp0_ticks_i[5]
port 156 nsew signal input
flabel metal3 s 59200 25440 60000 25560 0 FreeSans 480 0 0 0 temp0_ticks_i[6]
port 157 nsew signal input
flabel metal3 s 59200 26256 60000 26376 0 FreeSans 480 0 0 0 temp0_ticks_i[7]
port 158 nsew signal input
flabel metal3 s 59200 27072 60000 27192 0 FreeSans 480 0 0 0 temp0_ticks_i[8]
port 159 nsew signal input
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 temp0_ticks_i[9]
port 160 nsew signal input
flabel metal3 s 59200 5856 60000 5976 0 FreeSans 480 0 0 0 temp1_dac_i[0]
port 161 nsew signal input
flabel metal3 s 59200 6672 60000 6792 0 FreeSans 480 0 0 0 temp1_dac_i[1]
port 162 nsew signal input
flabel metal3 s 59200 7488 60000 7608 0 FreeSans 480 0 0 0 temp1_dac_i[2]
port 163 nsew signal input
flabel metal3 s 59200 8304 60000 8424 0 FreeSans 480 0 0 0 temp1_dac_i[3]
port 164 nsew signal input
flabel metal3 s 59200 9120 60000 9240 0 FreeSans 480 0 0 0 temp1_dac_i[4]
port 165 nsew signal input
flabel metal3 s 59200 9936 60000 10056 0 FreeSans 480 0 0 0 temp1_dac_i[5]
port 166 nsew signal input
flabel metal3 s 59200 30336 60000 30456 0 FreeSans 480 0 0 0 temp1_ticks_i[0]
port 167 nsew signal input
flabel metal3 s 59200 38496 60000 38616 0 FreeSans 480 0 0 0 temp1_ticks_i[10]
port 168 nsew signal input
flabel metal3 s 59200 39312 60000 39432 0 FreeSans 480 0 0 0 temp1_ticks_i[11]
port 169 nsew signal input
flabel metal3 s 59200 31152 60000 31272 0 FreeSans 480 0 0 0 temp1_ticks_i[1]
port 170 nsew signal input
flabel metal3 s 59200 31968 60000 32088 0 FreeSans 480 0 0 0 temp1_ticks_i[2]
port 171 nsew signal input
flabel metal3 s 59200 32784 60000 32904 0 FreeSans 480 0 0 0 temp1_ticks_i[3]
port 172 nsew signal input
flabel metal3 s 59200 33600 60000 33720 0 FreeSans 480 0 0 0 temp1_ticks_i[4]
port 173 nsew signal input
flabel metal3 s 59200 34416 60000 34536 0 FreeSans 480 0 0 0 temp1_ticks_i[5]
port 174 nsew signal input
flabel metal3 s 59200 35232 60000 35352 0 FreeSans 480 0 0 0 temp1_ticks_i[6]
port 175 nsew signal input
flabel metal3 s 59200 36048 60000 36168 0 FreeSans 480 0 0 0 temp1_ticks_i[7]
port 176 nsew signal input
flabel metal3 s 59200 36864 60000 36984 0 FreeSans 480 0 0 0 temp1_ticks_i[8]
port 177 nsew signal input
flabel metal3 s 59200 37680 60000 37800 0 FreeSans 480 0 0 0 temp1_ticks_i[9]
port 178 nsew signal input
flabel metal3 s 59200 10752 60000 10872 0 FreeSans 480 0 0 0 temp2_dac_i[0]
port 179 nsew signal input
flabel metal3 s 59200 11568 60000 11688 0 FreeSans 480 0 0 0 temp2_dac_i[1]
port 180 nsew signal input
flabel metal3 s 59200 12384 60000 12504 0 FreeSans 480 0 0 0 temp2_dac_i[2]
port 181 nsew signal input
flabel metal3 s 59200 13200 60000 13320 0 FreeSans 480 0 0 0 temp2_dac_i[3]
port 182 nsew signal input
flabel metal3 s 59200 14016 60000 14136 0 FreeSans 480 0 0 0 temp2_dac_i[4]
port 183 nsew signal input
flabel metal3 s 59200 14832 60000 14952 0 FreeSans 480 0 0 0 temp2_dac_i[5]
port 184 nsew signal input
flabel metal3 s 59200 40128 60000 40248 0 FreeSans 480 0 0 0 temp2_ticks_i[0]
port 185 nsew signal input
flabel metal3 s 59200 48288 60000 48408 0 FreeSans 480 0 0 0 temp2_ticks_i[10]
port 186 nsew signal input
flabel metal3 s 59200 49104 60000 49224 0 FreeSans 480 0 0 0 temp2_ticks_i[11]
port 187 nsew signal input
flabel metal3 s 59200 40944 60000 41064 0 FreeSans 480 0 0 0 temp2_ticks_i[1]
port 188 nsew signal input
flabel metal3 s 59200 41760 60000 41880 0 FreeSans 480 0 0 0 temp2_ticks_i[2]
port 189 nsew signal input
flabel metal3 s 59200 42576 60000 42696 0 FreeSans 480 0 0 0 temp2_ticks_i[3]
port 190 nsew signal input
flabel metal3 s 59200 43392 60000 43512 0 FreeSans 480 0 0 0 temp2_ticks_i[4]
port 191 nsew signal input
flabel metal3 s 59200 44208 60000 44328 0 FreeSans 480 0 0 0 temp2_ticks_i[5]
port 192 nsew signal input
flabel metal3 s 59200 45024 60000 45144 0 FreeSans 480 0 0 0 temp2_ticks_i[6]
port 193 nsew signal input
flabel metal3 s 59200 45840 60000 45960 0 FreeSans 480 0 0 0 temp2_ticks_i[7]
port 194 nsew signal input
flabel metal3 s 59200 46656 60000 46776 0 FreeSans 480 0 0 0 temp2_ticks_i[8]
port 195 nsew signal input
flabel metal3 s 59200 47472 60000 47592 0 FreeSans 480 0 0 0 temp2_ticks_i[9]
port 196 nsew signal input
flabel metal3 s 59200 15648 60000 15768 0 FreeSans 480 0 0 0 temp3_dac_i[0]
port 197 nsew signal input
flabel metal3 s 59200 16464 60000 16584 0 FreeSans 480 0 0 0 temp3_dac_i[1]
port 198 nsew signal input
flabel metal3 s 59200 17280 60000 17400 0 FreeSans 480 0 0 0 temp3_dac_i[2]
port 199 nsew signal input
flabel metal3 s 59200 18096 60000 18216 0 FreeSans 480 0 0 0 temp3_dac_i[3]
port 200 nsew signal input
flabel metal3 s 59200 18912 60000 19032 0 FreeSans 480 0 0 0 temp3_dac_i[4]
port 201 nsew signal input
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 temp3_dac_i[5]
port 202 nsew signal input
flabel metal3 s 59200 49920 60000 50040 0 FreeSans 480 0 0 0 temp3_ticks_i[0]
port 203 nsew signal input
flabel metal3 s 59200 58080 60000 58200 0 FreeSans 480 0 0 0 temp3_ticks_i[10]
port 204 nsew signal input
flabel metal3 s 59200 58896 60000 59016 0 FreeSans 480 0 0 0 temp3_ticks_i[11]
port 205 nsew signal input
flabel metal3 s 59200 50736 60000 50856 0 FreeSans 480 0 0 0 temp3_ticks_i[1]
port 206 nsew signal input
flabel metal3 s 59200 51552 60000 51672 0 FreeSans 480 0 0 0 temp3_ticks_i[2]
port 207 nsew signal input
flabel metal3 s 59200 52368 60000 52488 0 FreeSans 480 0 0 0 temp3_ticks_i[3]
port 208 nsew signal input
flabel metal3 s 59200 53184 60000 53304 0 FreeSans 480 0 0 0 temp3_ticks_i[4]
port 209 nsew signal input
flabel metal3 s 59200 54000 60000 54120 0 FreeSans 480 0 0 0 temp3_ticks_i[5]
port 210 nsew signal input
flabel metal3 s 59200 54816 60000 54936 0 FreeSans 480 0 0 0 temp3_ticks_i[6]
port 211 nsew signal input
flabel metal3 s 59200 55632 60000 55752 0 FreeSans 480 0 0 0 temp3_ticks_i[7]
port 212 nsew signal input
flabel metal3 s 59200 56448 60000 56568 0 FreeSans 480 0 0 0 temp3_ticks_i[8]
port 213 nsew signal input
flabel metal3 s 59200 57264 60000 57384 0 FreeSans 480 0 0 0 temp3_ticks_i[9]
port 214 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 temp_dac_o[0]
port 215 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 temp_dac_o[1]
port 216 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 temp_dac_o[2]
port 217 nsew signal tristate
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 temp_dac_o[3]
port 218 nsew signal tristate
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 temp_dac_o[4]
port 219 nsew signal tristate
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 temp_dac_o[5]
port 220 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 temp_sel_i[0]
port 221 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 temp_sel_i[1]
port 222 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 temp_ticks_o[0]
port 223 nsew signal tristate
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 temp_ticks_o[10]
port 224 nsew signal tristate
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 temp_ticks_o[11]
port 225 nsew signal tristate
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 temp_ticks_o[1]
port 226 nsew signal tristate
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 temp_ticks_o[2]
port 227 nsew signal tristate
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 temp_ticks_o[3]
port 228 nsew signal tristate
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 temp_ticks_o[4]
port 229 nsew signal tristate
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 temp_ticks_o[5]
port 230 nsew signal tristate
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 temp_ticks_o[6]
port 231 nsew signal tristate
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 temp_ticks_o[7]
port 232 nsew signal tristate
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 temp_ticks_o[8]
port 233 nsew signal tristate
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 temp_ticks_o[9]
port 234 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 235 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 235 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 236 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 236 nsew ground bidirectional
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal1 7912 18190 7912 18190 0 _000_
rlabel metal1 8096 19278 8096 19278 0 _001_
rlabel metal1 8464 12886 8464 12886 0 _002_
rlabel metal2 15318 23426 15318 23426 0 _003_
rlabel metal1 9384 23766 9384 23766 0 _004_
rlabel metal1 11914 23154 11914 23154 0 _005_
rlabel metal1 9614 20366 9614 20366 0 _006_
rlabel metal1 12650 26758 12650 26758 0 _007_
rlabel metal1 12236 14450 12236 14450 0 _008_
rlabel metal2 15962 23936 15962 23936 0 _009_
rlabel metal1 19780 18598 19780 18598 0 _010_
rlabel metal1 18377 18870 18377 18870 0 _011_
rlabel metal1 18860 13158 18860 13158 0 _012_
rlabel metal2 9062 11492 9062 11492 0 _013_
rlabel metal2 16974 6018 16974 6018 0 _014_
rlabel metal2 20746 11016 20746 11016 0 _015_
rlabel metal1 4186 3604 4186 3604 0 _016_
rlabel metal1 5152 2958 5152 2958 0 _017_
rlabel metal1 8234 2958 8234 2958 0 _018_
rlabel metal2 2714 5984 2714 5984 0 _019_
rlabel metal1 4560 6970 4560 6970 0 _020_
rlabel metal2 6670 8126 6670 8126 0 _021_
rlabel metal1 4968 9010 4968 9010 0 _022_
rlabel metal2 8326 8670 8326 8670 0 _023_
rlabel metal2 11638 5916 11638 5916 0 _024_
rlabel metal1 15962 8534 15962 8534 0 _025_
rlabel metal2 18354 3230 18354 3230 0 _026_
rlabel metal1 16376 5270 16376 5270 0 _027_
rlabel metal1 18768 5338 18768 5338 0 _028_
rlabel metal1 19918 2890 19918 2890 0 _029_
rlabel metal1 19918 3434 19918 3434 0 _030_
rlabel metal1 14122 3128 14122 3128 0 _031_
rlabel metal2 3910 13702 3910 13702 0 _032_
rlabel metal1 5480 12410 5480 12410 0 _033_
rlabel metal2 2530 18394 2530 18394 0 _034_
rlabel metal2 4278 15334 4278 15334 0 _035_
rlabel metal2 2530 16796 2530 16796 0 _036_
rlabel metal1 4554 11662 4554 11662 0 _037_
rlabel metal2 4738 19788 4738 19788 0 _038_
rlabel metal1 9476 25670 9476 25670 0 _039_
rlabel metal2 13202 22474 13202 22474 0 _040_
rlabel metal2 15686 21148 15686 21148 0 _041_
rlabel metal2 13478 11866 13478 11866 0 _042_
rlabel metal1 17894 13362 17894 13362 0 _043_
rlabel metal2 21482 18088 21482 18088 0 _044_
rlabel metal1 18768 9962 18768 9962 0 _045_
rlabel metal2 21758 7820 21758 7820 0 _046_
rlabel metal2 19642 9248 19642 9248 0 _047_
rlabel metal2 5566 24582 5566 24582 0 _048_
rlabel metal1 9062 22542 9062 22542 0 _049_
rlabel metal1 4830 20366 4830 20366 0 _050_
rlabel metal1 2530 23188 2530 23188 0 _051_
rlabel metal1 4744 22202 4744 22202 0 _052_
rlabel metal2 15594 24412 15594 24412 0 _053_
rlabel metal1 6992 15062 6992 15062 0 _054_
rlabel metal1 13432 20842 13432 20842 0 _055_
rlabel metal1 12052 15402 12052 15402 0 _056_
rlabel metal1 13708 17714 13708 17714 0 _057_
rlabel metal2 16054 18972 16054 18972 0 _058_
rlabel metal2 19458 15980 19458 15980 0 _059_
rlabel metal2 19458 14144 19458 14144 0 _060_
rlabel metal1 17112 8058 17112 8058 0 _061_
rlabel metal1 18400 6358 18400 6358 0 _062_
rlabel metal2 13478 13090 13478 13090 0 _063_
rlabel metal2 32430 54094 32430 54094 0 _064_
rlabel metal2 31878 53618 31878 53618 0 _065_
rlabel metal2 31970 53312 31970 53312 0 _066_
rlabel metal2 32338 54264 32338 54264 0 _067_
rlabel viali 30408 56338 30408 56338 0 _068_
rlabel metal2 28474 56372 28474 56372 0 _069_
rlabel metal2 28290 54468 28290 54468 0 _070_
rlabel metal2 25898 55930 25898 55930 0 _071_
rlabel via1 32979 56338 32979 56338 0 _072_
rlabel metal1 39422 56372 39422 56372 0 _073_
rlabel metal1 33258 55692 33258 55692 0 _074_
rlabel metal1 41607 55726 41607 55726 0 _075_
rlabel metal2 41906 54978 41906 54978 0 _076_
rlabel metal2 42182 55250 42182 55250 0 _077_
rlabel viali 33441 55726 33441 55726 0 _078_
rlabel via2 35834 56355 35834 56355 0 _079_
rlabel metal1 32315 55590 32315 55590 0 _080_
rlabel metal1 28290 56270 28290 56270 0 _081_
rlabel metal1 26220 55930 26220 55930 0 _082_
rlabel metal1 21942 56338 21942 56338 0 _083_
rlabel metal1 25760 56338 25760 56338 0 _084_
rlabel metal2 43470 56576 43470 56576 0 _085_
rlabel viali 33349 56338 33349 56338 0 _086_
rlabel metal1 30038 56168 30038 56168 0 _087_
rlabel metal1 24242 55930 24242 55930 0 _088_
rlabel metal2 23322 55930 23322 55930 0 _089_
rlabel metal2 23138 55930 23138 55930 0 _090_
rlabel metal1 37904 54570 37904 54570 0 _091_
rlabel metal1 36616 54298 36616 54298 0 _092_
rlabel metal1 35190 54536 35190 54536 0 _093_
rlabel via1 25180 54162 25180 54162 0 _094_
rlabel metal1 23782 54264 23782 54264 0 _095_
rlabel metal2 23598 54332 23598 54332 0 _096_
rlabel metal2 35282 55488 35282 55488 0 _097_
rlabel viali 35465 55726 35465 55726 0 _098_
rlabel metal2 34546 55148 34546 55148 0 _099_
rlabel metal1 27572 54162 27572 54162 0 _100_
rlabel metal2 27094 53754 27094 53754 0 _101_
rlabel metal2 23414 53754 23414 53754 0 _102_
rlabel metal1 37858 55624 37858 55624 0 _103_
rlabel via1 35741 56338 35741 56338 0 _104_
rlabel via2 29854 56389 29854 56389 0 _105_
rlabel metal1 28244 55930 28244 55930 0 _106_
rlabel metal2 29946 55930 29946 55930 0 _107_
rlabel metal1 21873 55658 21873 55658 0 _108_
rlabel metal2 36662 56270 36662 56270 0 _109_
rlabel metal1 38364 55930 38364 55930 0 _110_
rlabel metal2 30222 56457 30222 56457 0 _111_
rlabel viali 30039 56333 30039 56333 0 _112_
rlabel metal1 31188 56338 31188 56338 0 _113_
rlabel metal2 21666 57392 21666 57392 0 _114_
rlabel metal1 57408 6426 57408 6426 0 _115_
rlabel metal2 56994 5882 56994 5882 0 _116_
rlabel metal2 58282 4522 58282 4522 0 _117_
rlabel metal1 56350 3536 56350 3536 0 _118_
rlabel metal1 58374 3026 58374 3026 0 _119_
rlabel metal1 40664 3502 40664 3502 0 _120_
rlabel metal2 55338 11084 55338 11084 0 _121_
rlabel metal1 57224 4046 57224 4046 0 _122_
rlabel metal1 50554 26350 50554 26350 0 _123_
rlabel metal1 58052 23154 58052 23154 0 _124_
rlabel metal2 57546 20679 57546 20679 0 _125_
rlabel metal1 57454 3026 57454 3026 0 _126_
rlabel metal1 48438 3502 48438 3502 0 _127_
rlabel metal1 55522 32402 55522 32402 0 _128_
rlabel metal1 54602 34714 54602 34714 0 _129_
rlabel metal2 52394 34782 52394 34782 0 _130_
rlabel metal1 57684 4114 57684 4114 0 _131_
rlabel metal1 54740 3162 54740 3162 0 _132_
rlabel metal1 55752 4114 55752 4114 0 _133_
rlabel metal1 56810 3502 56810 3502 0 _134_
rlabel metal1 20608 18054 20608 18054 0 _135_
rlabel metal1 19504 24378 19504 24378 0 _136_
rlabel metal1 6164 26962 6164 26962 0 _137_
rlabel metal1 7176 27438 7176 27438 0 _138_
rlabel metal1 8556 26962 8556 26962 0 _139_
rlabel metal2 9154 25466 9154 25466 0 _140_
rlabel metal2 7222 26044 7222 26044 0 _141_
rlabel metal1 10212 28050 10212 28050 0 _142_
rlabel metal2 9890 28220 9890 28220 0 _143_
rlabel metal2 12374 27132 12374 27132 0 _144_
rlabel metal2 13018 26554 13018 26554 0 _145_
rlabel metal1 17112 26214 17112 26214 0 _146_
rlabel metal1 19872 18734 19872 18734 0 _147_
rlabel metal2 20286 18564 20286 18564 0 _148_
rlabel metal1 19964 13294 19964 13294 0 _149_
rlabel metal2 19918 11322 19918 11322 0 _150_
rlabel metal2 22586 6460 22586 6460 0 _151_
rlabel metal2 22586 11322 22586 11322 0 _152_
rlabel metal2 23230 3298 23230 3298 0 _153_
rlabel metal1 23506 3570 23506 3570 0 _154_
rlabel metal1 2438 4012 2438 4012 0 _155_
rlabel metal1 3496 3162 3496 3162 0 _156_
rlabel metal1 3220 4114 3220 4114 0 _157_
rlabel metal1 3220 3026 3220 3026 0 _158_
rlabel metal2 2530 6460 2530 6460 0 _159_
rlabel metal1 3128 7378 3128 7378 0 _160_
rlabel metal2 2990 8636 2990 8636 0 _161_
rlabel metal1 3128 9554 3128 9554 0 _162_
rlabel metal1 8878 8942 8878 8942 0 _163_
rlabel metal2 19458 6460 19458 6460 0 _164_
rlabel metal1 19136 8466 19136 8466 0 _165_
rlabel metal1 19320 3502 19320 3502 0 _166_
rlabel metal2 19826 6086 19826 6086 0 _167_
rlabel metal1 19688 5202 19688 5202 0 _168_
rlabel metal2 20562 3196 20562 3196 0 _169_
rlabel metal2 22126 3706 22126 3706 0 _170_
rlabel metal2 22402 3196 22402 3196 0 _171_
rlabel metal1 21436 16694 21436 16694 0 _172_
rlabel metal1 2162 18224 2162 18224 0 _173_
rlabel metal1 2530 13906 2530 13906 0 _174_
rlabel metal1 2714 12138 2714 12138 0 _175_
rlabel metal2 2714 18564 2714 18564 0 _176_
rlabel metal1 2530 14994 2530 14994 0 _177_
rlabel metal1 2530 17170 2530 17170 0 _178_
rlabel metal1 3266 11662 3266 11662 0 _179_
rlabel metal1 2530 20434 2530 20434 0 _180_
rlabel metal1 9936 25874 9936 25874 0 _181_
rlabel metal1 13616 25874 13616 25874 0 _182_
rlabel metal1 18584 22610 18584 22610 0 _183_
rlabel metal2 19826 12410 19826 12410 0 _184_
rlabel metal1 20010 13906 20010 13906 0 _185_
rlabel metal1 21712 16762 21712 16762 0 _186_
rlabel metal2 19918 10234 19918 10234 0 _187_
rlabel metal2 22586 8636 22586 8636 0 _188_
rlabel metal2 22678 9724 22678 9724 0 _189_
rlabel metal1 22218 17510 22218 17510 0 _190_
rlabel metal2 2162 25262 2162 25262 0 _191_
rlabel metal2 2438 25466 2438 25466 0 _192_
rlabel metal1 5244 26350 5244 26350 0 _193_
rlabel metal2 3726 26044 3726 26044 0 _194_
rlabel metal2 2346 23290 2346 23290 0 _195_
rlabel metal2 2714 22916 2714 22916 0 _196_
rlabel metal1 14582 28050 14582 28050 0 _197_
rlabel metal2 6578 28730 6578 28730 0 _198_
rlabel metal1 11454 26962 11454 26962 0 _199_
rlabel metal2 14766 26758 14766 26758 0 _200_
rlabel metal2 15962 26044 15962 26044 0 _201_
rlabel metal1 19044 20434 19044 20434 0 _202_
rlabel metal1 19550 17510 19550 17510 0 _203_
rlabel metal2 22218 14212 22218 14212 0 _204_
rlabel metal1 19872 7854 19872 7854 0 _205_
rlabel metal2 22126 7242 22126 7242 0 _206_
rlabel metal1 22586 12614 22586 12614 0 _207_
rlabel metal2 13018 14348 13018 14348 0 clknet_0_reg_wr_i
rlabel metal2 9614 3298 9614 3298 0 clknet_3_0__leaf_reg_wr_i
rlabel metal1 6532 13294 6532 13294 0 clknet_3_1__leaf_reg_wr_i
rlabel metal1 18400 3502 18400 3502 0 clknet_3_2__leaf_reg_wr_i
rlabel metal1 17986 13260 17986 13260 0 clknet_3_3__leaf_reg_wr_i
rlabel metal2 9200 16626 9200 16626 0 clknet_3_4__leaf_reg_wr_i
rlabel metal1 7774 19380 7774 19380 0 clknet_3_5__leaf_reg_wr_i
rlabel metal1 14536 17646 14536 17646 0 clknet_3_6__leaf_reg_wr_i
rlabel metal2 12466 22848 12466 22848 0 clknet_3_7__leaf_reg_wr_i
rlabel metal1 56488 2414 56488 2414 0 loopback_i
rlabel metal2 57546 1520 57546 1520 0 loopback_o
rlabel metal1 1932 57426 1932 57426 0 mux0_i[0]
rlabel metal1 3174 57426 3174 57426 0 mux0_i[1]
rlabel metal1 4324 57426 4324 57426 0 mux0_i[2]
rlabel metal1 5796 57426 5796 57426 0 mux0_i[3]
rlabel metal1 6716 57426 6716 57426 0 mux0_i[4]
rlabel metal1 8234 57426 8234 57426 0 mux0_i[5]
rlabel metal1 9108 57426 9108 57426 0 mux1_i[0]
rlabel metal1 10304 57426 10304 57426 0 mux1_i[1]
rlabel metal1 11316 57494 11316 57494 0 mux1_i[2]
rlabel metal1 12696 57426 12696 57426 0 mux1_i[3]
rlabel metal1 13800 57494 13800 57494 0 mux1_i[4]
rlabel metal1 15088 57426 15088 57426 0 mux1_i[5]
rlabel metal1 16721 57426 16721 57426 0 mux2_i[0]
rlabel metal1 17480 57426 17480 57426 0 mux2_i[1]
rlabel metal1 18676 57426 18676 57426 0 mux2_i[2]
rlabel metal1 19964 57426 19964 57426 0 mux2_i[3]
rlabel metal1 21068 57426 21068 57426 0 mux2_i[4]
rlabel metal1 22264 57426 22264 57426 0 mux2_i[5]
rlabel metal1 23460 57426 23460 57426 0 mux3_i[0]
rlabel metal1 24656 57426 24656 57426 0 mux3_i[1]
rlabel metal1 25622 57562 25622 57562 0 mux3_i[2]
rlabel metal1 26818 57562 26818 57562 0 mux3_i[3]
rlabel metal1 28244 57426 28244 57426 0 mux3_i[4]
rlabel metal1 29302 57562 29302 57562 0 mux3_i[5]
rlabel metal1 30636 57426 30636 57426 0 mux4_i[0]
rlabel metal1 32062 57426 32062 57426 0 mux4_i[1]
rlabel metal1 33028 57426 33028 57426 0 mux4_i[2]
rlabel metal1 34224 57562 34224 57562 0 mux4_i[3]
rlabel metal1 35558 57426 35558 57426 0 mux4_i[4]
rlabel metal1 36708 57426 36708 57426 0 mux4_i[5]
rlabel metal1 37904 57426 37904 57426 0 mux5_i[0]
rlabel metal1 39100 57426 39100 57426 0 mux5_i[1]
rlabel metal1 40296 57426 40296 57426 0 mux5_i[2]
rlabel metal2 41354 58320 41354 58320 0 mux5_i[3]
rlabel metal2 42688 57426 42688 57426 0 mux5_i[4]
rlabel metal1 43884 57426 43884 57426 0 mux5_i[5]
rlabel metal1 45172 57426 45172 57426 0 mux6_i[0]
rlabel metal1 46276 57426 46276 57426 0 mux6_i[1]
rlabel metal1 47656 57426 47656 57426 0 mux6_i[2]
rlabel metal1 48668 57426 48668 57426 0 mux6_i[3]
rlabel metal1 50140 57426 50140 57426 0 mux6_i[4]
rlabel metal1 51152 57426 51152 57426 0 mux6_i[5]
rlabel metal1 52256 57426 52256 57426 0 mux7_i[0]
rlabel metal1 53452 57426 53452 57426 0 mux7_i[1]
rlabel metal1 54648 57426 54648 57426 0 mux7_i[2]
rlabel metal1 55844 57426 55844 57426 0 mux7_i[3]
rlabel metal1 57040 57426 57040 57426 0 mux7_i[4]
rlabel metal1 58236 57426 58236 57426 0 mux7_i[5]
rlabel metal1 24564 2346 24564 2346 0 mux_adr_i[0]
rlabel metal1 25622 2346 25622 2346 0 mux_adr_i[1]
rlabel metal2 26634 1520 26634 1520 0 mux_adr_i[2]
rlabel metal1 27876 2822 27876 2822 0 mux_o[0]
rlabel metal2 28842 1520 28842 1520 0 mux_o[1]
rlabel metal2 29946 1520 29946 1520 0 mux_o[2]
rlabel metal2 31050 1520 31050 1520 0 mux_o[3]
rlabel metal2 32154 1520 32154 1520 0 mux_o[4]
rlabel metal2 33258 1520 33258 1520 0 mux_o[5]
rlabel metal1 57086 2618 57086 2618 0 net1
rlabel metal1 21022 54570 21022 54570 0 net10
rlabel metal1 58236 32198 58236 32198 0 net100
rlabel metal1 58098 33286 58098 33286 0 net101
rlabel metal2 56626 33286 56626 33286 0 net102
rlabel metal2 58374 33660 58374 33660 0 net103
rlabel metal1 56258 34612 56258 34612 0 net104
rlabel metal2 58190 35564 58190 35564 0 net105
rlabel metal1 57822 36890 57822 36890 0 net106
rlabel metal1 56672 37910 56672 37910 0 net107
rlabel via1 57615 5746 57615 5746 0 net108
rlabel metal1 56120 6630 56120 6630 0 net109
rlabel metal1 21022 54230 21022 54230 0 net11
rlabel via1 57615 7922 57615 7922 0 net110
rlabel metal1 58052 9962 58052 9962 0 net111
rlabel metal1 56889 11662 56889 11662 0 net112
rlabel via1 57349 13362 57349 13362 0 net113
rlabel metal1 57776 40358 57776 40358 0 net114
rlabel metal1 59018 48518 59018 48518 0 net115
rlabel metal1 58512 49062 58512 49062 0 net116
rlabel metal3 57753 40052 57753 40052 0 net117
rlabel metal1 58834 41990 58834 41990 0 net118
rlabel metal1 57592 42534 57592 42534 0 net119
rlabel metal2 18998 56474 18998 56474 0 net12
rlabel metal1 58972 43622 58972 43622 0 net120
rlabel metal1 58420 44166 58420 44166 0 net121
rlabel metal1 57730 45254 57730 45254 0 net122
rlabel metal1 58466 45798 58466 45798 0 net123
rlabel metal1 58880 47158 58880 47158 0 net124
rlabel metal1 57086 47430 57086 47430 0 net125
rlabel metal1 57592 8262 57592 8262 0 net126
rlabel metal1 56718 6834 56718 6834 0 net127
rlabel metal1 58466 17510 58466 17510 0 net128
rlabel metal1 57822 18054 57822 18054 0 net129
rlabel metal2 20838 57052 20838 57052 0 net13
rlabel metal1 57408 19482 57408 19482 0 net130
rlabel metal1 58144 19686 58144 19686 0 net131
rlabel metal1 58650 50150 58650 50150 0 net132
rlabel metal1 58328 44302 58328 44302 0 net133
rlabel metal1 57822 56678 57822 56678 0 net134
rlabel metal1 58558 50694 58558 50694 0 net135
rlabel metal1 58604 51782 58604 51782 0 net136
rlabel metal1 58742 52598 58742 52598 0 net137
rlabel metal1 58926 53414 58926 53414 0 net138
rlabel metal1 58696 53958 58696 53958 0 net139
rlabel metal2 17066 56950 17066 56950 0 net14
rlabel metal1 58282 55386 58282 55386 0 net140
rlabel metal1 58374 55590 58374 55590 0 net141
rlabel metal1 58144 56678 58144 56678 0 net142
rlabel metal1 56856 56678 56856 56678 0 net143
rlabel metal1 55614 2380 55614 2380 0 net144
rlabel metal2 36386 2210 36386 2210 0 net145
rlabel metal1 58052 2414 58052 2414 0 net146
rlabel metal1 26910 56134 26910 56134 0 net147
rlabel metal1 23736 55862 23736 55862 0 net148
rlabel metal1 27094 4114 27094 4114 0 net149
rlabel metal2 22034 57018 22034 57018 0 net15
rlabel metal1 31050 2414 31050 2414 0 net150
rlabel metal2 32338 2754 32338 2754 0 net151
rlabel metal1 33304 3162 33304 3162 0 net152
rlabel metal2 2530 3876 2530 3876 0 net153
rlabel via1 16698 13413 16698 13413 0 net154
rlabel metal1 1978 13294 1978 13294 0 net155
rlabel metal2 2438 12920 2438 12920 0 net156
rlabel metal1 1886 14960 1886 14960 0 net157
rlabel metal2 16422 3876 16422 3876 0 net158
rlabel metal1 1748 16558 1748 16558 0 net159
rlabel metal2 18906 55658 18906 55658 0 net16
rlabel metal1 2622 4046 2622 4046 0 net160
rlabel metal1 2576 3502 2576 3502 0 net161
rlabel metal2 2346 6222 2346 6222 0 net162
rlabel metal2 4094 7106 4094 7106 0 net163
rlabel metal1 1886 7888 1886 7888 0 net164
rlabel metal2 2438 9316 2438 9316 0 net165
rlabel metal1 9568 9010 9568 9010 0 net166
rlabel metal1 1886 10608 1886 10608 0 net167
rlabel metal1 2530 10438 2530 10438 0 net168
rlabel metal1 2070 17170 2070 17170 0 net169
rlabel metal2 22310 57052 22310 57052 0 net17
rlabel metal1 2300 24582 2300 24582 0 net170
rlabel metal2 19366 14144 19366 14144 0 net171
rlabel metal2 21206 17714 21206 17714 0 net172
rlabel metal1 2162 28050 2162 28050 0 net173
rlabel metal1 2162 29138 2162 29138 0 net174
rlabel metal1 2162 29614 2162 29614 0 net175
rlabel metal1 2070 12206 2070 12206 0 net176
rlabel metal1 2254 18156 2254 18156 0 net177
rlabel metal1 1978 19822 1978 19822 0 net178
rlabel metal1 2208 17714 2208 17714 0 net179
rlabel metal2 28658 56848 28658 56848 0 net18
rlabel metal1 2254 21522 2254 21522 0 net180
rlabel metal2 1886 21420 1886 21420 0 net181
rlabel metal1 1886 23188 1886 23188 0 net182
rlabel metal2 14306 25194 14306 25194 0 net183
rlabel metal2 2438 23936 2438 23936 0 net184
rlabel metal1 2530 25806 2530 25806 0 net185
rlabel metal1 2162 38930 2162 38930 0 net186
rlabel metal1 2944 39270 2944 39270 0 net187
rlabel metal1 3082 40358 3082 40358 0 net188
rlabel metal1 2990 40902 2990 40902 0 net189
rlabel metal2 28934 56712 28934 56712 0 net19
rlabel metal1 2484 41990 2484 41990 0 net190
rlabel metal1 4370 42534 4370 42534 0 net191
rlabel metal1 4278 26486 4278 26486 0 net192
rlabel metal1 3266 32402 3266 32402 0 net193
rlabel via1 2438 23630 2438 23630 0 net194
rlabel metal1 2392 22746 2392 22746 0 net195
rlabel metal1 1886 34544 1886 34544 0 net196
rlabel metal1 2162 35666 2162 35666 0 net197
rlabel metal1 2162 36142 2162 36142 0 net198
rlabel metal1 2484 37094 2484 37094 0 net199
rlabel metal2 2254 57630 2254 57630 0 net2
rlabel metal2 25070 56814 25070 56814 0 net20
rlabel metal1 2530 37638 2530 37638 0 net200
rlabel metal1 3864 43622 3864 43622 0 net201
rlabel metal1 19136 20570 19136 20570 0 net202
rlabel metal1 18078 18394 18078 18394 0 net203
rlabel metal1 2162 53550 2162 53550 0 net204
rlabel metal1 3634 53958 3634 53958 0 net205
rlabel metal1 2990 55250 2990 55250 0 net206
rlabel metal1 2116 55726 2116 55726 0 net207
rlabel metal1 1932 44370 1932 44370 0 net208
rlabel metal1 2162 45458 2162 45458 0 net209
rlabel metal1 24978 55794 24978 55794 0 net21
rlabel metal1 2116 45934 2116 45934 0 net210
rlabel metal1 4554 46954 4554 46954 0 net211
rlabel metal1 2162 47634 2162 47634 0 net212
rlabel metal1 2162 48722 2162 48722 0 net213
rlabel metal2 2438 48960 2438 48960 0 net214
rlabel metal2 2438 50048 2438 50048 0 net215
rlabel metal2 16790 23596 16790 23596 0 net216
rlabel metal2 37766 2754 37766 2754 0 net217
rlabel metal1 38594 2414 38594 2414 0 net218
rlabel metal2 39238 2652 39238 2652 0 net219
rlabel metal1 25116 54706 25116 54706 0 net22
rlabel metal2 40342 2890 40342 2890 0 net220
rlabel metal1 53452 10438 53452 10438 0 net221
rlabel metal2 58190 3128 58190 3128 0 net222
rlabel metal1 44114 3162 44114 3162 0 net223
rlabel metal2 55522 2890 55522 2890 0 net224
rlabel metal1 55798 2448 55798 2448 0 net225
rlabel metal2 44850 4658 44850 4658 0 net226
rlabel metal2 57270 18938 57270 18938 0 net227
rlabel metal1 47886 2448 47886 2448 0 net228
rlabel metal1 48024 3366 48024 3366 0 net229
rlabel metal1 26910 54162 26910 54162 0 net23
rlabel metal1 51980 32334 51980 32334 0 net230
rlabel metal1 52716 2822 52716 2822 0 net231
rlabel metal1 51428 2414 51428 2414 0 net232
rlabel metal2 53406 3196 53406 3196 0 net233
rlabel metal1 54004 2414 54004 2414 0 net234
rlabel metal1 9437 6358 9437 6358 0 net235
rlabel metal2 5198 12823 5198 12823 0 net236
rlabel metal2 16238 11934 16238 11934 0 net237
rlabel metal2 14858 9180 14858 9180 0 net238
rlabel metal1 9423 20502 9423 20502 0 net239
rlabel metal2 28566 56508 28566 56508 0 net24
rlabel metal2 5290 19550 5290 19550 0 net240
rlabel metal2 16698 14858 16698 14858 0 net241
rlabel metal2 16054 21386 16054 21386 0 net242
rlabel metal1 14352 3502 14352 3502 0 net243
rlabel metal2 29762 57052 29762 57052 0 net25
rlabel metal2 33166 56508 33166 56508 0 net26
rlabel metal1 32798 56406 32798 56406 0 net27
rlabel metal1 35466 54706 35466 54706 0 net28
rlabel metal1 35006 55658 35006 55658 0 net29
rlabel metal2 3450 56474 3450 56474 0 net3
rlabel metal2 35466 56814 35466 56814 0 net30
rlabel metal2 36570 56814 36570 56814 0 net31
rlabel metal1 36478 55760 36478 55760 0 net32
rlabel metal1 38502 56372 38502 56372 0 net33
rlabel metal2 37674 55726 37674 55726 0 net34
rlabel metal1 38962 56848 38962 56848 0 net35
rlabel metal2 40526 56814 40526 56814 0 net36
rlabel metal2 40066 56576 40066 56576 0 net37
rlabel viali 41813 56338 41813 56338 0 net38
rlabel viali 44021 56814 44021 56814 0 net39
rlabel metal1 17618 57528 17618 57528 0 net4
rlabel viali 43837 55726 43837 55726 0 net40
rlabel viali 43929 55250 43929 55250 0 net41
rlabel viali 42089 55726 42089 55726 0 net42
rlabel viali 43837 56338 43837 56338 0 net43
rlabel metal2 52210 56814 52210 56814 0 net44
rlabel metal2 53406 56950 53406 56950 0 net45
rlabel metal2 54602 56406 54602 56406 0 net46
rlabel metal2 54694 56270 54694 56270 0 net47
rlabel metal1 56097 57290 56097 57290 0 net48
rlabel metal2 58190 56746 58190 56746 0 net49
rlabel metal2 5750 55386 5750 55386 0 net5
rlabel metal1 26818 2618 26818 2618 0 net50
rlabel metal1 26151 2414 26151 2414 0 net51
rlabel metal1 32246 55250 32246 55250 0 net52
rlabel metal2 4830 2176 4830 2176 0 net53
rlabel metal2 5934 2074 5934 2074 0 net54
rlabel metal1 2208 3026 2208 3026 0 net55
rlabel metal1 18676 2482 18676 2482 0 net56
rlabel metal1 20102 17578 20102 17578 0 net57
rlabel metal1 20332 2482 20332 2482 0 net58
rlabel metal1 20378 3366 20378 3366 0 net59
rlabel metal2 6946 56576 6946 56576 0 net6
rlabel metal1 22724 4182 22724 4182 0 net60
rlabel metal1 23092 2618 23092 2618 0 net61
rlabel metal1 2530 4250 2530 4250 0 net62
rlabel metal1 2438 3366 2438 3366 0 net63
rlabel metal2 10258 2108 10258 2108 0 net64
rlabel metal1 4278 2278 4278 2278 0 net65
rlabel metal1 8326 2550 8326 2550 0 net66
rlabel metal2 13570 2142 13570 2142 0 net67
rlabel metal1 12558 2482 12558 2482 0 net68
rlabel metal1 15548 25126 15548 25126 0 net69
rlabel metal2 8326 56338 8326 56338 0 net7
rlabel metal1 17986 2550 17986 2550 0 net70
rlabel metal1 3680 2618 3680 2618 0 net71
rlabel metal2 56718 4420 56718 4420 0 net72
rlabel metal1 56718 2822 56718 2822 0 net73
rlabel metal1 57132 2278 57132 2278 0 net74
rlabel metal2 57454 8364 57454 8364 0 net75
rlabel metal2 58282 9316 58282 9316 0 net76
rlabel metal1 58374 5338 58374 5338 0 net77
rlabel metal1 58236 21114 58236 21114 0 net78
rlabel metal2 57638 37332 57638 37332 0 net79
rlabel metal2 17894 56678 17894 56678 0 net8
rlabel metal2 59110 35020 59110 35020 0 net80
rlabel metal2 58190 23460 58190 23460 0 net81
rlabel metal1 58466 21862 58466 21862 0 net82
rlabel metal1 57500 22746 57500 22746 0 net83
rlabel metal1 56626 32538 56626 32538 0 net84
rlabel metal1 58420 32878 58420 32878 0 net85
rlabel metal1 56718 26010 56718 26010 0 net86
rlabel metal1 58420 35054 58420 35054 0 net87
rlabel metal1 57592 37094 57592 37094 0 net88
rlabel metal1 57868 37638 57868 37638 0 net89
rlabel metal1 19366 56984 19366 56984 0 net9
rlabel metal1 56810 5746 56810 5746 0 net90
rlabel metal1 57868 6630 57868 6630 0 net91
rlabel metal1 57408 7514 57408 7514 0 net92
rlabel metal1 58098 8330 58098 8330 0 net93
rlabel metal1 58144 9146 58144 9146 0 net94
rlabel metal1 58328 9418 58328 9418 0 net95
rlabel metal1 58420 26418 58420 26418 0 net96
rlabel metal1 57178 39066 57178 39066 0 net97
rlabel metal1 57546 38318 57546 38318 0 net98
rlabel metal1 58328 25330 58328 25330 0 net99
rlabel metal3 1188 4284 1188 4284 0 reg0_o[0]
rlabel metal3 1188 12444 1188 12444 0 reg0_o[10]
rlabel metal3 1188 13260 1188 13260 0 reg0_o[11]
rlabel via2 1702 14059 1702 14059 0 reg0_o[12]
rlabel metal3 1188 14892 1188 14892 0 reg0_o[13]
rlabel metal3 1188 15708 1188 15708 0 reg0_o[14]
rlabel metal2 1702 16473 1702 16473 0 reg0_o[15]
rlabel metal3 1188 5100 1188 5100 0 reg0_o[1]
rlabel via2 1702 5899 1702 5899 0 reg0_o[2]
rlabel metal2 1702 6579 1702 6579 0 reg0_o[3]
rlabel metal3 1556 7548 1556 7548 0 reg0_o[4]
rlabel metal2 1702 8211 1702 8211 0 reg0_o[5]
rlabel metal2 1702 8891 1702 8891 0 reg0_o[6]
rlabel metal3 1188 9996 1188 9996 0 reg0_o[7]
rlabel via2 1702 10795 1702 10795 0 reg0_o[8]
rlabel metal2 1702 11475 1702 11475 0 reg0_o[9]
rlabel via2 1702 17323 1702 17323 0 reg1_o[0]
rlabel via2 1702 25483 1702 25483 0 reg1_o[10]
rlabel metal3 1188 26316 1188 26316 0 reg1_o[11]
rlabel metal3 1188 27132 1188 27132 0 reg1_o[12]
rlabel metal3 1188 27948 1188 27948 0 reg1_o[13]
rlabel metal3 1188 28764 1188 28764 0 reg1_o[14]
rlabel metal3 1188 29580 1188 29580 0 reg1_o[15]
rlabel metal3 1188 18156 1188 18156 0 reg1_o[1]
rlabel metal3 1188 18972 1188 18972 0 reg1_o[2]
rlabel metal3 1188 19788 1188 19788 0 reg1_o[3]
rlabel via2 1702 20587 1702 20587 0 reg1_o[4]
rlabel metal3 1188 21420 1188 21420 0 reg1_o[5]
rlabel via2 1702 22219 1702 22219 0 reg1_o[6]
rlabel metal3 1188 23052 1188 23052 0 reg1_o[7]
rlabel metal3 1188 23868 1188 23868 0 reg1_o[8]
rlabel metal3 1188 24684 1188 24684 0 reg1_o[9]
rlabel metal3 1188 30396 1188 30396 0 reg2_o[0]
rlabel metal3 1188 38556 1188 38556 0 reg2_o[10]
rlabel metal3 1188 39372 1188 39372 0 reg2_o[11]
rlabel metal3 1188 40188 1188 40188 0 reg2_o[12]
rlabel metal3 1188 41004 1188 41004 0 reg2_o[13]
rlabel metal3 1188 41820 1188 41820 0 reg2_o[14]
rlabel metal3 1188 42636 1188 42636 0 reg2_o[15]
rlabel metal3 1188 31212 1188 31212 0 reg2_o[1]
rlabel metal3 1188 32028 1188 32028 0 reg2_o[2]
rlabel metal3 1188 32844 1188 32844 0 reg2_o[3]
rlabel metal3 1188 33660 1188 33660 0 reg2_o[4]
rlabel metal3 1188 34476 1188 34476 0 reg2_o[5]
rlabel metal3 1188 35292 1188 35292 0 reg2_o[6]
rlabel metal3 1188 36108 1188 36108 0 reg2_o[7]
rlabel metal3 1188 36924 1188 36924 0 reg2_o[8]
rlabel metal3 1188 37740 1188 37740 0 reg2_o[9]
rlabel metal3 1188 43452 1188 43452 0 reg3_o[0]
rlabel metal3 1188 51612 1188 51612 0 reg3_o[10]
rlabel metal3 1188 52428 1188 52428 0 reg3_o[11]
rlabel metal3 1188 53244 1188 53244 0 reg3_o[12]
rlabel metal3 1188 54060 1188 54060 0 reg3_o[13]
rlabel metal3 1188 54876 1188 54876 0 reg3_o[14]
rlabel metal3 1188 55692 1188 55692 0 reg3_o[15]
rlabel metal3 1188 44268 1188 44268 0 reg3_o[1]
rlabel metal3 1188 45084 1188 45084 0 reg3_o[2]
rlabel metal3 1188 45900 1188 45900 0 reg3_o[3]
rlabel metal3 1188 46716 1188 46716 0 reg3_o[4]
rlabel metal3 1188 47532 1188 47532 0 reg3_o[5]
rlabel metal3 1188 48348 1188 48348 0 reg3_o[6]
rlabel metal3 1188 49164 1188 49164 0 reg3_o[7]
rlabel metal3 1188 49980 1188 49980 0 reg3_o[8]
rlabel metal3 1188 50796 1188 50796 0 reg3_o[9]
rlabel metal1 4600 2414 4600 2414 0 reg_adr_i[0]
rlabel metal1 5704 2414 5704 2414 0 reg_adr_i[1]
rlabel metal2 6762 1571 6762 1571 0 reg_dat_i[0]
rlabel metal1 17848 2414 17848 2414 0 reg_dat_i[10]
rlabel metal1 17710 2958 17710 2958 0 reg_dat_i[11]
rlabel metal2 20010 1435 20010 1435 0 reg_dat_i[12]
rlabel metal2 21390 3740 21390 3740 0 reg_dat_i[13]
rlabel metal1 22310 2380 22310 2380 0 reg_dat_i[14]
rlabel metal1 23552 2414 23552 2414 0 reg_dat_i[15]
rlabel metal1 8004 2346 8004 2346 0 reg_dat_i[1]
rlabel metal1 8924 2414 8924 2414 0 reg_dat_i[2]
rlabel metal1 10212 2346 10212 2346 0 reg_dat_i[3]
rlabel metal1 11132 2346 11132 2346 0 reg_dat_i[4]
rlabel metal1 12328 2414 12328 2414 0 reg_dat_i[5]
rlabel metal1 12788 2346 12788 2346 0 reg_dat_i[6]
rlabel metal1 14628 2346 14628 2346 0 reg_dat_i[7]
rlabel metal1 15686 2346 15686 2346 0 reg_dat_i[8]
rlabel metal1 16836 2346 16836 2346 0 reg_dat_i[9]
rlabel metal1 11454 12818 11454 12818 0 reg_wr_i
rlabel metal2 2438 3162 2438 3162 0 rst_n_i
rlabel metal1 56718 3026 56718 3026 0 temp0_dac_i[0]
rlabel metal2 56074 2431 56074 2431 0 temp0_dac_i[1]
rlabel metal2 57546 2533 57546 2533 0 temp0_dac_i[2]
rlabel metal2 57730 4029 57730 4029 0 temp0_dac_i[3]
rlabel metal2 58374 4437 58374 4437 0 temp0_dac_i[4]
rlabel metal2 58374 5151 58374 5151 0 temp0_dac_i[5]
rlabel metal2 58374 20757 58374 20757 0 temp0_ticks_i[0]
rlabel metal2 58374 28645 58374 28645 0 temp0_ticks_i[10]
rlabel metal1 58144 29138 58144 29138 0 temp0_ticks_i[11]
rlabel metal2 58374 21471 58374 21471 0 temp0_ticks_i[1]
rlabel metal1 58052 21998 58052 21998 0 temp0_ticks_i[2]
rlabel metal2 58374 22831 58374 22831 0 temp0_ticks_i[3]
rlabel metal2 58374 24021 58374 24021 0 temp0_ticks_i[4]
rlabel metal2 58374 24735 58374 24735 0 temp0_ticks_i[5]
rlabel metal2 57546 25687 57546 25687 0 temp0_ticks_i[6]
rlabel metal2 58374 26095 58374 26095 0 temp0_ticks_i[7]
rlabel via2 58374 27115 58374 27115 0 temp0_ticks_i[8]
rlabel metal2 58374 27999 58374 27999 0 temp0_ticks_i[9]
rlabel metal2 58374 6103 58374 6103 0 temp1_dac_i[0]
rlabel via2 58374 6749 58374 6749 0 temp1_dac_i[1]
rlabel metal2 58374 7463 58374 7463 0 temp1_dac_i[2]
rlabel metal2 58374 8415 58374 8415 0 temp1_dac_i[3]
rlabel metal2 58374 9061 58374 9061 0 temp1_dac_i[4]
rlabel metal1 58006 9554 58006 9554 0 temp1_dac_i[5]
rlabel metal2 58190 30311 58190 30311 0 temp1_ticks_i[0]
rlabel metal2 58374 38743 58374 38743 0 temp1_ticks_i[10]
rlabel via2 58374 39389 58374 39389 0 temp1_ticks_i[11]
rlabel metal2 58190 31263 58190 31263 0 temp1_ticks_i[1]
rlabel via2 58374 32011 58374 32011 0 temp1_ticks_i[2]
rlabel metal1 58144 33490 58144 33490 0 temp1_ticks_i[3]
rlabel metal1 58420 33966 58420 33966 0 temp1_ticks_i[4]
rlabel metal1 58052 34578 58052 34578 0 temp1_ticks_i[5]
rlabel metal2 58374 35479 58374 35479 0 temp1_ticks_i[6]
rlabel via2 58374 36125 58374 36125 0 temp1_ticks_i[7]
rlabel metal2 58374 36839 58374 36839 0 temp1_ticks_i[8]
rlabel metal2 58374 37791 58374 37791 0 temp1_ticks_i[9]
rlabel metal1 58420 11118 58420 11118 0 temp2_dac_i[0]
rlabel metal2 58374 11679 58374 11679 0 temp2_dac_i[1]
rlabel metal2 58374 12325 58374 12325 0 temp2_dac_i[2]
rlabel metal2 58374 13039 58374 13039 0 temp2_dac_i[3]
rlabel metal2 58374 14229 58374 14229 0 temp2_dac_i[4]
rlabel metal2 58374 14943 58374 14943 0 temp2_dac_i[5]
rlabel metal2 58374 40341 58374 40341 0 temp2_ticks_i[0]
rlabel metal2 58374 48535 58374 48535 0 temp2_ticks_i[10]
rlabel via2 58374 49181 58374 49181 0 temp2_ticks_i[11]
rlabel metal3 58842 41004 58842 41004 0 temp2_ticks_i[1]
rlabel metal2 58374 42007 58374 42007 0 temp2_ticks_i[2]
rlabel via2 58374 42653 58374 42653 0 temp2_ticks_i[3]
rlabel metal2 58374 43605 58374 43605 0 temp2_ticks_i[4]
rlabel metal2 58374 44319 58374 44319 0 temp2_ticks_i[5]
rlabel metal2 58374 45271 58374 45271 0 temp2_ticks_i[6]
rlabel via2 58374 45917 58374 45917 0 temp2_ticks_i[7]
rlabel metal2 58374 46869 58374 46869 0 temp2_ticks_i[8]
rlabel metal2 58374 47583 58374 47583 0 temp2_ticks_i[9]
rlabel via2 58374 15691 58374 15691 0 temp3_dac_i[0]
rlabel via2 58374 16541 58374 16541 0 temp3_dac_i[1]
rlabel metal2 58374 17493 58374 17493 0 temp3_dac_i[2]
rlabel metal2 58374 18207 58374 18207 0 temp3_dac_i[3]
rlabel via2 58374 18955 58374 18955 0 temp3_dac_i[4]
rlabel via2 58374 19805 58374 19805 0 temp3_dac_i[5]
rlabel metal2 58374 50133 58374 50133 0 temp3_ticks_i[0]
rlabel metal1 58420 56338 58420 56338 0 temp3_ticks_i[10]
rlabel metal2 57546 57885 57546 57885 0 temp3_ticks_i[11]
rlabel metal2 58374 50847 58374 50847 0 temp3_ticks_i[1]
rlabel metal2 58374 51799 58374 51799 0 temp3_ticks_i[2]
rlabel via2 58374 52445 58374 52445 0 temp3_ticks_i[3]
rlabel metal2 58374 53397 58374 53397 0 temp3_ticks_i[4]
rlabel metal2 58374 54111 58374 54111 0 temp3_ticks_i[5]
rlabel metal1 57960 55250 57960 55250 0 temp3_ticks_i[6]
rlabel via2 58374 55709 58374 55709 0 temp3_ticks_i[7]
rlabel metal2 58374 56661 58374 56661 0 temp3_ticks_i[8]
rlabel metal2 57086 57069 57086 57069 0 temp3_ticks_i[9]
rlabel metal2 36570 1520 36570 1520 0 temp_dac_o[0]
rlabel metal2 37674 1520 37674 1520 0 temp_dac_o[1]
rlabel metal2 38778 1520 38778 1520 0 temp_dac_o[2]
rlabel metal2 39882 1520 39882 1520 0 temp_dac_o[3]
rlabel metal2 40986 1520 40986 1520 0 temp_dac_o[4]
rlabel metal2 42090 1520 42090 1520 0 temp_dac_o[5]
rlabel metal2 34362 1520 34362 1520 0 temp_sel_i[0]
rlabel metal1 36064 2414 36064 2414 0 temp_sel_i[1]
rlabel metal2 43194 1520 43194 1520 0 temp_ticks_o[0]
rlabel metal2 54234 1520 54234 1520 0 temp_ticks_o[10]
rlabel metal2 55338 1520 55338 1520 0 temp_ticks_o[11]
rlabel metal2 44298 1520 44298 1520 0 temp_ticks_o[1]
rlabel metal2 45402 1520 45402 1520 0 temp_ticks_o[2]
rlabel metal2 46506 1520 46506 1520 0 temp_ticks_o[3]
rlabel metal2 47610 1520 47610 1520 0 temp_ticks_o[4]
rlabel metal2 48714 1520 48714 1520 0 temp_ticks_o[5]
rlabel metal2 49818 1520 49818 1520 0 temp_ticks_o[6]
rlabel metal2 50922 1520 50922 1520 0 temp_ticks_o[7]
rlabel metal2 52026 1520 52026 1520 0 temp_ticks_o[8]
rlabel metal2 53130 1520 53130 1520 0 temp_ticks_o[9]
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
