magic
tech sky130A
magscale 1 2
timestamp 1670943006
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 1104 2128 28888 27792
<< metal2 >>
rect 3790 0 3846 800
rect 11242 0 11298 800
rect 18694 0 18750 800
rect 26146 0 26202 800
<< obsm2 >>
rect 1490 856 28500 28393
rect 1490 800 3734 856
rect 3902 800 11186 856
rect 11354 800 18638 856
rect 18806 800 26090 856
rect 26258 800 28500 856
<< metal3 >>
rect 29200 28296 30000 28416
rect 0 27072 800 27192
rect 29200 25848 30000 25968
rect 29200 23400 30000 23520
rect 0 22176 800 22296
rect 29200 20952 30000 21072
rect 29200 18504 30000 18624
rect 0 17280 800 17400
rect 29200 16056 30000 16176
rect 29200 13608 30000 13728
rect 0 12384 800 12504
rect 29200 11160 30000 11280
rect 29200 8712 30000 8832
rect 0 7488 800 7608
rect 29200 6264 30000 6384
rect 29200 3816 30000 3936
rect 0 2592 800 2712
rect 29200 1368 30000 1488
<< obsm3 >>
rect 800 28216 29120 28389
rect 800 27272 29200 28216
rect 880 26992 29200 27272
rect 800 26048 29200 26992
rect 800 25768 29120 26048
rect 800 23600 29200 25768
rect 800 23320 29120 23600
rect 800 22376 29200 23320
rect 880 22096 29200 22376
rect 800 21152 29200 22096
rect 800 20872 29120 21152
rect 800 18704 29200 20872
rect 800 18424 29120 18704
rect 800 17480 29200 18424
rect 880 17200 29200 17480
rect 800 16256 29200 17200
rect 800 15976 29120 16256
rect 800 13808 29200 15976
rect 800 13528 29120 13808
rect 800 12584 29200 13528
rect 880 12304 29200 12584
rect 800 11360 29200 12304
rect 800 11080 29120 11360
rect 800 8912 29200 11080
rect 800 8632 29120 8912
rect 800 7688 29200 8632
rect 880 7408 29200 7688
rect 800 6464 29200 7408
rect 800 6184 29120 6464
rect 800 4016 29200 6184
rect 800 3736 29120 4016
rect 800 2792 29200 3736
rect 880 2512 29200 2792
rect 800 1568 29200 2512
rect 800 1395 29120 1568
<< metal4 >>
rect 3344 2128 3664 27792
rect 5744 2128 6064 27792
rect 8144 2128 8464 27792
rect 10544 2128 10864 27792
rect 12944 2128 13264 27792
rect 15344 2128 15664 27792
rect 17744 2128 18064 27792
rect 20144 2128 20464 27792
rect 22544 2128 22864 27792
rect 24944 2128 25264 27792
rect 27344 2128 27664 27792
<< labels >>
rlabel metal2 s 3790 0 3846 800 6 clk
port 1 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 conversion_finished_out
port 2 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 rst_n
port 3 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 start_conv_in
port 4 nsew signal input
rlabel metal3 s 29200 1368 30000 1488 6 tick_result_out[0]
port 5 nsew signal output
rlabel metal3 s 29200 25848 30000 25968 6 tick_result_out[10]
port 6 nsew signal output
rlabel metal3 s 29200 28296 30000 28416 6 tick_result_out[11]
port 7 nsew signal output
rlabel metal3 s 29200 3816 30000 3936 6 tick_result_out[1]
port 8 nsew signal output
rlabel metal3 s 29200 6264 30000 6384 6 tick_result_out[2]
port 9 nsew signal output
rlabel metal3 s 29200 8712 30000 8832 6 tick_result_out[3]
port 10 nsew signal output
rlabel metal3 s 29200 11160 30000 11280 6 tick_result_out[4]
port 11 nsew signal output
rlabel metal3 s 29200 13608 30000 13728 6 tick_result_out[5]
port 12 nsew signal output
rlabel metal3 s 29200 16056 30000 16176 6 tick_result_out[6]
port 13 nsew signal output
rlabel metal3 s 29200 18504 30000 18624 6 tick_result_out[7]
port 14 nsew signal output
rlabel metal3 s 29200 20952 30000 21072 6 tick_result_out[8]
port 15 nsew signal output
rlabel metal3 s 29200 23400 30000 23520 6 tick_result_out[9]
port 16 nsew signal output
rlabel metal4 s 3344 2128 3664 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 8144 2128 8464 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 17744 2128 18064 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 22544 2128 22864 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 27344 2128 27664 27792 6 vccd1
port 17 nsew power bidirectional
rlabel metal3 s 0 2592 800 2712 6 vdac_result_out[0]
port 18 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 vdac_result_out[1]
port 19 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 vdac_result_out[2]
port 20 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 vdac_result_out[3]
port 21 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 vdac_result_out[4]
port 22 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 vdac_result_out[5]
port 23 nsew signal output
rlabel metal4 s 5744 2128 6064 27792 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 10544 2128 10864 27792 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 15344 2128 15664 27792 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 20144 2128 20464 27792 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 24944 2128 25264 27792 6 vssd1
port 24 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1482648
string GDS_FILE /foss/designs/openlane/tempsense/runs/foo/results/signoff/tempsense.magic.gds
string GDS_START 366644
<< end >>

