magic
tech sky130A
magscale 1 2
timestamp 1670618896
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 1104 1708 59694 57712
<< metal2 >>
rect 1858 59200 1914 60000
rect 3054 59200 3110 60000
rect 4250 59200 4306 60000
rect 5446 59200 5502 60000
rect 6642 59200 6698 60000
rect 7838 59200 7894 60000
rect 9034 59200 9090 60000
rect 10230 59200 10286 60000
rect 11426 59200 11482 60000
rect 12622 59200 12678 60000
rect 13818 59200 13874 60000
rect 15014 59200 15070 60000
rect 16210 59200 16266 60000
rect 17406 59200 17462 60000
rect 18602 59200 18658 60000
rect 19798 59200 19854 60000
rect 20994 59200 21050 60000
rect 22190 59200 22246 60000
rect 23386 59200 23442 60000
rect 24582 59200 24638 60000
rect 25778 59200 25834 60000
rect 26974 59200 27030 60000
rect 28170 59200 28226 60000
rect 29366 59200 29422 60000
rect 30562 59200 30618 60000
rect 31758 59200 31814 60000
rect 32954 59200 33010 60000
rect 34150 59200 34206 60000
rect 35346 59200 35402 60000
rect 36542 59200 36598 60000
rect 37738 59200 37794 60000
rect 38934 59200 38990 60000
rect 40130 59200 40186 60000
rect 41326 59200 41382 60000
rect 42522 59200 42578 60000
rect 43718 59200 43774 60000
rect 44914 59200 44970 60000
rect 46110 59200 46166 60000
rect 47306 59200 47362 60000
rect 48502 59200 48558 60000
rect 49698 59200 49754 60000
rect 50894 59200 50950 60000
rect 52090 59200 52146 60000
rect 53286 59200 53342 60000
rect 54482 59200 54538 60000
rect 55678 59200 55734 60000
rect 56874 59200 56930 60000
rect 58070 59200 58126 60000
rect 2318 0 2374 800
rect 3422 0 3478 800
rect 4526 0 4582 800
rect 5630 0 5686 800
rect 6734 0 6790 800
rect 7838 0 7894 800
rect 8942 0 8998 800
rect 10046 0 10102 800
rect 11150 0 11206 800
rect 12254 0 12310 800
rect 13358 0 13414 800
rect 14462 0 14518 800
rect 15566 0 15622 800
rect 16670 0 16726 800
rect 17774 0 17830 800
rect 18878 0 18934 800
rect 19982 0 20038 800
rect 21086 0 21142 800
rect 22190 0 22246 800
rect 23294 0 23350 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26606 0 26662 800
rect 27710 0 27766 800
rect 28814 0 28870 800
rect 29918 0 29974 800
rect 31022 0 31078 800
rect 32126 0 32182 800
rect 33230 0 33286 800
rect 34334 0 34390 800
rect 35438 0 35494 800
rect 36542 0 36598 800
rect 37646 0 37702 800
rect 38750 0 38806 800
rect 39854 0 39910 800
rect 40958 0 41014 800
rect 42062 0 42118 800
rect 43166 0 43222 800
rect 44270 0 44326 800
rect 45374 0 45430 800
rect 46478 0 46534 800
rect 47582 0 47638 800
rect 48686 0 48742 800
rect 49790 0 49846 800
rect 50894 0 50950 800
rect 51998 0 52054 800
rect 53102 0 53158 800
rect 54206 0 54262 800
rect 55310 0 55366 800
rect 56414 0 56470 800
rect 57518 0 57574 800
<< obsm2 >>
rect 1674 59144 1802 59200
rect 1970 59144 2998 59200
rect 3166 59144 4194 59200
rect 4362 59144 5390 59200
rect 5558 59144 6586 59200
rect 6754 59144 7782 59200
rect 7950 59144 8978 59200
rect 9146 59144 10174 59200
rect 10342 59144 11370 59200
rect 11538 59144 12566 59200
rect 12734 59144 13762 59200
rect 13930 59144 14958 59200
rect 15126 59144 16154 59200
rect 16322 59144 17350 59200
rect 17518 59144 18546 59200
rect 18714 59144 19742 59200
rect 19910 59144 20938 59200
rect 21106 59144 22134 59200
rect 22302 59144 23330 59200
rect 23498 59144 24526 59200
rect 24694 59144 25722 59200
rect 25890 59144 26918 59200
rect 27086 59144 28114 59200
rect 28282 59144 29310 59200
rect 29478 59144 30506 59200
rect 30674 59144 31702 59200
rect 31870 59144 32898 59200
rect 33066 59144 34094 59200
rect 34262 59144 35290 59200
rect 35458 59144 36486 59200
rect 36654 59144 37682 59200
rect 37850 59144 38878 59200
rect 39046 59144 40074 59200
rect 40242 59144 41270 59200
rect 41438 59144 42466 59200
rect 42634 59144 43662 59200
rect 43830 59144 44858 59200
rect 45026 59144 46054 59200
rect 46222 59144 47250 59200
rect 47418 59144 48446 59200
rect 48614 59144 49642 59200
rect 49810 59144 50838 59200
rect 51006 59144 52034 59200
rect 52202 59144 53230 59200
rect 53398 59144 54426 59200
rect 54594 59144 55622 59200
rect 55790 59144 56818 59200
rect 56986 59144 58014 59200
rect 58182 59144 59688 59200
rect 1674 856 59688 59144
rect 1674 734 2262 856
rect 2430 734 3366 856
rect 3534 734 4470 856
rect 4638 734 5574 856
rect 5742 734 6678 856
rect 6846 734 7782 856
rect 7950 734 8886 856
rect 9054 734 9990 856
rect 10158 734 11094 856
rect 11262 734 12198 856
rect 12366 734 13302 856
rect 13470 734 14406 856
rect 14574 734 15510 856
rect 15678 734 16614 856
rect 16782 734 17718 856
rect 17886 734 18822 856
rect 18990 734 19926 856
rect 20094 734 21030 856
rect 21198 734 22134 856
rect 22302 734 23238 856
rect 23406 734 24342 856
rect 24510 734 25446 856
rect 25614 734 26550 856
rect 26718 734 27654 856
rect 27822 734 28758 856
rect 28926 734 29862 856
rect 30030 734 30966 856
rect 31134 734 32070 856
rect 32238 734 33174 856
rect 33342 734 34278 856
rect 34446 734 35382 856
rect 35550 734 36486 856
rect 36654 734 37590 856
rect 37758 734 38694 856
rect 38862 734 39798 856
rect 39966 734 40902 856
rect 41070 734 42006 856
rect 42174 734 43110 856
rect 43278 734 44214 856
rect 44382 734 45318 856
rect 45486 734 46422 856
rect 46590 734 47526 856
rect 47694 734 48630 856
rect 48798 734 49734 856
rect 49902 734 50838 856
rect 51006 734 51942 856
rect 52110 734 53046 856
rect 53214 734 54150 856
rect 54318 734 55254 856
rect 55422 734 56358 856
rect 56526 734 57462 856
rect 57630 734 59688 856
<< metal3 >>
rect 59200 58896 60000 59016
rect 59200 58080 60000 58200
rect 59200 57264 60000 57384
rect 59200 56448 60000 56568
rect 0 55632 800 55752
rect 59200 55632 60000 55752
rect 0 54816 800 54936
rect 59200 54816 60000 54936
rect 0 54000 800 54120
rect 59200 54000 60000 54120
rect 0 53184 800 53304
rect 59200 53184 60000 53304
rect 0 52368 800 52488
rect 59200 52368 60000 52488
rect 0 51552 800 51672
rect 59200 51552 60000 51672
rect 0 50736 800 50856
rect 59200 50736 60000 50856
rect 0 49920 800 50040
rect 59200 49920 60000 50040
rect 0 49104 800 49224
rect 59200 49104 60000 49224
rect 0 48288 800 48408
rect 59200 48288 60000 48408
rect 0 47472 800 47592
rect 59200 47472 60000 47592
rect 0 46656 800 46776
rect 59200 46656 60000 46776
rect 0 45840 800 45960
rect 59200 45840 60000 45960
rect 0 45024 800 45144
rect 59200 45024 60000 45144
rect 0 44208 800 44328
rect 59200 44208 60000 44328
rect 0 43392 800 43512
rect 59200 43392 60000 43512
rect 0 42576 800 42696
rect 59200 42576 60000 42696
rect 0 41760 800 41880
rect 59200 41760 60000 41880
rect 0 40944 800 41064
rect 59200 40944 60000 41064
rect 0 40128 800 40248
rect 59200 40128 60000 40248
rect 0 39312 800 39432
rect 59200 39312 60000 39432
rect 0 38496 800 38616
rect 59200 38496 60000 38616
rect 0 37680 800 37800
rect 59200 37680 60000 37800
rect 0 36864 800 36984
rect 59200 36864 60000 36984
rect 0 36048 800 36168
rect 59200 36048 60000 36168
rect 0 35232 800 35352
rect 59200 35232 60000 35352
rect 0 34416 800 34536
rect 59200 34416 60000 34536
rect 0 33600 800 33720
rect 59200 33600 60000 33720
rect 0 32784 800 32904
rect 59200 32784 60000 32904
rect 0 31968 800 32088
rect 59200 31968 60000 32088
rect 0 31152 800 31272
rect 59200 31152 60000 31272
rect 0 30336 800 30456
rect 59200 30336 60000 30456
rect 0 29520 800 29640
rect 59200 29520 60000 29640
rect 0 28704 800 28824
rect 59200 28704 60000 28824
rect 0 27888 800 28008
rect 59200 27888 60000 28008
rect 0 27072 800 27192
rect 59200 27072 60000 27192
rect 0 26256 800 26376
rect 59200 26256 60000 26376
rect 0 25440 800 25560
rect 59200 25440 60000 25560
rect 0 24624 800 24744
rect 59200 24624 60000 24744
rect 0 23808 800 23928
rect 59200 23808 60000 23928
rect 0 22992 800 23112
rect 59200 22992 60000 23112
rect 0 22176 800 22296
rect 59200 22176 60000 22296
rect 0 21360 800 21480
rect 59200 21360 60000 21480
rect 0 20544 800 20664
rect 59200 20544 60000 20664
rect 0 19728 800 19848
rect 59200 19728 60000 19848
rect 0 18912 800 19032
rect 59200 18912 60000 19032
rect 0 18096 800 18216
rect 59200 18096 60000 18216
rect 0 17280 800 17400
rect 59200 17280 60000 17400
rect 0 16464 800 16584
rect 59200 16464 60000 16584
rect 0 15648 800 15768
rect 59200 15648 60000 15768
rect 0 14832 800 14952
rect 59200 14832 60000 14952
rect 0 14016 800 14136
rect 59200 14016 60000 14136
rect 0 13200 800 13320
rect 59200 13200 60000 13320
rect 0 12384 800 12504
rect 59200 12384 60000 12504
rect 0 11568 800 11688
rect 59200 11568 60000 11688
rect 0 10752 800 10872
rect 59200 10752 60000 10872
rect 0 9936 800 10056
rect 59200 9936 60000 10056
rect 0 9120 800 9240
rect 59200 9120 60000 9240
rect 0 8304 800 8424
rect 59200 8304 60000 8424
rect 0 7488 800 7608
rect 59200 7488 60000 7608
rect 0 6672 800 6792
rect 59200 6672 60000 6792
rect 0 5856 800 5976
rect 59200 5856 60000 5976
rect 0 5040 800 5160
rect 59200 5040 60000 5160
rect 0 4224 800 4344
rect 59200 4224 60000 4344
rect 59200 3408 60000 3528
rect 59200 2592 60000 2712
rect 59200 1776 60000 1896
rect 59200 960 60000 1080
<< obsm3 >>
rect 800 58816 59120 58989
rect 800 58280 59200 58816
rect 800 58000 59120 58280
rect 800 57464 59200 58000
rect 800 57184 59120 57464
rect 800 56648 59200 57184
rect 800 56368 59120 56648
rect 800 55832 59200 56368
rect 880 55552 59120 55832
rect 800 55016 59200 55552
rect 880 54736 59120 55016
rect 800 54200 59200 54736
rect 880 53920 59120 54200
rect 800 53384 59200 53920
rect 880 53104 59120 53384
rect 800 52568 59200 53104
rect 880 52288 59120 52568
rect 800 51752 59200 52288
rect 880 51472 59120 51752
rect 800 50936 59200 51472
rect 880 50656 59120 50936
rect 800 50120 59200 50656
rect 880 49840 59120 50120
rect 800 49304 59200 49840
rect 880 49024 59120 49304
rect 800 48488 59200 49024
rect 880 48208 59120 48488
rect 800 47672 59200 48208
rect 880 47392 59120 47672
rect 800 46856 59200 47392
rect 880 46576 59120 46856
rect 800 46040 59200 46576
rect 880 45760 59120 46040
rect 800 45224 59200 45760
rect 880 44944 59120 45224
rect 800 44408 59200 44944
rect 880 44128 59120 44408
rect 800 43592 59200 44128
rect 880 43312 59120 43592
rect 800 42776 59200 43312
rect 880 42496 59120 42776
rect 800 41960 59200 42496
rect 880 41680 59120 41960
rect 800 41144 59200 41680
rect 880 40864 59120 41144
rect 800 40328 59200 40864
rect 880 40048 59120 40328
rect 800 39512 59200 40048
rect 880 39232 59120 39512
rect 800 38696 59200 39232
rect 880 38416 59120 38696
rect 800 37880 59200 38416
rect 880 37600 59120 37880
rect 800 37064 59200 37600
rect 880 36784 59120 37064
rect 800 36248 59200 36784
rect 880 35968 59120 36248
rect 800 35432 59200 35968
rect 880 35152 59120 35432
rect 800 34616 59200 35152
rect 880 34336 59120 34616
rect 800 33800 59200 34336
rect 880 33520 59120 33800
rect 800 32984 59200 33520
rect 880 32704 59120 32984
rect 800 32168 59200 32704
rect 880 31888 59120 32168
rect 800 31352 59200 31888
rect 880 31072 59120 31352
rect 800 30536 59200 31072
rect 880 30256 59120 30536
rect 800 29720 59200 30256
rect 880 29440 59120 29720
rect 800 28904 59200 29440
rect 880 28624 59120 28904
rect 800 28088 59200 28624
rect 880 27808 59120 28088
rect 800 27272 59200 27808
rect 880 26992 59120 27272
rect 800 26456 59200 26992
rect 880 26176 59120 26456
rect 800 25640 59200 26176
rect 880 25360 59120 25640
rect 800 24824 59200 25360
rect 880 24544 59120 24824
rect 800 24008 59200 24544
rect 880 23728 59120 24008
rect 800 23192 59200 23728
rect 880 22912 59120 23192
rect 800 22376 59200 22912
rect 880 22096 59120 22376
rect 800 21560 59200 22096
rect 880 21280 59120 21560
rect 800 20744 59200 21280
rect 880 20464 59120 20744
rect 800 19928 59200 20464
rect 880 19648 59120 19928
rect 800 19112 59200 19648
rect 880 18832 59120 19112
rect 800 18296 59200 18832
rect 880 18016 59120 18296
rect 800 17480 59200 18016
rect 880 17200 59120 17480
rect 800 16664 59200 17200
rect 880 16384 59120 16664
rect 800 15848 59200 16384
rect 880 15568 59120 15848
rect 800 15032 59200 15568
rect 880 14752 59120 15032
rect 800 14216 59200 14752
rect 880 13936 59120 14216
rect 800 13400 59200 13936
rect 880 13120 59120 13400
rect 800 12584 59200 13120
rect 880 12304 59120 12584
rect 800 11768 59200 12304
rect 880 11488 59120 11768
rect 800 10952 59200 11488
rect 880 10672 59120 10952
rect 800 10136 59200 10672
rect 880 9856 59120 10136
rect 800 9320 59200 9856
rect 880 9040 59120 9320
rect 800 8504 59200 9040
rect 880 8224 59120 8504
rect 800 7688 59200 8224
rect 880 7408 59120 7688
rect 800 6872 59200 7408
rect 880 6592 59120 6872
rect 800 6056 59200 6592
rect 880 5776 59120 6056
rect 800 5240 59200 5776
rect 880 4960 59120 5240
rect 800 4424 59200 4960
rect 880 4144 59120 4424
rect 800 3608 59200 4144
rect 800 3328 59120 3608
rect 800 2792 59200 3328
rect 800 2512 59120 2792
rect 800 1976 59200 2512
rect 800 1696 59120 1976
rect 800 1160 59200 1696
rect 800 987 59120 1160
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< labels >>
rlabel metal2 s 56414 0 56470 800 6 loopback_i
port 1 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 loopback_o
port 2 nsew signal output
rlabel metal2 s 1858 59200 1914 60000 6 mux0_i[0]
port 3 nsew signal input
rlabel metal2 s 3054 59200 3110 60000 6 mux0_i[1]
port 4 nsew signal input
rlabel metal2 s 4250 59200 4306 60000 6 mux0_i[2]
port 5 nsew signal input
rlabel metal2 s 5446 59200 5502 60000 6 mux0_i[3]
port 6 nsew signal input
rlabel metal2 s 6642 59200 6698 60000 6 mux0_i[4]
port 7 nsew signal input
rlabel metal2 s 7838 59200 7894 60000 6 mux0_i[5]
port 8 nsew signal input
rlabel metal2 s 9034 59200 9090 60000 6 mux1_i[0]
port 9 nsew signal input
rlabel metal2 s 10230 59200 10286 60000 6 mux1_i[1]
port 10 nsew signal input
rlabel metal2 s 11426 59200 11482 60000 6 mux1_i[2]
port 11 nsew signal input
rlabel metal2 s 12622 59200 12678 60000 6 mux1_i[3]
port 12 nsew signal input
rlabel metal2 s 13818 59200 13874 60000 6 mux1_i[4]
port 13 nsew signal input
rlabel metal2 s 15014 59200 15070 60000 6 mux1_i[5]
port 14 nsew signal input
rlabel metal2 s 16210 59200 16266 60000 6 mux2_i[0]
port 15 nsew signal input
rlabel metal2 s 17406 59200 17462 60000 6 mux2_i[1]
port 16 nsew signal input
rlabel metal2 s 18602 59200 18658 60000 6 mux2_i[2]
port 17 nsew signal input
rlabel metal2 s 19798 59200 19854 60000 6 mux2_i[3]
port 18 nsew signal input
rlabel metal2 s 20994 59200 21050 60000 6 mux2_i[4]
port 19 nsew signal input
rlabel metal2 s 22190 59200 22246 60000 6 mux2_i[5]
port 20 nsew signal input
rlabel metal2 s 23386 59200 23442 60000 6 mux3_i[0]
port 21 nsew signal input
rlabel metal2 s 24582 59200 24638 60000 6 mux3_i[1]
port 22 nsew signal input
rlabel metal2 s 25778 59200 25834 60000 6 mux3_i[2]
port 23 nsew signal input
rlabel metal2 s 26974 59200 27030 60000 6 mux3_i[3]
port 24 nsew signal input
rlabel metal2 s 28170 59200 28226 60000 6 mux3_i[4]
port 25 nsew signal input
rlabel metal2 s 29366 59200 29422 60000 6 mux3_i[5]
port 26 nsew signal input
rlabel metal2 s 30562 59200 30618 60000 6 mux4_i[0]
port 27 nsew signal input
rlabel metal2 s 31758 59200 31814 60000 6 mux4_i[1]
port 28 nsew signal input
rlabel metal2 s 32954 59200 33010 60000 6 mux4_i[2]
port 29 nsew signal input
rlabel metal2 s 34150 59200 34206 60000 6 mux4_i[3]
port 30 nsew signal input
rlabel metal2 s 35346 59200 35402 60000 6 mux4_i[4]
port 31 nsew signal input
rlabel metal2 s 36542 59200 36598 60000 6 mux4_i[5]
port 32 nsew signal input
rlabel metal2 s 37738 59200 37794 60000 6 mux5_i[0]
port 33 nsew signal input
rlabel metal2 s 38934 59200 38990 60000 6 mux5_i[1]
port 34 nsew signal input
rlabel metal2 s 40130 59200 40186 60000 6 mux5_i[2]
port 35 nsew signal input
rlabel metal2 s 41326 59200 41382 60000 6 mux5_i[3]
port 36 nsew signal input
rlabel metal2 s 42522 59200 42578 60000 6 mux5_i[4]
port 37 nsew signal input
rlabel metal2 s 43718 59200 43774 60000 6 mux5_i[5]
port 38 nsew signal input
rlabel metal2 s 44914 59200 44970 60000 6 mux6_i[0]
port 39 nsew signal input
rlabel metal2 s 46110 59200 46166 60000 6 mux6_i[1]
port 40 nsew signal input
rlabel metal2 s 47306 59200 47362 60000 6 mux6_i[2]
port 41 nsew signal input
rlabel metal2 s 48502 59200 48558 60000 6 mux6_i[3]
port 42 nsew signal input
rlabel metal2 s 49698 59200 49754 60000 6 mux6_i[4]
port 43 nsew signal input
rlabel metal2 s 50894 59200 50950 60000 6 mux6_i[5]
port 44 nsew signal input
rlabel metal2 s 52090 59200 52146 60000 6 mux7_i[0]
port 45 nsew signal input
rlabel metal2 s 53286 59200 53342 60000 6 mux7_i[1]
port 46 nsew signal input
rlabel metal2 s 54482 59200 54538 60000 6 mux7_i[2]
port 47 nsew signal input
rlabel metal2 s 55678 59200 55734 60000 6 mux7_i[3]
port 48 nsew signal input
rlabel metal2 s 56874 59200 56930 60000 6 mux7_i[4]
port 49 nsew signal input
rlabel metal2 s 58070 59200 58126 60000 6 mux7_i[5]
port 50 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 mux_adr_i[0]
port 51 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 mux_adr_i[1]
port 52 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 mux_adr_i[2]
port 53 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 mux_o[0]
port 54 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 mux_o[1]
port 55 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 mux_o[2]
port 56 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 mux_o[3]
port 57 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 mux_o[4]
port 58 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 mux_o[5]
port 59 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 reg0_o[0]
port 60 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 reg0_o[10]
port 61 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 reg0_o[11]
port 62 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 reg0_o[12]
port 63 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 reg0_o[13]
port 64 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 reg0_o[14]
port 65 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 reg0_o[15]
port 66 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 reg0_o[1]
port 67 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 reg0_o[2]
port 68 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 reg0_o[3]
port 69 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 reg0_o[4]
port 70 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 reg0_o[5]
port 71 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 reg0_o[6]
port 72 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 reg0_o[7]
port 73 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 reg0_o[8]
port 74 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 reg0_o[9]
port 75 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 reg1_o[0]
port 76 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 reg1_o[10]
port 77 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 reg1_o[11]
port 78 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 reg1_o[12]
port 79 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 reg1_o[13]
port 80 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 reg1_o[14]
port 81 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 reg1_o[15]
port 82 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 reg1_o[1]
port 83 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 reg1_o[2]
port 84 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 reg1_o[3]
port 85 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 reg1_o[4]
port 86 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 reg1_o[5]
port 87 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 reg1_o[6]
port 88 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 reg1_o[7]
port 89 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 reg1_o[8]
port 90 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 reg1_o[9]
port 91 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 reg2_o[0]
port 92 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 reg2_o[10]
port 93 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 reg2_o[11]
port 94 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 reg2_o[12]
port 95 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 reg2_o[13]
port 96 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 reg2_o[14]
port 97 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 reg2_o[15]
port 98 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 reg2_o[1]
port 99 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 reg2_o[2]
port 100 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 reg2_o[3]
port 101 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 reg2_o[4]
port 102 nsew signal output
rlabel metal3 s 0 34416 800 34536 6 reg2_o[5]
port 103 nsew signal output
rlabel metal3 s 0 35232 800 35352 6 reg2_o[6]
port 104 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 reg2_o[7]
port 105 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 reg2_o[8]
port 106 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 reg2_o[9]
port 107 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 reg3_o[0]
port 108 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 reg3_o[10]
port 109 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 reg3_o[11]
port 110 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 reg3_o[12]
port 111 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 reg3_o[13]
port 112 nsew signal output
rlabel metal3 s 0 54816 800 54936 6 reg3_o[14]
port 113 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 reg3_o[15]
port 114 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 reg3_o[1]
port 115 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 reg3_o[2]
port 116 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 reg3_o[3]
port 117 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 reg3_o[4]
port 118 nsew signal output
rlabel metal3 s 0 47472 800 47592 6 reg3_o[5]
port 119 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 reg3_o[6]
port 120 nsew signal output
rlabel metal3 s 0 49104 800 49224 6 reg3_o[7]
port 121 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 reg3_o[8]
port 122 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 reg3_o[9]
port 123 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 reg_adr_i[0]
port 124 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 reg_adr_i[1]
port 125 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 reg_dat_i[0]
port 126 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 reg_dat_i[10]
port 127 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 reg_dat_i[11]
port 128 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 reg_dat_i[12]
port 129 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 reg_dat_i[13]
port 130 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 reg_dat_i[14]
port 131 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 reg_dat_i[15]
port 132 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 reg_dat_i[1]
port 133 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 reg_dat_i[2]
port 134 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 reg_dat_i[3]
port 135 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 reg_dat_i[4]
port 136 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 reg_dat_i[5]
port 137 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 reg_dat_i[6]
port 138 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 reg_dat_i[7]
port 139 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 reg_dat_i[8]
port 140 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 reg_dat_i[9]
port 141 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 reg_wr_i
port 142 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 rst_n_i
port 143 nsew signal input
rlabel metal3 s 59200 960 60000 1080 6 temp0_dac_i[0]
port 144 nsew signal input
rlabel metal3 s 59200 1776 60000 1896 6 temp0_dac_i[1]
port 145 nsew signal input
rlabel metal3 s 59200 2592 60000 2712 6 temp0_dac_i[2]
port 146 nsew signal input
rlabel metal3 s 59200 3408 60000 3528 6 temp0_dac_i[3]
port 147 nsew signal input
rlabel metal3 s 59200 4224 60000 4344 6 temp0_dac_i[4]
port 148 nsew signal input
rlabel metal3 s 59200 5040 60000 5160 6 temp0_dac_i[5]
port 149 nsew signal input
rlabel metal3 s 59200 20544 60000 20664 6 temp0_ticks_i[0]
port 150 nsew signal input
rlabel metal3 s 59200 28704 60000 28824 6 temp0_ticks_i[10]
port 151 nsew signal input
rlabel metal3 s 59200 29520 60000 29640 6 temp0_ticks_i[11]
port 152 nsew signal input
rlabel metal3 s 59200 21360 60000 21480 6 temp0_ticks_i[1]
port 153 nsew signal input
rlabel metal3 s 59200 22176 60000 22296 6 temp0_ticks_i[2]
port 154 nsew signal input
rlabel metal3 s 59200 22992 60000 23112 6 temp0_ticks_i[3]
port 155 nsew signal input
rlabel metal3 s 59200 23808 60000 23928 6 temp0_ticks_i[4]
port 156 nsew signal input
rlabel metal3 s 59200 24624 60000 24744 6 temp0_ticks_i[5]
port 157 nsew signal input
rlabel metal3 s 59200 25440 60000 25560 6 temp0_ticks_i[6]
port 158 nsew signal input
rlabel metal3 s 59200 26256 60000 26376 6 temp0_ticks_i[7]
port 159 nsew signal input
rlabel metal3 s 59200 27072 60000 27192 6 temp0_ticks_i[8]
port 160 nsew signal input
rlabel metal3 s 59200 27888 60000 28008 6 temp0_ticks_i[9]
port 161 nsew signal input
rlabel metal3 s 59200 5856 60000 5976 6 temp1_dac_i[0]
port 162 nsew signal input
rlabel metal3 s 59200 6672 60000 6792 6 temp1_dac_i[1]
port 163 nsew signal input
rlabel metal3 s 59200 7488 60000 7608 6 temp1_dac_i[2]
port 164 nsew signal input
rlabel metal3 s 59200 8304 60000 8424 6 temp1_dac_i[3]
port 165 nsew signal input
rlabel metal3 s 59200 9120 60000 9240 6 temp1_dac_i[4]
port 166 nsew signal input
rlabel metal3 s 59200 9936 60000 10056 6 temp1_dac_i[5]
port 167 nsew signal input
rlabel metal3 s 59200 30336 60000 30456 6 temp1_ticks_i[0]
port 168 nsew signal input
rlabel metal3 s 59200 38496 60000 38616 6 temp1_ticks_i[10]
port 169 nsew signal input
rlabel metal3 s 59200 39312 60000 39432 6 temp1_ticks_i[11]
port 170 nsew signal input
rlabel metal3 s 59200 31152 60000 31272 6 temp1_ticks_i[1]
port 171 nsew signal input
rlabel metal3 s 59200 31968 60000 32088 6 temp1_ticks_i[2]
port 172 nsew signal input
rlabel metal3 s 59200 32784 60000 32904 6 temp1_ticks_i[3]
port 173 nsew signal input
rlabel metal3 s 59200 33600 60000 33720 6 temp1_ticks_i[4]
port 174 nsew signal input
rlabel metal3 s 59200 34416 60000 34536 6 temp1_ticks_i[5]
port 175 nsew signal input
rlabel metal3 s 59200 35232 60000 35352 6 temp1_ticks_i[6]
port 176 nsew signal input
rlabel metal3 s 59200 36048 60000 36168 6 temp1_ticks_i[7]
port 177 nsew signal input
rlabel metal3 s 59200 36864 60000 36984 6 temp1_ticks_i[8]
port 178 nsew signal input
rlabel metal3 s 59200 37680 60000 37800 6 temp1_ticks_i[9]
port 179 nsew signal input
rlabel metal3 s 59200 10752 60000 10872 6 temp2_dac_i[0]
port 180 nsew signal input
rlabel metal3 s 59200 11568 60000 11688 6 temp2_dac_i[1]
port 181 nsew signal input
rlabel metal3 s 59200 12384 60000 12504 6 temp2_dac_i[2]
port 182 nsew signal input
rlabel metal3 s 59200 13200 60000 13320 6 temp2_dac_i[3]
port 183 nsew signal input
rlabel metal3 s 59200 14016 60000 14136 6 temp2_dac_i[4]
port 184 nsew signal input
rlabel metal3 s 59200 14832 60000 14952 6 temp2_dac_i[5]
port 185 nsew signal input
rlabel metal3 s 59200 40128 60000 40248 6 temp2_ticks_i[0]
port 186 nsew signal input
rlabel metal3 s 59200 48288 60000 48408 6 temp2_ticks_i[10]
port 187 nsew signal input
rlabel metal3 s 59200 49104 60000 49224 6 temp2_ticks_i[11]
port 188 nsew signal input
rlabel metal3 s 59200 40944 60000 41064 6 temp2_ticks_i[1]
port 189 nsew signal input
rlabel metal3 s 59200 41760 60000 41880 6 temp2_ticks_i[2]
port 190 nsew signal input
rlabel metal3 s 59200 42576 60000 42696 6 temp2_ticks_i[3]
port 191 nsew signal input
rlabel metal3 s 59200 43392 60000 43512 6 temp2_ticks_i[4]
port 192 nsew signal input
rlabel metal3 s 59200 44208 60000 44328 6 temp2_ticks_i[5]
port 193 nsew signal input
rlabel metal3 s 59200 45024 60000 45144 6 temp2_ticks_i[6]
port 194 nsew signal input
rlabel metal3 s 59200 45840 60000 45960 6 temp2_ticks_i[7]
port 195 nsew signal input
rlabel metal3 s 59200 46656 60000 46776 6 temp2_ticks_i[8]
port 196 nsew signal input
rlabel metal3 s 59200 47472 60000 47592 6 temp2_ticks_i[9]
port 197 nsew signal input
rlabel metal3 s 59200 15648 60000 15768 6 temp3_dac_i[0]
port 198 nsew signal input
rlabel metal3 s 59200 16464 60000 16584 6 temp3_dac_i[1]
port 199 nsew signal input
rlabel metal3 s 59200 17280 60000 17400 6 temp3_dac_i[2]
port 200 nsew signal input
rlabel metal3 s 59200 18096 60000 18216 6 temp3_dac_i[3]
port 201 nsew signal input
rlabel metal3 s 59200 18912 60000 19032 6 temp3_dac_i[4]
port 202 nsew signal input
rlabel metal3 s 59200 19728 60000 19848 6 temp3_dac_i[5]
port 203 nsew signal input
rlabel metal3 s 59200 49920 60000 50040 6 temp3_ticks_i[0]
port 204 nsew signal input
rlabel metal3 s 59200 58080 60000 58200 6 temp3_ticks_i[10]
port 205 nsew signal input
rlabel metal3 s 59200 58896 60000 59016 6 temp3_ticks_i[11]
port 206 nsew signal input
rlabel metal3 s 59200 50736 60000 50856 6 temp3_ticks_i[1]
port 207 nsew signal input
rlabel metal3 s 59200 51552 60000 51672 6 temp3_ticks_i[2]
port 208 nsew signal input
rlabel metal3 s 59200 52368 60000 52488 6 temp3_ticks_i[3]
port 209 nsew signal input
rlabel metal3 s 59200 53184 60000 53304 6 temp3_ticks_i[4]
port 210 nsew signal input
rlabel metal3 s 59200 54000 60000 54120 6 temp3_ticks_i[5]
port 211 nsew signal input
rlabel metal3 s 59200 54816 60000 54936 6 temp3_ticks_i[6]
port 212 nsew signal input
rlabel metal3 s 59200 55632 60000 55752 6 temp3_ticks_i[7]
port 213 nsew signal input
rlabel metal3 s 59200 56448 60000 56568 6 temp3_ticks_i[8]
port 214 nsew signal input
rlabel metal3 s 59200 57264 60000 57384 6 temp3_ticks_i[9]
port 215 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 temp_dac_o[0]
port 216 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 temp_dac_o[1]
port 217 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 temp_dac_o[2]
port 218 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 temp_dac_o[3]
port 219 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 temp_dac_o[4]
port 220 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 temp_dac_o[5]
port 221 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 temp_sel_i[0]
port 222 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 temp_sel_i[1]
port 223 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 temp_ticks_o[0]
port 224 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 temp_ticks_o[10]
port 225 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 temp_ticks_o[11]
port 226 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 temp_ticks_o[1]
port 227 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 temp_ticks_o[2]
port 228 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 temp_ticks_o[3]
port 229 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 temp_ticks_o[4]
port 230 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 temp_ticks_o[5]
port 231 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 temp_ticks_o[6]
port 232 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 temp_ticks_o[7]
port 233 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 temp_ticks_o[8]
port 234 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 temp_ticks_o[9]
port 235 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 236 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 236 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 237 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 237 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2608062
string GDS_FILE /home/harald/mpw8-submission/openlane/config_reg_mux/runs/22_12_09_21_46/results/signoff/config_reg_mux.magic.gds
string GDS_START 270676
<< end >>

